LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L3WROM IS
    PORT (
        weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
        address : IN unsigned(weightsbitsAddress(3) DOWNTO 0));
END L3WROM;

ARCHITECTURE RTL OF L3WROM IS

    TYPE ROM_mem IS ARRAY (0 TO 2047) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem := (0=>"100110110",
    1=>"000110110",
    2=>"011011011",
    3=>"100100100",
    4=>"010111111",
    5=>"001001010",
    6=>"110110110",
    7=>"011010010",
    8=>"110010110",
    9=>"011001010",
    10=>"010011011",
    11=>"001001010",
    12=>"000010000",
    13=>"000100101",
    14=>"001001001",
    15=>"010110110",
    16=>"110110110",
    17=>"101101001",
    18=>"100001011",
    19=>"001111010",
    20=>"001001001",
    21=>"110110110",
    22=>"110110100",
    23=>"001101001",
    24=>"001001011",
    25=>"100100101",
    26=>"001001011",
    27=>"100100000",
    28=>"011000011",
    29=>"110110110",
    30=>"001000011",
    31=>"011011011",
    32=>"100100111",
    33=>"000100101",
    34=>"111000000",
    35=>"000000111",
    36=>"000111011",
    37=>"000111100",
    38=>"101111111",
    39=>"000100110",
    40=>"111000000",
    41=>"000000001",
    42=>"010000111",
    43=>"101000000",
    44=>"000001000",
    45=>"100001000",
    46=>"011001111",
    47=>"001011101",
    48=>"110010000",
    49=>"000111111",
    50=>"001101100",
    51=>"111000000",
    52=>"100000111",
    53=>"000111111",
    54=>"101111100",
    55=>"110001000",
    56=>"100001111",
    57=>"111100000",
    58=>"000111111",
    59=>"000010000",
    60=>"001100010",
    61=>"010000010",
    62=>"111010111",
    63=>"101001001",
    64=>"011001001",
    65=>"001011011",
    66=>"100100100",
    67=>"100101101",
    68=>"111001001",
    69=>"011011000",
    70=>"111101111",
    71=>"100100111",
    72=>"011001001",
    73=>"100100100",
    74=>"101111111",
    75=>"000000100",
    76=>"000000000",
    77=>"011000000",
    78=>"100110110",
    79=>"001101011",
    80=>"111111001",
    81=>"010001010",
    82=>"110000100",
    83=>"011011011",
    84=>"001001001",
    85=>"101100100",
    86=>"101111111",
    87=>"000100100",
    88=>"001001011",
    89=>"010010011",
    90=>"011011001",
    91=>"000000000",
    92=>"010011011",
    93=>"011001101",
    94=>"000100110",
    95=>"110101001",
    96=>"000000000",
    97=>"000010000",
    98=>"001101111",
    99=>"010000010",
    100=>"010111111",
    101=>"000000000",
    102=>"100100100",
    103=>"100100000",
    104=>"010101000",
    105=>"000110000",
    106=>"010110011",
    107=>"000111000",
    108=>"001001000",
    109=>"100101011",
    110=>"000111011",
    111=>"011011100",
    112=>"010101110",
    113=>"000010010",
    114=>"010110000",
    115=>"110111000",
    116=>"000100000",
    117=>"000110011",
    118=>"000000000",
    119=>"001100000",
    120=>"110000000",
    121=>"000001101",
    122=>"101111111",
    123=>"011011000",
    124=>"011011110",
    125=>"000000100",
    126=>"111000111",
    127=>"000000000",
    128=>"100101111",
    129=>"100101100",
    130=>"000000001",
    131=>"000000000",
    132=>"111101000",
    133=>"000001001",
    134=>"110111111",
    135=>"000100111",
    136=>"001000000",
    137=>"000100100",
    138=>"001000011",
    139=>"100100110",
    140=>"101001111",
    141=>"100000100",
    142=>"000000000",
    143=>"011111110",
    144=>"001101101",
    145=>"000100100",
    146=>"010000000",
    147=>"111111111",
    148=>"010001000",
    149=>"000000000",
    150=>"100101111",
    151=>"000000100",
    152=>"111110000",
    153=>"110111111",
    154=>"111111111",
    155=>"010111111",
    156=>"000000000",
    157=>"001111111",
    158=>"001001111",
    159=>"111110000",
    160=>"000111111",
    161=>"000000111",
    162=>"001001000",
    163=>"111110111",
    164=>"001001001",
    165=>"110011001",
    166=>"000111111",
    167=>"000110110",
    168=>"010111011",
    169=>"111001000",
    170=>"000000000",
    171=>"011001000",
    172=>"011000000",
    173=>"111110100",
    174=>"000110010",
    175=>"110111111",
    176=>"011011001",
    177=>"111100100",
    178=>"000000100",
    179=>"110111011",
    180=>"011001001",
    181=>"100110111",
    182=>"111111111",
    183=>"011000000",
    184=>"011000100",
    185=>"110110111",
    186=>"000000000",
    187=>"110110111",
    188=>"111011000",
    189=>"000111011",
    190=>"111000000",
    191=>"111001000",
    192=>"011100001",
    193=>"100101000",
    194=>"011100000",
    195=>"100101011",
    196=>"000001110",
    197=>"000111110",
    198=>"111111000",
    199=>"111111100",
    200=>"000111100",
    201=>"100001111",
    202=>"000111100",
    203=>"000110100",
    204=>"000001000",
    205=>"100001111",
    206=>"000001111",
    207=>"011001000",
    208=>"001111100",
    209=>"110000011",
    210=>"000011110",
    211=>"000011110",
    212=>"001110000",
    213=>"011100000",
    214=>"000000011",
    215=>"000000111",
    216=>"001110100",
    217=>"110000011",
    218=>"011110000",
    219=>"000000001",
    220=>"111000111",
    221=>"011110000",
    222=>"000011110",
    223=>"011100110",
    224=>"101001001",
    225=>"101101100",
    226=>"011100011",
    227=>"000000000",
    228=>"110000101",
    229=>"100100110",
    230=>"111000000",
    231=>"111101001",
    232=>"100000000",
    233=>"010110110",
    234=>"111111111",
    235=>"100000001",
    236=>"101000001",
    237=>"000000000",
    238=>"111111111",
    239=>"000001011",
    240=>"101001011",
    241=>"011010110",
    242=>"110101000",
    243=>"000000000",
    244=>"110101101",
    245=>"000000001",
    246=>"100001001",
    247=>"111110110",
    248=>"111111111",
    249=>"000110100",
    250=>"111110100",
    251=>"000000001",
    252=>"010100111",
    253=>"101001001",
    254=>"000111111",
    255=>"110110110",
    256=>"111001000",
    257=>"000101111",
    258=>"100110111",
    259=>"011000100",
    260=>"000000000",
    261=>"100100111",
    262=>"100111011",
    263=>"001001111",
    264=>"110111011",
    265=>"011001100",
    266=>"111111111",
    267=>"001001000",
    268=>"011000000",
    269=>"011111101",
    270=>"011001100",
    271=>"111001001",
    272=>"000000000",
    273=>"000011001",
    274=>"001100110",
    275=>"100110111",
    276=>"001000000",
    277=>"011001100",
    278=>"111101101",
    279=>"111100100",
    280=>"100110111",
    281=>"100110011",
    282=>"000110011",
    283=>"000100110",
    284=>"100110111",
    285=>"001000010",
    286=>"000000111",
    287=>"111001010",
    288=>"000101001",
    289=>"100101100",
    290=>"001000000",
    291=>"000000000",
    292=>"001101111",
    293=>"000101001",
    294=>"100000111",
    295=>"101101101",
    296=>"111111101",
    297=>"001101101",
    298=>"000000100",
    299=>"000000000",
    300=>"101001000",
    301=>"011001011",
    302=>"000000000",
    303=>"000100111",
    304=>"011010111",
    305=>"101000111",
    306=>"000101101",
    307=>"111101101",
    308=>"000001101",
    309=>"011111111",
    310=>"000000000",
    311=>"000000011",
    312=>"100100010",
    313=>"000000100",
    314=>"000100100",
    315=>"101000010",
    316=>"010001110",
    317=>"101100101",
    318=>"000000010",
    319=>"111111111",
    320=>"100001011",
    321=>"100001011",
    322=>"011010001",
    323=>"110111111",
    324=>"110000000",
    325=>"100101111",
    326=>"011111111",
    327=>"001001011",
    328=>"111111000",
    329=>"110100111",
    330=>"100110110",
    331=>"000001001",
    332=>"100100000",
    333=>"011111110",
    334=>"011111111",
    335=>"011001011",
    336=>"000111011",
    337=>"000001001",
    338=>"111100010",
    339=>"111111111",
    340=>"100000000",
    341=>"000000000",
    342=>"001001001",
    343=>"011110110",
    344=>"100001000",
    345=>"000000000",
    346=>"100000001",
    347=>"110111110",
    348=>"000000000",
    349=>"100000100",
    350=>"110111111",
    351=>"111000010",
    352=>"011001001",
    353=>"100100110",
    354=>"000000000",
    355=>"110110110",
    356=>"001000100",
    357=>"000100110",
    358=>"110110001",
    359=>"011011001",
    360=>"100110100",
    361=>"011011001",
    362=>"010011110",
    363=>"011011001",
    364=>"001001101",
    365=>"010000010",
    366=>"101101111",
    367=>"101100101",
    368=>"000110111",
    369=>"011000110",
    370=>"110011000",
    371=>"100000100",
    372=>"100100110",
    373=>"111011000",
    374=>"001000001",
    375=>"011010010",
    376=>"111101111",
    377=>"111001111",
    378=>"000101100",
    379=>"011111001",
    380=>"100110110",
    381=>"001100101",
    382=>"010011010",
    383=>"001101100",
    384=>"000010010",
    385=>"000011000",
    386=>"100100000",
    387=>"001011110",
    388=>"111111011",
    389=>"000010010",
    390=>"001011101",
    391=>"000011000",
    392=>"110000000",
    393=>"010111000",
    394=>"000010000",
    395=>"000110000",
    396=>"010010000",
    397=>"010010010",
    398=>"001011000",
    399=>"010110010",
    400=>"000011000",
    401=>"010010010",
    402=>"000011000",
    403=>"111011010",
    404=>"000011000",
    405=>"000011000",
    406=>"010010010",
    407=>"000110000",
    408=>"000010011",
    409=>"001111000",
    410=>"100110001",
    411=>"000000010",
    412=>"100011001",
    413=>"000101001",
    414=>"111010111",
    415=>"000111010",
    416=>"111010010",
    417=>"010001011",
    418=>"100000010",
    419=>"001001100",
    420=>"111000011",
    421=>"001000011",
    422=>"111000111",
    423=>"010011001",
    424=>"011010000",
    425=>"000111001",
    426=>"110010011",
    427=>"110001000",
    428=>"000000000",
    429=>"011101100",
    430=>"111000111",
    431=>"000000110",
    432=>"010010110",
    433=>"101101101",
    434=>"011011000",
    435=>"101000011",
    436=>"000010010",
    437=>"111000000",
    438=>"101000101",
    439=>"000111000",
    440=>"100111011",
    441=>"011001100",
    442=>"110100001",
    443=>"011000100",
    444=>"000111000",
    445=>"110000111",
    446=>"000111001",
    447=>"000111011",
    448=>"100100110",
    449=>"011001001",
    450=>"010111001",
    451=>"110011011",
    452=>"001000000",
    453=>"011001000",
    454=>"110001101",
    455=>"100110110",
    456=>"111111000",
    457=>"100110110",
    458=>"111111111",
    459=>"001100100",
    460=>"000100100",
    461=>"010000010",
    462=>"101100011",
    463=>"111001101",
    464=>"010001110",
    465=>"010010010",
    466=>"111011001",
    467=>"111110000",
    468=>"011111010",
    469=>"111011010",
    470=>"011000100",
    471=>"001110000",
    472=>"011111110",
    473=>"101101111",
    474=>"000100100",
    475=>"111011011",
    476=>"011011101",
    477=>"100101100",
    478=>"000000110",
    479=>"010010000",
    480=>"100100110",
    481=>"101101000",
    482=>"111111101",
    483=>"111111111",
    484=>"000000001",
    485=>"101111111",
    486=>"111000100",
    487=>"101111001",
    488=>"000000000",
    489=>"111101001",
    490=>"111111111",
    491=>"101001000",
    492=>"110000000",
    493=>"111111111",
    494=>"110101001",
    495=>"011101110",
    496=>"000000000",
    497=>"100000100",
    498=>"111000000",
    499=>"100101011",
    500=>"100001011",
    501=>"100011101",
    502=>"001101101",
    503=>"000000000",
    504=>"111111111",
    505=>"001100110",
    506=>"101011010",
    507=>"011101110",
    508=>"001000000",
    509=>"000000000",
    510=>"000000000",
    511=>"110111001",
    512=>"100001111",
    513=>"000101101",
    514=>"011100100",
    515=>"110001000",
    516=>"100111000",
    517=>"111011000",
    518=>"111000000",
    519=>"110110101",
    520=>"101111000",
    521=>"010000111",
    522=>"111110000",
    523=>"100000000",
    524=>"000001000",
    525=>"001000001",
    526=>"111100110",
    527=>"111001001",
    528=>"111001000",
    529=>"000110111",
    530=>"110111000",
    531=>"010000010",
    532=>"111000010",
    533=>"111000000",
    534=>"000111111",
    535=>"000111111",
    536=>"100110111",
    537=>"111001101",
    538=>"111111010",
    539=>"111001000",
    540=>"000111111",
    541=>"111000000",
    542=>"000111111",
    543=>"000000110",
    544=>"010010010",
    545=>"010000010",
    546=>"100010011",
    547=>"001000101",
    548=>"111010100",
    549=>"011000010",
    550=>"111111000",
    551=>"010010011",
    552=>"111000000",
    553=>"000010010",
    554=>"111111111",
    555=>"000000011",
    556=>"000000001",
    557=>"011011111",
    558=>"000000011",
    559=>"011001000",
    560=>"011011001",
    561=>"001000100",
    562=>"110110011",
    563=>"111111111",
    564=>"000000011",
    565=>"111111110",
    566=>"010000111",
    567=>"000000000",
    568=>"001111111",
    569=>"000010000",
    570=>"100000100",
    571=>"111111111",
    572=>"000000000",
    573=>"101101000",
    574=>"000000000",
    575=>"010101111",
    576=>"100100100",
    577=>"010011001",
    578=>"101100110",
    579=>"011001001",
    580=>"100110110",
    581=>"010001001",
    582=>"101110110",
    583=>"000011001",
    584=>"110010000",
    585=>"010000001",
    586=>"100110111",
    587=>"010010000",
    588=>"001100000",
    589=>"011011000",
    590=>"001001100",
    591=>"110010001",
    592=>"100110110",
    593=>"011001100",
    594=>"011001001",
    595=>"010010010",
    596=>"000001011",
    597=>"001001001",
    598=>"100100110",
    599=>"011101100",
    600=>"100100111",
    601=>"110011001",
    602=>"100110111",
    603=>"110001000",
    604=>"011000001",
    605=>"100110010",
    606=>"010000001",
    607=>"011011011",
    608=>"000100101",
    609=>"001100001",
    610=>"011100000",
    611=>"100001111",
    612=>"001110100",
    613=>"001110100",
    614=>"100011010",
    615=>"000110001",
    616=>"001011100",
    617=>"001110000",
    618=>"111110000",
    619=>"011100000",
    620=>"001000000",
    621=>"101001111",
    622=>"111000001",
    623=>"010010101",
    624=>"000100000",
    625=>"100001111",
    626=>"011110000",
    627=>"110100011",
    628=>"111100000",
    629=>"001011110",
    630=>"110000001",
    631=>"100000110",
    632=>"000100100",
    633=>"100001111",
    634=>"010110100",
    635=>"000001100",
    636=>"000011110",
    637=>"010110010",
    638=>"000001101",
    639=>"011100001",
    640=>"011011010",
    641=>"011001011",
    642=>"000011011",
    643=>"000100100",
    644=>"110011010",
    645=>"100100111",
    646=>"111011001",
    647=>"000100110",
    648=>"101101110",
    649=>"001100011",
    650=>"110111001",
    651=>"000000011",
    652=>"000000000",
    653=>"100110010",
    654=>"100100110",
    655=>"010011000",
    656=>"101101010",
    657=>"111011000",
    658=>"100111111",
    659=>"001010011",
    660=>"100100100",
    661=>"000110110",
    662=>"011011011",
    663=>"100011000",
    664=>"000011001",
    665=>"101110010",
    666=>"010000000",
    667=>"000100110",
    668=>"000111111",
    669=>"010010011",
    670=>"000011000",
    671=>"000100110",
    672=>"000010010",
    673=>"011011111",
    674=>"000000011",
    675=>"111111111",
    676=>"111110111",
    677=>"011101101",
    678=>"001000000",
    679=>"000111111",
    680=>"000000010",
    681=>"010111011",
    682=>"110100011",
    683=>"111111011",
    684=>"111111111",
    685=>"000000010",
    686=>"100110111",
    687=>"100111011",
    688=>"000000000",
    689=>"100010110",
    690=>"111111101",
    691=>"111111001",
    692=>"011001001",
    693=>"111111111",
    694=>"000000100",
    695=>"000111111",
    696=>"101110110",
    697=>"010011101",
    698=>"111111001",
    699=>"000000000",
    700=>"000100001",
    701=>"001011100",
    702=>"110011111",
    703=>"110111011",
    704=>"011111101",
    705=>"101100101",
    706=>"001000001",
    707=>"000000000",
    708=>"101100000",
    709=>"101100100",
    710=>"111111111",
    711=>"100101001",
    712=>"111000110",
    713=>"101101001",
    714=>"001010010",
    715=>"100100000",
    716=>"100000000",
    717=>"000000000",
    718=>"001000000",
    719=>"001001001",
    720=>"001011111",
    721=>"111011011",
    722=>"100100101",
    723=>"000000111",
    724=>"001000001",
    725=>"101111000",
    726=>"001000001",
    727=>"000000100",
    728=>"000000000",
    729=>"100000100",
    730=>"100000000",
    731=>"000110111",
    732=>"001001000",
    733=>"010010111",
    734=>"001000000",
    735=>"110100100",
    736=>"000000111",
    737=>"111100000",
    738=>"110000001",
    739=>"111101001",
    740=>"111111011",
    741=>"111000000",
    742=>"111100000",
    743=>"000000111",
    744=>"101101001",
    745=>"000010111",
    746=>"010110010",
    747=>"000001111",
    748=>"010001011",
    749=>"101011111",
    750=>"011111101",
    751=>"000000111",
    752=>"100000100",
    753=>"111000001",
    754=>"001010100",
    755=>"111101111",
    756=>"001000110",
    757=>"100000001",
    758=>"001000001",
    759=>"100000000",
    760=>"010111111",
    761=>"000011000",
    762=>"111110010",
    763=>"100110101",
    764=>"001000001",
    765=>"100001001",
    766=>"000011101",
    767=>"100000011",
    768=>"001101101",
    769=>"101100100",
    770=>"000000000",
    771=>"100000100",
    772=>"101111101",
    773=>"111010110",
    774=>"101101101",
    775=>"101100111",
    776=>"111111111",
    777=>"000000011",
    778=>"000000000",
    779=>"101100111",
    780=>"000000000",
    781=>"000000000",
    782=>"111100111",
    783=>"000110000",
    784=>"111111111",
    785=>"111000011",
    786=>"001000100",
    787=>"111001100",
    788=>"011111101",
    789=>"100111101",
    790=>"001000101",
    791=>"111000111",
    792=>"000000000",
    793=>"111001111",
    794=>"011011011",
    795=>"000000000",
    796=>"111000111",
    797=>"101101100",
    798=>"110111111",
    799=>"111000111",
    800=>"010010010",
    801=>"010010011",
    802=>"111110001",
    803=>"000000000",
    804=>"000001000",
    805=>"010011011",
    806=>"100100101",
    807=>"000011111",
    808=>"000000000",
    809=>"000011111",
    810=>"001000001",
    811=>"000000001",
    812=>"010000010",
    813=>"101100000",
    814=>"111111111",
    815=>"110111111",
    816=>"110100000",
    817=>"111100000",
    818=>"001001011",
    819=>"100100000",
    820=>"010000100",
    821=>"011001001",
    822=>"111100000",
    823=>"111100001",
    824=>"000000000",
    825=>"011111111",
    826=>"111110101",
    827=>"010001100",
    828=>"111011011",
    829=>"000101000",
    830=>"111100110",
    831=>"011111111",
    832=>"011110011",
    833=>"011110000",
    834=>"111111111",
    835=>"000000000",
    836=>"011111110",
    837=>"000010001",
    838=>"000111111",
    839=>"011010000",
    840=>"011011111",
    841=>"010000011",
    842=>"011111111",
    843=>"111000001",
    844=>"110000000",
    845=>"100000000",
    846=>"000011111",
    847=>"010100000",
    848=>"100101101",
    849=>"111000000",
    850=>"010000001",
    851=>"111111111",
    852=>"010110101",
    853=>"000001011",
    854=>"111110000",
    855=>"111100000",
    856=>"011011111",
    857=>"000000000",
    858=>"001011111",
    859=>"000000000",
    860=>"111000001",
    861=>"000111111",
    862=>"110000001",
    863=>"111000000",
    864=>"001001001",
    865=>"000001011",
    866=>"011011101",
    867=>"100111010",
    868=>"000111000",
    869=>"111100000",
    870=>"011110100",
    871=>"000011011",
    872=>"101100101",
    873=>"111100100",
    874=>"001111100",
    875=>"111010000",
    876=>"001111000",
    877=>"001111100",
    878=>"000100100",
    879=>"000000101",
    880=>"111110000",
    881=>"111100100",
    882=>"000111110",
    883=>"000000111",
    884=>"000001111",
    885=>"000000001",
    886=>"001011011",
    887=>"011100010",
    888=>"110111110",
    889=>"100101001",
    890=>"100100101",
    891=>"010101110",
    892=>"111110000",
    893=>"100101100",
    894=>"010110100",
    895=>"011001011",
    896=>"010000000",
    897=>"000000000",
    898=>"000001001",
    899=>"011111111",
    900=>"000000101",
    901=>"000000000",
    902=>"000010010",
    903=>"010000000",
    904=>"111000000",
    905=>"010111000",
    906=>"100011001",
    907=>"000000000",
    908=>"011111101",
    909=>"111110011",
    910=>"110110011",
    911=>"000110000",
    912=>"010100001",
    913=>"000011010",
    914=>"111111111",
    915=>"000000111",
    916=>"011111111",
    917=>"010110110",
    918=>"001000101",
    919=>"100110011",
    920=>"111011010",
    921=>"000100110",
    922=>"111011110",
    923=>"101000000",
    924=>"010011000",
    925=>"010011111",
    926=>"000101100",
    927=>"111011000",
    928=>"101100101",
    929=>"101000101",
    930=>"000000000",
    931=>"001101100",
    932=>"000000000",
    933=>"111001001",
    934=>"100000111",
    935=>"101000100",
    936=>"111000000",
    937=>"101000100",
    938=>"111111111",
    939=>"001000000",
    940=>"001000000",
    941=>"110010011",
    942=>"001001000",
    943=>"001000001",
    944=>"100111111",
    945=>"001000101",
    946=>"111101101",
    947=>"000000000",
    948=>"000000000",
    949=>"001000000",
    950=>"111111111",
    951=>"100100100",
    952=>"110110110",
    953=>"101101101",
    954=>"100000000",
    955=>"101101011",
    956=>"011001001",
    957=>"010010010",
    958=>"111111111",
    959=>"001000001",
    960=>"010000101",
    961=>"000000110",
    962=>"011100100",
    963=>"000111001",
    964=>"011100010",
    965=>"000110011",
    966=>"000111110",
    967=>"000100111",
    968=>"011110011",
    969=>"011000111",
    970=>"000001000",
    971=>"000000111",
    972=>"000000001",
    973=>"100000000",
    974=>"111111000",
    975=>"000100011",
    976=>"000110011",
    977=>"111001100",
    978=>"111101000",
    979=>"001000111",
    980=>"000011001",
    981=>"100111000",
    982=>"001000111",
    983=>"111001100",
    984=>"111001100",
    985=>"001000111",
    986=>"001000111",
    987=>"000111011",
    988=>"100000111",
    989=>"000111001",
    990=>"000001001",
    991=>"110001111",
    992=>"011001111",
    993=>"000100010",
    994=>"110110001",
    995=>"001100110",
    996=>"000000000",
    997=>"011001110",
    998=>"000000011",
    999=>"000001111",
    1000=>"111011111",
    1001=>"100000000",
    1002=>"111001001",
    1003=>"000000000",
    1004=>"111111010",
    1005=>"011111110",
    1006=>"010001001",
    1007=>"100110110",
    1008=>"010010010",
    1009=>"000001110",
    1010=>"011001011",
    1011=>"000011010",
    1012=>"111111111",
    1013=>"111111000",
    1014=>"100100111",
    1015=>"111111001",
    1016=>"110000001",
    1017=>"101110110",
    1018=>"110100111",
    1019=>"011101011",
    1020=>"001011100",
    1021=>"011000011",
    1022=>"101110011",
    1023=>"111111011",
    1024=>"111101100",
    1025=>"101101000",
    1026=>"100011111",
    1027=>"011111110",
    1028=>"111100000",
    1029=>"001111101",
    1030=>"011111100",
    1031=>"111100000",
    1032=>"111100000",
    1033=>"110111000",
    1034=>"110100001",
    1035=>"110100101",
    1036=>"100000000",
    1037=>"111111010",
    1038=>"000011111",
    1039=>"011101101",
    1040=>"000000000",
    1041=>"011011011",
    1042=>"100000011",
    1043=>"111111111",
    1044=>"100111111",
    1045=>"100100111",
    1046=>"111110111",
    1047=>"111010100",
    1048=>"110111010",
    1049=>"011011000",
    1050=>"110111111",
    1051=>"001000100",
    1052=>"111011000",
    1053=>"100101101",
    1054=>"001110010",
    1055=>"110100000",
    1056=>"011001101",
    1057=>"011100100",
    1058=>"011011001",
    1059=>"000000100",
    1060=>"110011111",
    1061=>"011011000",
    1062=>"110111011",
    1063=>"011101000",
    1064=>"111001000",
    1065=>"111111000",
    1066=>"111111011",
    1067=>"011001000",
    1068=>"001000000",
    1069=>"001100110",
    1070=>"111111111",
    1071=>"011001000",
    1072=>"110000110",
    1073=>"110111110",
    1074=>"001100110",
    1075=>"001000000",
    1076=>"000000001",
    1077=>"110111111",
    1078=>"011000101",
    1079=>"001100111",
    1080=>"111111111",
    1081=>"000000000",
    1082=>"000000100",
    1083=>"011000100",
    1084=>"001000010",
    1085=>"011000110",
    1086=>"010000010",
    1087=>"011011000",
    1088=>"011001010",
    1089=>"111100110",
    1090=>"101001000",
    1091=>"100111000",
    1092=>"000110111",
    1093=>"011000111",
    1094=>"111011100",
    1095=>"000110111",
    1096=>"011000110",
    1097=>"110010110",
    1098=>"000011000",
    1099=>"000100111",
    1100=>"000100000",
    1101=>"100000110",
    1102=>"111000000",
    1103=>"000100111",
    1104=>"010111111",
    1105=>"111001000",
    1106=>"101111011",
    1107=>"000111001",
    1108=>"000111001",
    1109=>"000010110",
    1110=>"110011000",
    1111=>"111011000",
    1112=>"111011100",
    1113=>"000100001",
    1114=>"111011000",
    1115=>"010100111",
    1116=>"111010000",
    1117=>"010110001",
    1118=>"111101010",
    1119=>"001110010",
    1120=>"000111111",
    1121=>"101000001",
    1122=>"011111100",
    1123=>"100110001",
    1124=>"000011010",
    1125=>"100110110",
    1126=>"111001111",
    1127=>"110010000",
    1128=>"001111111",
    1129=>"110110010",
    1130=>"001001100",
    1131=>"000110110",
    1132=>"010111111",
    1133=>"111011011",
    1134=>"100110010",
    1135=>"110100111",
    1136=>"000010010",
    1137=>"111100111",
    1138=>"010011111",
    1139=>"100111011",
    1140=>"110111000",
    1141=>"010111011",
    1142=>"111111111",
    1143=>"000111111",
    1144=>"011000100",
    1145=>"110111111",
    1146=>"100100000",
    1147=>"110010001",
    1148=>"100110010",
    1149=>"111111001",
    1150=>"100010111",
    1151=>"000110010",
    1152=>"010000100",
    1153=>"001001101",
    1154=>"010100101",
    1155=>"001000110",
    1156=>"101011110",
    1157=>"011000100",
    1158=>"100011011",
    1159=>"001100100",
    1160=>"111011100",
    1161=>"001000100",
    1162=>"001110000",
    1163=>"011000000",
    1164=>"100000000",
    1165=>"001100110",
    1166=>"010001011",
    1167=>"110011101",
    1168=>"011000100",
    1169=>"100011001",
    1170=>"001100110",
    1171=>"000100011",
    1172=>"011000100",
    1173=>"011100110",
    1174=>"000000011",
    1175=>"101110010",
    1176=>"010010101",
    1177=>"101110010",
    1178=>"000001001",
    1179=>"011001110",
    1180=>"011000101",
    1181=>"100101011",
    1182=>"010000100",
    1183=>"111110101",
    1184=>"000000111",
    1185=>"001001001",
    1186=>"000000000",
    1187=>"110011011",
    1188=>"001000000",
    1189=>"110110000",
    1190=>"010100101",
    1191=>"100100100",
    1192=>"000000000",
    1193=>"100100111",
    1194=>"000000000",
    1195=>"001000000",
    1196=>"001001001",
    1197=>"111111111",
    1198=>"110011011",
    1199=>"111111011",
    1200=>"011101101",
    1201=>"110010011",
    1202=>"101101110",
    1203=>"000000000",
    1204=>"001000100",
    1205=>"000000000",
    1206=>"001001101",
    1207=>"110110111",
    1208=>"000000000",
    1209=>"110111111",
    1210=>"000100100",
    1211=>"011001111",
    1212=>"110001111",
    1213=>"001001101",
    1214=>"110111110",
    1215=>"111111111",
    1216=>"110100101",
    1217=>"110000000",
    1218=>"100001011",
    1219=>"000100110",
    1220=>"111011110",
    1221=>"111100001",
    1222=>"001111110",
    1223=>"111001010",
    1224=>"110000000",
    1225=>"111000000",
    1226=>"100000011",
    1227=>"110100000",
    1228=>"010000001",
    1229=>"111111110",
    1230=>"100000001",
    1231=>"001000000",
    1232=>"111000110",
    1233=>"011111000",
    1234=>"110100010",
    1235=>"000000000",
    1236=>"000001011",
    1237=>"011111010",
    1238=>"110100100",
    1239=>"000000101",
    1240=>"001001010",
    1241=>"010111111",
    1242=>"101111111",
    1243=>"111110100",
    1244=>"111111011",
    1245=>"100000011",
    1246=>"100001001",
    1247=>"111001001",
    1248=>"110010011",
    1249=>"001001101",
    1250=>"100100110",
    1251=>"010010000",
    1252=>"100110011",
    1253=>"010011001",
    1254=>"100110110",
    1255=>"010011011",
    1256=>"101110110",
    1257=>"010011011",
    1258=>"100110111",
    1259=>"000001001",
    1260=>"000000100",
    1261=>"011001001",
    1262=>"110011001",
    1263=>"111011001",
    1264=>"101100110",
    1265=>"010010001",
    1266=>"100101111",
    1267=>"001101100",
    1268=>"100110011",
    1269=>"110010001",
    1270=>"000100110",
    1271=>"000100100",
    1272=>"100100111",
    1273=>"011001100",
    1274=>"001100110",
    1275=>"010001000",
    1276=>"001010010",
    1277=>"101110110",
    1278=>"010010001",
    1279=>"000000001",
    1280=>"100100111",
    1281=>"010010011",
    1282=>"011001101",
    1283=>"010010011",
    1284=>"100100110",
    1285=>"100010110",
    1286=>"111101111",
    1287=>"110010010",
    1288=>"111011000",
    1289=>"100100101",
    1290=>"001000100",
    1291=>"010010110",
    1292=>"010000000",
    1293=>"100000001",
    1294=>"001001001",
    1295=>"101001001",
    1296=>"001001001",
    1297=>"000100110",
    1298=>"101001101",
    1299=>"011001001",
    1300=>"010010110",
    1301=>"000010010",
    1302=>"101101001",
    1303=>"001011010",
    1304=>"010010000",
    1305=>"100100100",
    1306=>"110110110",
    1307=>"110100101",
    1308=>"100100100",
    1309=>"101101101",
    1310=>"010101010",
    1311=>"001000001",
    1312=>"100000000",
    1313=>"100110100",
    1314=>"101111101",
    1315=>"111111111",
    1316=>"001101101",
    1317=>"000000000",
    1318=>"000001111",
    1319=>"000101000",
    1320=>"011101110",
    1321=>"000101000",
    1322=>"111111111",
    1323=>"000001100",
    1324=>"111111111",
    1325=>"110111101",
    1326=>"000100001",
    1327=>"000000100",
    1328=>"111111111",
    1329=>"111101100",
    1330=>"100111100",
    1331=>"110000000",
    1332=>"110101110",
    1333=>"000000000",
    1334=>"101100000",
    1335=>"011000000",
    1336=>"111111110",
    1337=>"000001000",
    1338=>"100001110",
    1339=>"101111111",
    1340=>"111011111",
    1341=>"000111001",
    1342=>"111011111",
    1343=>"110111110",
    1344=>"100101100",
    1345=>"111001001",
    1346=>"011000110",
    1347=>"110010111",
    1348=>"000010110",
    1349=>"000100110",
    1350=>"100100111",
    1351=>"111001001",
    1352=>"110100010",
    1353=>"100100111",
    1354=>"110110111",
    1355=>"000100111",
    1356=>"000100100",
    1357=>"000010011",
    1358=>"001000110",
    1359=>"001000111",
    1360=>"001111101",
    1361=>"101100111",
    1362=>"100110101",
    1363=>"000101001",
    1364=>"000000000",
    1365=>"010000110",
    1366=>"111011000",
    1367=>"110101100",
    1368=>"100001011",
    1369=>"011100100",
    1370=>"000000010",
    1371=>"110111000",
    1372=>"100110101",
    1373=>"000000111",
    1374=>"011001010",
    1375=>"010110100",
    1376=>"011111111",
    1377=>"001000111",
    1378=>"000000001",
    1379=>"111000100",
    1380=>"111111000",
    1381=>"101001101",
    1382=>"111111110",
    1383=>"111000110",
    1384=>"001100000",
    1385=>"000000111",
    1386=>"111100011",
    1387=>"000000100",
    1388=>"111000000",
    1389=>"101111111",
    1390=>"100100000",
    1391=>"111001101",
    1392=>"111111010",
    1393=>"000000001",
    1394=>"000100000",
    1395=>"111111011",
    1396=>"111000000",
    1397=>"111000000",
    1398=>"011111111",
    1399=>"110100100",
    1400=>"101101111",
    1401=>"000101000",
    1402=>"000000000",
    1403=>"001111011",
    1404=>"000001101",
    1405=>"111111000",
    1406=>"000011011",
    1407=>"100000000",
    1408=>"011011000",
    1409=>"010011001",
    1410=>"011000000",
    1411=>"100100110",
    1412=>"011011001",
    1413=>"100010110",
    1414=>"011011101",
    1415=>"001111000",
    1416=>"100011011",
    1417=>"100101010",
    1418=>"011001000",
    1419=>"100010000",
    1420=>"000000011",
    1421=>"100100100",
    1422=>"100100110",
    1423=>"101101101",
    1424=>"011011011",
    1425=>"100100110",
    1426=>"000011001",
    1427=>"101101101",
    1428=>"000001100",
    1429=>"001011011",
    1430=>"011011001",
    1431=>"000100010",
    1432=>"000101100",
    1433=>"100000110",
    1434=>"111001100",
    1435=>"000000011",
    1436=>"101100100",
    1437=>"011011001",
    1438=>"100100100",
    1439=>"110100110",
    1440=>"100100000",
    1441=>"001001111",
    1442=>"110110100",
    1443=>"111100001",
    1444=>"000000101",
    1445=>"001001011",
    1446=>"000001111",
    1447=>"110100000",
    1448=>"001111111",
    1449=>"111110100",
    1450=>"000001110",
    1451=>"110100000",
    1452=>"111010000",
    1453=>"111111101",
    1454=>"100000101",
    1455=>"110000101",
    1456=>"100100001",
    1457=>"111100001",
    1458=>"011010100",
    1459=>"100000001",
    1460=>"000000100",
    1461=>"010110000",
    1462=>"000001011",
    1463=>"101111110",
    1464=>"000001011",
    1465=>"110110000",
    1466=>"011011110",
    1467=>"111111100",
    1468=>"111000000",
    1469=>"000101111",
    1470=>"110010000",
    1471=>"001011010",
    1472=>"010111000",
    1473=>"000011011",
    1474=>"000100000",
    1475=>"000100100",
    1476=>"000100000",
    1477=>"010000111",
    1478=>"010111011",
    1479=>"000011010",
    1480=>"000000000",
    1481=>"001001001",
    1482=>"000000000",
    1483=>"000000100",
    1484=>"000000000",
    1485=>"111111111",
    1486=>"110111011",
    1487=>"001001001",
    1488=>"000000000",
    1489=>"000101111",
    1490=>"000111111",
    1491=>"000000101",
    1492=>"011011011",
    1493=>"001111110",
    1494=>"111111010",
    1495=>"100100111",
    1496=>"111111101",
    1497=>"001111111",
    1498=>"101111101",
    1499=>"000000000",
    1500=>"011111001",
    1501=>"101010000",
    1502=>"000000111",
    1503=>"111111111",
    1504=>"111100000",
    1505=>"001100100",
    1506=>"110110010",
    1507=>"001001111",
    1508=>"010000001",
    1509=>"100111111",
    1510=>"111100100",
    1511=>"111100101",
    1512=>"001001001",
    1513=>"111110100",
    1514=>"011011000",
    1515=>"000000001",
    1516=>"000000011",
    1517=>"001001011",
    1518=>"100101100",
    1519=>"001010111",
    1520=>"000011011",
    1521=>"100110110",
    1522=>"000000001",
    1523=>"011000111",
    1524=>"000011011",
    1525=>"001001011",
    1526=>"111100100",
    1527=>"100100111",
    1528=>"010001100",
    1529=>"000011110",
    1530=>"110110001",
    1531=>"001011010",
    1532=>"100101111",
    1533=>"111001100",
    1534=>"000111111",
    1535=>"000010010",
    1536=>"000000001",
    1537=>"110111000",
    1538=>"100010010",
    1539=>"101011111",
    1540=>"000000001",
    1541=>"000000000",
    1542=>"010111000",
    1543=>"110011000",
    1544=>"111000000",
    1545=>"000000000",
    1546=>"110111011",
    1547=>"000000001",
    1548=>"000000011",
    1549=>"011010101",
    1550=>"011011000",
    1551=>"000011000",
    1552=>"010000000",
    1553=>"000000000",
    1554=>"100111011",
    1555=>"001111111",
    1556=>"010111111",
    1557=>"110011000",
    1558=>"111000000",
    1559=>"100100110",
    1560=>"010010010",
    1561=>"101101110",
    1562=>"110110100",
    1563=>"011000000",
    1564=>"001001001",
    1565=>"011001000",
    1566=>"000111111",
    1567=>"001001111",
    1568=>"000110010",
    1569=>"100000110",
    1570=>"111111111",
    1571=>"001000000",
    1572=>"000000000",
    1573=>"000100110",
    1574=>"111000000",
    1575=>"000110111",
    1576=>"000101010",
    1577=>"111111100",
    1578=>"111001000",
    1579=>"000111111",
    1580=>"000001010",
    1581=>"101111010",
    1582=>"000110110",
    1583=>"010000000",
    1584=>"110010111",
    1585=>"101110000",
    1586=>"000010111",
    1587=>"111111110",
    1588=>"100111111",
    1589=>"000000111",
    1590=>"111100000",
    1591=>"000110000",
    1592=>"101010001",
    1593=>"111110111",
    1594=>"000001001",
    1595=>"011000111",
    1596=>"000110110",
    1597=>"111001101",
    1598=>"101010000",
    1599=>"000110100",
    1600=>"111000000",
    1601=>"100000110",
    1602=>"000000000",
    1603=>"011111011",
    1604=>"100000100",
    1605=>"011001001",
    1606=>"111110000",
    1607=>"000101111",
    1608=>"111110100",
    1609=>"000001111",
    1610=>"000000000",
    1611=>"000100100",
    1612=>"000000100",
    1613=>"011111111",
    1614=>"010111100",
    1615=>"111011100",
    1616=>"100100100",
    1617=>"001001111",
    1618=>"011100000",
    1619=>"010110111",
    1620=>"000000101",
    1621=>"110111110",
    1622=>"011000111",
    1623=>"000100111",
    1624=>"000000001",
    1625=>"111111111",
    1626=>"100100100",
    1627=>"111110110",
    1628=>"001000111",
    1629=>"110110100",
    1630=>"000000111",
    1631=>"001001111",
    1632=>"111001111",
    1633=>"100100111",
    1634=>"110100000",
    1635=>"101111110",
    1636=>"010100100",
    1637=>"001100110",
    1638=>"111110111",
    1639=>"111000001",
    1640=>"101001001",
    1641=>"100011001",
    1642=>"110011001",
    1643=>"001000011",
    1644=>"001000000",
    1645=>"101111000",
    1646=>"001110110",
    1647=>"000010111",
    1648=>"110011110",
    1649=>"100110110",
    1650=>"100001000",
    1651=>"111011000",
    1652=>"000001001",
    1653=>"001000010",
    1654=>"111100100",
    1655=>"010011111",
    1656=>"100111001",
    1657=>"000001110",
    1658=>"110110001",
    1659=>"000100110",
    1660=>"000111000",
    1661=>"111000011",
    1662=>"000000100",
    1663=>"000001001",
    1664=>"000000001",
    1665=>"000010010",
    1666=>"100000011",
    1667=>"011010111",
    1668=>"010001011",
    1669=>"000111010",
    1670=>"100000000",
    1671=>"000000001",
    1672=>"111010000",
    1673=>"000000000",
    1674=>"100001110",
    1675=>"000001001",
    1676=>"010010111",
    1677=>"001100100",
    1678=>"110111111",
    1679=>"000000000",
    1680=>"110111110",
    1681=>"010010000",
    1682=>"110100110",
    1683=>"011001011",
    1684=>"010000000",
    1685=>"010110110",
    1686=>"100000101",
    1687=>"100100010",
    1688=>"110011011",
    1689=>"110110000",
    1690=>"111111111",
    1691=>"001000000",
    1692=>"011011000",
    1693=>"000101001",
    1694=>"000001100",
    1695=>"000010000",
    1696=>"001001101",
    1697=>"001001100",
    1698=>"000000000",
    1699=>"010110111",
    1700=>"001001110",
    1701=>"011011110",
    1702=>"100101101",
    1703=>"011011010",
    1704=>"110001001",
    1705=>"001001011",
    1706=>"001010100",
    1707=>"001011010",
    1708=>"000010000",
    1709=>"100000001",
    1710=>"011011011",
    1711=>"100110100",
    1712=>"011011101",
    1713=>"111110110",
    1714=>"001111001",
    1715=>"010010110",
    1716=>"010010110",
    1717=>"100100000",
    1718=>"101100100",
    1719=>"000000010",
    1720=>"010010010",
    1721=>"100001001",
    1722=>"011010110",
    1723=>"110001001",
    1724=>"111111111",
    1725=>"100101001",
    1726=>"000000010",
    1727=>"000000100",
    1728=>"101101101",
    1729=>"101001101",
    1730=>"000100010",
    1731=>"111011000",
    1732=>"000101110",
    1733=>"100100100",
    1734=>"011011011",
    1735=>"100100100",
    1736=>"110110100",
    1737=>"100101111",
    1738=>"000110110",
    1739=>"100100100",
    1740=>"100100100",
    1741=>"111000000",
    1742=>"011001011",
    1743=>"000100000",
    1744=>"100100100",
    1745=>"011011011",
    1746=>"110110110",
    1747=>"001001011",
    1748=>"000100110",
    1749=>"011110000",
    1750=>"111001101",
    1751=>"111001111",
    1752=>"001111110",
    1753=>"111011000",
    1754=>"001001111",
    1755=>"111110000",
    1756=>"000101001",
    1757=>"110100100",
    1758=>"000110110",
    1759=>"000100000",
    1760=>"000011000",
    1761=>"001010101",
    1762=>"100000011",
    1763=>"111111111",
    1764=>"100001011",
    1765=>"010011010",
    1766=>"001001111",
    1767=>"101100101",
    1768=>"101111111",
    1769=>"110111111",
    1770=>"000000000",
    1771=>"110100000",
    1772=>"000000000",
    1773=>"000000000",
    1774=>"111111111",
    1775=>"000100110",
    1776=>"000000000",
    1777=>"110111000",
    1778=>"000000000",
    1779=>"111111111",
    1780=>"101111100",
    1781=>"111111111",
    1782=>"011111000",
    1783=>"000100000",
    1784=>"000000000",
    1785=>"111111111",
    1786=>"111110111",
    1787=>"010000000",
    1788=>"110011000",
    1789=>"000000010",
    1790=>"110101000",
    1791=>"111110001",
    1792=>"111110000",
    1793=>"000000111",
    1794=>"000000111",
    1795=>"101011001",
    1796=>"000111111",
    1797=>"000000111",
    1798=>"111011000",
    1799=>"111100000",
    1800=>"001100000",
    1801=>"111011000",
    1802=>"001001000",
    1803=>"110000001",
    1804=>"000000100",
    1805=>"001111101",
    1806=>"011011011",
    1807=>"000110111",
    1808=>"000111101",
    1809=>"100000111",
    1810=>"001000100",
    1811=>"011111111",
    1812=>"001010111",
    1813=>"100000111",
    1814=>"110100000",
    1815=>"000010100",
    1816=>"111011100",
    1817=>"110110001",
    1818=>"111000101",
    1819=>"000110000",
    1820=>"000000110",
    1821=>"101111100",
    1822=>"000111000",
    1823=>"000011011",
    1824=>"000110111",
    1825=>"110100100",
    1826=>"110011010",
    1827=>"101110111",
    1828=>"000001010",
    1829=>"000001011",
    1830=>"111011100",
    1831=>"100100110",
    1832=>"100001000",
    1833=>"000001011",
    1834=>"011111011",
    1835=>"011001001",
    1836=>"001001001",
    1837=>"010110010",
    1838=>"001100001",
    1839=>"011111001",
    1840=>"111101100",
    1841=>"010100010",
    1842=>"101000110",
    1843=>"000001011",
    1844=>"100000100",
    1845=>"000000000",
    1846=>"000110110",
    1847=>"010000001",
    1848=>"011010011",
    1849=>"010001000",
    1850=>"001000001",
    1851=>"001111010",
    1852=>"110101000",
    1853=>"001000000",
    1854=>"101011110",
    1855=>"000011111",
    1856=>"111001011",
    1857=>"110100000",
    1858=>"100100000",
    1859=>"001011111",
    1860=>"010110100",
    1861=>"010100100",
    1862=>"001011110",
    1863=>"101101000",
    1864=>"011011000",
    1865=>"110110001",
    1866=>"110100000",
    1867=>"110100000",
    1868=>"010000000",
    1869=>"001001111",
    1870=>"111110110",
    1871=>"001001110",
    1872=>"001001011",
    1873=>"110101101",
    1874=>"000100100",
    1875=>"110110100",
    1876=>"110100000",
    1877=>"001001011",
    1878=>"001011011",
    1879=>"110110101",
    1880=>"110100100",
    1881=>"001011110",
    1882=>"110100000",
    1883=>"011011111",
    1884=>"100001111",
    1885=>"001011011",
    1886=>"000100100",
    1887=>"110100000",
    1888=>"001001001",
    1889=>"110100100",
    1890=>"110110110",
    1891=>"010001001",
    1892=>"100100000",
    1893=>"110100100",
    1894=>"101101111",
    1895=>"011011011",
    1896=>"001101100",
    1897=>"001011011",
    1898=>"001011100",
    1899=>"010110000",
    1900=>"010000000",
    1901=>"101101110",
    1902=>"100000101",
    1903=>"110011111",
    1904=>"110100001",
    1905=>"010100011",
    1906=>"001010010",
    1907=>"001001001",
    1908=>"001011000",
    1909=>"010100001",
    1910=>"100100001",
    1911=>"111011011",
    1912=>"000001000",
    1913=>"110110110",
    1914=>"011011110",
    1915=>"111111111",
    1916=>"110000000",
    1917=>"101101001",
    1918=>"010010100",
    1919=>"100001001",
    1920=>"110011111",
    1921=>"101100110",
    1922=>"111011011",
    1923=>"011100111",
    1924=>"010011001",
    1925=>"000000110",
    1926=>"110111101",
    1927=>"101001000",
    1928=>"010001101",
    1929=>"110001100",
    1930=>"111111001",
    1931=>"101101110",
    1932=>"000000000",
    1933=>"000100100",
    1934=>"111111111",
    1935=>"111011101",
    1936=>"010111001",
    1937=>"011011111",
    1938=>"100001010",
    1939=>"011111100",
    1940=>"001011111",
    1941=>"101100111",
    1942=>"101111111",
    1943=>"000100000",
    1944=>"100000001",
    1945=>"111111110",
    1946=>"111011011",
    1947=>"011000110",
    1948=>"000000000",
    1949=>"110110100",
    1950=>"000000000",
    1951=>"111110001",
    1952=>"010110000",
    1953=>"000110101",
    1954=>"111110110",
    1955=>"000000000",
    1956=>"111111110",
    1957=>"011110100",
    1958=>"100101001",
    1959=>"011110110",
    1960=>"001111110",
    1961=>"011011110",
    1962=>"111111101",
    1963=>"010111100",
    1964=>"001000000",
    1965=>"000000001",
    1966=>"111111111",
    1967=>"000000001",
    1968=>"010111000",
    1969=>"010111111",
    1970=>"000000100",
    1971=>"111110110",
    1972=>"011111110",
    1973=>"000000000",
    1974=>"111111001",
    1975=>"011111111",
    1976=>"111111110",
    1977=>"000000001",
    1978=>"111111111",
    1979=>"000000000",
    1980=>"110110110",
    1981=>"111001000",
    1982=>"010110110",
    1983=>"000110000",
    1984=>"001011101",
    1985=>"000111100",
    1986=>"010010100",
    1987=>"100100001",
    1988=>"101011010",
    1989=>"010010110",
    1990=>"101101111",
    1991=>"011111000",
    1992=>"110100100",
    1993=>"001011110",
    1994=>"000000000",
    1995=>"000010000",
    1996=>"010000000",
    1997=>"100001001",
    1998=>"010110101",
    1999=>"100101001",
    2000=>"110101101",
    2001=>"001001010",
    2002=>"000110010",
    2003=>"110110100",
    2004=>"000101101",
    2005=>"101001011",
    2006=>"001001111",
    2007=>"010100000",
    2008=>"011110100",
    2009=>"101001010",
    2010=>"101001010",
    2011=>"111001011",
    2012=>"000101010",
    2013=>"100101001",
    2014=>"110010100",
    2015=>"011010100",
    2016=>"111000000",
    2017=>"011111010",
    2018=>"001011111",
    2019=>"000000000",
    2020=>"111110000",
    2021=>"000000001",
    2022=>"110110000",
    2023=>"111111000",
    2024=>"100101001",
    2025=>"001000000",
    2026=>"100000000",
    2027=>"111111111",
    2028=>"001001001",
    2029=>"000001001",
    2030=>"111100100",
    2031=>"111001001",
    2032=>"101000110",
    2033=>"011110110",
    2034=>"111101101",
    2035=>"001001000",
    2036=>"000000000",
    2037=>"111111111",
    2038=>"111110000",
    2039=>"000001001",
    2040=>"000100100",
    2041=>"011000001",
    2042=>"011101111",
    2043=>"101101000",
    2044=>"100100110",
    2045=>"111110000",
    2046=>"101011111",
    2047=>"101000010");

BEGIN
    weight <= ROM_content(to_integer(address));
END RTL;