LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L3BNROM IS
    PORT (
        coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); -- Instruction bus
        address : IN unsigned(5 DOWNTO 0));
END L3BNROM;

ARCHITECTURE RTL OF L3BNROM IS

    TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem :=
    (0=>"0000010111001111"&"0011110000110110",
    1=>"0000001010110001"&"0010100110111000",
    2=>"0000010101110001"&"0011001100000001",
    3=>"0011011001110011"&"0010000001001110",
    4=>"0000110011010010"&"0010100011100011",
    5=>"1111111001101011"&"0011000101001100",
    6=>"0000001010111110"&"0010110010111001",
    7=>"0001010010111101"&"0010101101101101",
    8=>"0000111010011001"&"0011100010010001",
    9=>"0010111000001110"&"0011000010011001",
    10=>"0000011110010110"&"0010110101101001",
    11=>"0000111111111001"&"0011100011110100",
    12=>"0011010110100000"&"0110100011001111",
    13=>"0000100001101001"&"0101011111010011",
    14=>"0000010001001100"&"0011101101001000",
    15=>"0000101101100101"&"0010010000000010",
    16=>"1111101111110111"&"0011000110110010",
    17=>"0001111001011000"&"0010101110111111",
    18=>"0000001110010111"&"0011000111001001",
    19=>"0000011011100110"&"0011010100100101",
    20=>"0000100001110101"&"0100000000111100",
    21=>"1111011101101010"&"0001001010100010",
    22=>"1111111010001101"&"0011100000001111",
    23=>"0000110100100100"&"0011010110001000",
    24=>"0000001010101010"&"0010111111001110",
    25=>"0001010010110010"&"0011000001111111",
    26=>"0000101111000001"&"0010101011101010",
    27=>"0001110011010000"&"0100101010110010",
    28=>"0001001000010000"&"0010101011111000",
    29=>"0011011001111011"&"0010100011111100",
    30=>"0000110001111111"&"0010101010110111",
    31=>"0000011100110111"&"0001101111100000",
    32=>"1111100001000000"&"0010101111111111",
    33=>"0001001010011010"&"0010100111101011",
    34=>"0000000110001110"&"0011000011010011",
    35=>"1011001000111101"&"0011110101110010",
    36=>"0000011001000110"&"0011010010110110",
    37=>"0001010011111111"&"0010101100010011",
    38=>"0001011001011010"&"0010110110100010",
    39=>"1111110100010100"&"0010101110101110",
    40=>"0000001110100110"&"0011000011111001",
    41=>"0000100110011001"&"0001100001010101",
    42=>"0001011110001110"&"0100010001111010",
    43=>"0001011011011111"&"0010110100100000",
    44=>"1111111111010000"&"0011001100001110",
    45=>"0000110011101100"&"0011010100001000",
    46=>"0000111100111111"&"0011001101101111",
    47=>"0000010010110101"&"0011100010110000",
    48=>"0010010101000011"&"0001110101000000",
    49=>"0000001101100011"&"0010011000100011",
    50=>"1111111110011010"&"0010111000110110",
    51=>"0000000100100000"&"0011101011011001",
    52=>"0010001001111001"&"0001101001111000",
    53=>"1111100001111101"&"0011011010110000",
    54=>"0000010010100011"&"0100000100100000",
    55=>"1111011110010000"&"0010101101110101",
    56=>"0000001011011010"&"0011010011010101",
    57=>"0010001001111111"&"0100010011001011",
    58=>"0000001100101001"&"0011000101111010",
    59=>"0001000101101101"&"0011011010001010",
    60=>"1111010010001000"&"0010100001101000",
    61=>"1101110011101111"&"0011011101100000",
    62=>"0000101110001010"&"0010111100100001",
    63=>"1111110111100010"&"0001110000101010");
    
BEGIN
    coefs <= ROM_content(to_integer(address));
END RTL;