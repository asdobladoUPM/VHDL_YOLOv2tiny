LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L5BNROM IS
    PORT (
        coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); -- Instruction bus
        address : IN unsigned(7 DOWNTO 0));
END L5BNROM;

ARCHITECTURE RTL OF L5BNROM IS

    TYPE ROM_mem IS ARRAY (0 TO 255) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem :=
    (0=>"1111101000110111"&"0011100010110110",
    1=>"1111000011101010"&"0010110010101001",
    2=>"0001100111101110"&"0010111000001000",
    3=>"1111011111010010"&"0010111101001010",
    4=>"0000000000110010"&"0010110000111000",
    5=>"1101110101000011"&"0011101000010110",
    6=>"1111111110011010"&"0010011110101100",
    7=>"0001010001011010"&"0010111111101100",
    8=>"1110111001011111"&"0010111111000110",
    9=>"1110001111110000"&"0010100111111000",
    10=>"1111000100000000"&"0010011011111100",
    11=>"1101110011101100"&"0011001000010001",
    12=>"0001000101000100"&"0001111111000011",
    13=>"1111000010101000"&"0010101001011110",
    14=>"1111011011110001"&"0011110000101100",
    15=>"1111101101000011"&"0011010010100101",
    16=>"1111010000000110"&"0011001000110111",
    17=>"1111011010000111"&"0010011010110111",
    18=>"1111001011001110"&"0011010011000101",
    19=>"1110111010010000"&"0010101100110010",
    20=>"0001011011000000"&"0010110111101101",
    21=>"1111101001111010"&"0010001100011001",
    22=>"0000001110100110"&"0010100011111000",
    23=>"0000111000010101"&"0010010111101000",
    24=>"1100101100011001"&"0011010011111101",
    25=>"1111101011001011"&"0010110000001011",
    26=>"1110100100111010"&"0011011001001110",
    27=>"1111010100011010"&"0001111111110101",
    28=>"1110001001010100"&"0011100111000011",
    29=>"1111101011111011"&"0010100110110101",
    30=>"1110110011111011"&"0011100010110110",
    31=>"0001100001100101"&"0001111110111001",
    32=>"1110111011011100"&"0010010010011011",
    33=>"1110011011010011"&"0010110001000010",
    34=>"0000001101111001"&"0100011001111010",
    35=>"0000101100100010"&"0010111011110111",
    36=>"0000000100010110"&"0010101110001111",
    37=>"1110100101001101"&"0011100001001111",
    38=>"0001101001100110"&"0010000010011111",
    39=>"1111100011100000"&"0011001101100111",
    40=>"0001111101100111"&"0010011111001110",
    41=>"0000010100010011"&"0010111010111111",
    42=>"1110001011111011"&"0010100000010001",
    43=>"1111000100110100"&"0011001010011110",
    44=>"1111011100010100"&"0011010111001110",
    45=>"0000001001111111"&"0010111001010111",
    46=>"1111000111101001"&"0011010110001001",
    47=>"0000100011011100"&"0010100100000001",
    48=>"1111110101001101"&"0010100011111011",
    49=>"1111101011000111"&"0010101000010111",
    50=>"1111101001010110"&"0011101000100101",
    51=>"1111100101000101"&"0010101100001000",
    52=>"1110101011101000"&"0010100001000011",
    53=>"1111011101010111"&"0010011100110000",
    54=>"0000001110101100"&"0010000111001011",
    55=>"1111101100100100"&"0010001110011010",
    56=>"1111111000111000"&"0010100010010001",
    57=>"1111010001100000"&"0010000000001110",
    58=>"1110100110000001"&"0011000101010110",
    59=>"1111011010011100"&"0010101010110000",
    60=>"1111001000100111"&"0011100111000001",
    61=>"1111000101011011"&"0011001011010100",
    62=>"1010010001101000"&"0010001100111001",
    63=>"1111001010011001"&"0011100100110111",
    64=>"0000100010101011"&"0010110110011011",
    65=>"1110111000110111"&"0011011001011111",
    66=>"1111011100100100"&"0011000010011010",
    67=>"1111000001001010"&"0011101001101010",
    68=>"1111111010001000"&"0010101010010011",
    69=>"1111101010011111"&"0011101111110110",
    70=>"1110001011110011"&"0010111110100110",
    71=>"1110101110011110"&"0100000011011111",
    72=>"1111010100110010"&"0010101110110010",
    73=>"1100001000101100"&"0010111111110011",
    74=>"1111101011101001"&"0011010111010110",
    75=>"1101011111110101"&"0011001111111001",
    76=>"1111011010000111"&"0010011100011100",
    77=>"1111110011100000"&"0010101001011101",
    78=>"0000001000111000"&"0010101101101011",
    79=>"1111001100010000"&"0011010110011100",
    80=>"1111110010000111"&"0010010101100100",
    81=>"0000010011010100"&"0011000101101011",
    82=>"0000110101111100"&"0010101100001111",
    83=>"1111010101011001"&"0010111010111011",
    84=>"1111100001110011"&"0010101101110100",
    85=>"1111010111000011"&"0011000010000101",
    86=>"1111111110010101"&"0010111101010011",
    87=>"0001110010000000"&"0011010110111111",
    88=>"0000001000010101"&"0010111111110010",
    89=>"1111111010101111"&"0010111001110010",
    90=>"1111110001111000"&"0010011110110101",
    91=>"1111001000111101"&"0010110011101001",
    92=>"1111100110110101"&"0001110101001111",
    93=>"1111110111010100"&"0010101111011111",
    94=>"0001111010100011"&"0001110000110111",
    95=>"1110111010011100"&"0011101001000100",
    96=>"1110000001100001"&"0011001011011110",
    97=>"1110010101001101"&"0010111000011110",
    98=>"0000001100001001"&"0010101000111011",
    99=>"1111111001111110"&"0010111011111100",
    100=>"1111001011111110"&"0010101100011101",
    101=>"0000011010011111"&"0011001000001110",
    102=>"1111000101010000"&"0011010110001101",
    103=>"0000000100110100"&"0010010111101111",
    104=>"0000000001110100"&"0010100110110000",
    105=>"1111111101001001"&"0010011110111000",
    106=>"0000011111010101"&"0010100101011101",
    107=>"1111101110000011"&"0010110100001101",
    108=>"0000111010110010"&"0010101111100010",
    109=>"0001011100110100"&"0010000001000110",
    110=>"1111010100101101"&"0010001101000011",
    111=>"1110011010100100"&"0010110111100111",
    112=>"0000001011110000"&"0010110010110011",
    113=>"1111101000010101"&"0010011111001100",
    114=>"0000000101111101"&"0010001000101001",
    115=>"0001100000010011"&"0010101000101010",
    116=>"0000110100000110"&"0010010001000000",
    117=>"1011011010100100"&"0011001110001000",
    118=>"1111000111101100"&"0010111000010011",
    119=>"0000010100011101"&"0010111101000011",
    120=>"1111111000110101"&"0011001000111100",
    121=>"0000011110001010"&"0010011000111010",
    122=>"1111100010001110"&"0010110101010010",
    123=>"1111110101001011"&"0010100001011001",
    124=>"1110101000000101"&"0011100000110011",
    125=>"1111110001101000"&"0011000100110011",
    126=>"0000000101000101"&"0010011100101001",
    127=>"0001100110110001"&"0011000000101110",
    128=>"1111100110110101"&"0011000001010101",
    129=>"0000011110001101"&"0010110100110011",
    130=>"0000010010100110"&"0010011111000000",
    131=>"0000000100001110"&"0011010010001001",
    132=>"1111101100100111"&"0010101000111100",
    133=>"1111111001100111"&"0010101110010100",
    134=>"1110111011001110"&"0011011100110111",
    135=>"1110100100001110"&"0011000010110110",
    136=>"1111111100010011"&"0011000001011011",
    137=>"1111001100110001"&"0010110011110101",
    138=>"1111101011111000"&"0010011101001100",
    139=>"1111010100011100"&"0011010001110011",
    140=>"0000101100000101"&"0010011000001010",
    141=>"1110011110011101"&"0011010111000001",
    142=>"1110111101001110"&"0010101111000110",
    143=>"1010100111110001"&"0011100011101110",
    144=>"0000100110111110"&"0011010110110100",
    145=>"1111101100110101"&"0010101101111001",
    146=>"1111011001111010"&"0010110000101110",
    147=>"1110010001110100"&"0011000110011101",
    148=>"1110110010010110"&"0011011001001000",
    149=>"0000101110011101"&"0010010101010100",
    150=>"0000111110100100"&"0010000111010000",
    151=>"1111101010100111"&"0011000010011000",
    152=>"1111101111010011"&"0010100100010011",
    153=>"0000000010000001"&"0011101100101000",
    154=>"0000110110011001"&"0001110110101101",
    155=>"1111010000000110"&"0010111001101010",
    156=>"1111110111011011"&"0010110011010011",
    157=>"1110100001100000"&"0010110010111000",
    158=>"1111101010010010"&"0010110101100000",
    159=>"1100110111001111"&"0010101011111001",
    160=>"1111011010110011"&"0011110100100000",
    161=>"0000010011001111"&"0010100001111010",
    162=>"0000010001010000"&"0010010101001001",
    163=>"1110011100110010"&"0011111100101000",
    164=>"0000101000101100"&"0010111001011001",
    165=>"0000001011010000"&"0010100110100111",
    166=>"1111110010011011"&"0011100101111000",
    167=>"0000011001111011"&"0010100011001101",
    168=>"1111111001110111"&"0010110001000101",
    169=>"0000001001010000"&"0011010110100011",
    170=>"0000010001111010"&"0010100101000001",
    171=>"1101110001111010"&"0010100010000000",
    172=>"1111101100011010"&"0100011011101000",
    173=>"0000001100010111"&"0011000101011011",
    174=>"0000100111001111"&"0010100101011011",
    175=>"0000111101010100"&"0010010111100111",
    176=>"1110111110100001"&"0100011110011000",
    177=>"1111011111000100"&"0011011100110100",
    178=>"1111001000110111"&"0010100101000100",
    179=>"1111010111111011"&"0011000101110001",
    180=>"0000001011001100"&"0010111010111100",
    181=>"1110101111101001"&"0010111001100001",
    182=>"1110111001001100"&"0011011101111011",
    183=>"0000010110011011"&"0011010111010111",
    184=>"1110111010000001"&"0011010110110011",
    185=>"1111000010110010"&"0011011011110011",
    186=>"1111100000001000"&"0011000100000010",
    187=>"0000011000111101"&"0011000000000001",
    188=>"0000000010010000"&"0011000111100101",
    189=>"0000111010000000"&"0010110111000100",
    190=>"1111101101100010"&"0011101000001100",
    191=>"1111010010010101"&"0010100011001110",
    192=>"1111100000111100"&"0010001010000100",
    193=>"1110010010111101"&"0001111011010010",
    194=>"1111000001000100"&"0011011100000111",
    195=>"1111110010001011"&"0011110001000000",
    196=>"0000110001001110"&"0010101011011000",
    197=>"1110111110001111"&"0011111000011100",
    198=>"0000011111110110"&"0010011011100101",
    199=>"1111111101011010"&"0010111001110100",
    200=>"1110010111111011"&"0100000111001110",
    201=>"0000010101000101"&"0011000011011000",
    202=>"1111111011001100"&"0011010011100010",
    203=>"0000111110010111"&"0010010000001001",
    204=>"1111001100000110"&"0010010010101011",
    205=>"1110100111010000"&"0011011011101101",
    206=>"1110011100111010"&"0010100111111001",
    207=>"1111110001011011"&"0010110011000010",
    208=>"0001001111001001"&"0001111110011100",
    209=>"0000101110111100"&"0010110111101001",
    210=>"0000000010100011"&"0010111010010011",
    211=>"0000011101111011"&"0010100101101000",
    212=>"0000010101100000"&"0010001100100110",
    213=>"1111111001001100"&"0011000111011000",
    214=>"0001001100011101"&"0001110110011010",
    215=>"1111110010011110"&"0011000110100000",
    216=>"0001000110010000"&"0001100001010111",
    217=>"0000010101100001"&"0010011001111110",
    218=>"1110001101000010"&"0100110011101000",
    219=>"1111111111001110"&"0010010000101011",
    220=>"0000011111011111"&"0010101101110110",
    221=>"0000011110010000"&"0011010101100000",
    222=>"1111011111000001"&"0010110011110001",
    223=>"1111111100010001"&"0010101011000000",
    224=>"1111100111011110"&"0010011110001111",
    225=>"0000111111000110"&"0010101010110101",
    226=>"0001011011111010"&"0010010011100111",
    227=>"0000101111010011"&"0011001010011011",
    228=>"1101111101000110"&"0010100000001001",
    229=>"0000111110000100"&"0010001111101100",
    230=>"1111110111101100"&"0010010001111101",
    231=>"0000000001111110"&"0010100100110111",
    232=>"1111010000011101"&"0010110001111000",
    233=>"1111101101101110"&"0011001101111011",
    234=>"1111100001001001"&"0010011101001000",
    235=>"0000001000010110"&"0011001101000111",
    236=>"0001001111001010"&"0010001010011001",
    237=>"0000001111101111"&"0011001010010110",
    238=>"0000011010001011"&"0010111100111110",
    239=>"1101110000111011"&"0011001100111101",
    240=>"0000010010100110"&"0010000100100100",
    241=>"1111000010110110"&"0011101001010011",
    242=>"0000011000110110"&"0010110110111001",
    243=>"1111110100110000"&"0010011011011011",
    244=>"1111101010011110"&"0011000110100011",
    245=>"0001011111100101"&"0010010000001111",
    246=>"1101001101110011"&"0011001100111111",
    247=>"1110100001100101"&"0010110011001011",
    248=>"0000101001101011"&"0001111000011101",
    249=>"1111110010101110"&"0010101100011100",
    250=>"0000000010011100"&"0001111000110100",
    251=>"0000100110101001"&"0011000110111010",
    252=>"1111110010001100"&"0010000001101110",
    253=>"1111101110100000"&"0010000111011111",
    254=>"1111101011111110"&"0010111101101011",
    255=>"1111000000111000"&"0010011100011010");
    
BEGIN
    coefs <= ROM_content(to_integer(address));
END RTL;