LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L6WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(6) DOWNTO 0));
END L6WROM;

ARCHITECTURE RTL OF L6WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 131071) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"101100101",
1=>"110100011",
2=>"000100101",
3=>"111011011",
4=>"110110100",
5=>"000000111",
6=>"111100111",
7=>"011111101",
8=>"101101011",
9=>"100100000",
10=>"000010110",
11=>"110101011",
12=>"110111011",
13=>"000010011",
14=>"000100000",
15=>"011100111",
16=>"111100100",
17=>"110000010",
18=>"000111010",
19=>"000001011",
20=>"000110000",
21=>"111100111",
22=>"110100000",
23=>"010111111",
24=>"100000100",
25=>"011010001",
26=>"000010000",
27=>"000010011",
28=>"110100100",
29=>"101000010",
30=>"111100001",
31=>"111111000",
32=>"101100000",
33=>"100100100",
34=>"110011011",
35=>"111100111",
36=>"110100110",
37=>"111100111",
38=>"111100100",
39=>"011100000",
40=>"101111010",
41=>"110000000",
42=>"001101111",
43=>"110101111",
44=>"000111001",
45=>"011100111",
46=>"100110111",
47=>"110011010",
48=>"110000000",
49=>"111111111",
50=>"001111111",
51=>"000110000",
52=>"000111100",
53=>"100011011",
54=>"110100100",
55=>"101100100",
56=>"111111000",
57=>"111100101",
58=>"001010010",
59=>"100100010",
60=>"110010000",
61=>"011111010",
62=>"000000001",
63=>"101101100",
64=>"100110111",
65=>"110100001",
66=>"100110001",
67=>"011001000",
68=>"111000011",
69=>"110000000",
70=>"100100101",
71=>"011111000",
72=>"101100010",
73=>"010011011",
74=>"000011000",
75=>"101011000",
76=>"111100100",
77=>"001101000",
78=>"101101100",
79=>"001001101",
80=>"001011101",
81=>"011110111",
82=>"111000000",
83=>"000000000",
84=>"000100001",
85=>"001100000",
86=>"000110111",
87=>"001001101",
88=>"100010010",
89=>"100111101",
90=>"000000000",
91=>"000000000",
92=>"000111000",
93=>"100101100",
94=>"111111100",
95=>"111110101",
96=>"010110000",
97=>"101000111",
98=>"111100111",
99=>"010110110",
100=>"010010111",
101=>"000011000",
102=>"011011010",
103=>"101100110",
104=>"100110111",
105=>"111111011",
106=>"000100100",
107=>"111011100",
108=>"101100111",
109=>"011011000",
110=>"110100100",
111=>"010010011",
112=>"100111011",
113=>"100111011",
114=>"001100110",
115=>"000000000",
116=>"111100100",
117=>"000100000",
118=>"000001011",
119=>"011000011",
120=>"101011111",
121=>"000000001",
122=>"010010011",
123=>"011111000",
124=>"100100101",
125=>"010010011",
126=>"101100100",
127=>"000010101",
128=>"000101100",
129=>"111100000",
130=>"010111100",
131=>"100001001",
132=>"111101101",
133=>"110001000",
134=>"001001000",
135=>"100100000",
136=>"100111111",
137=>"000000000",
138=>"011010011",
139=>"011001100",
140=>"100111111",
141=>"000011011",
142=>"101101011",
143=>"000001001",
144=>"110111110",
145=>"111100100",
146=>"000001110",
147=>"111100001",
148=>"000011000",
149=>"100100100",
150=>"001011111",
151=>"010010110",
152=>"011011010",
153=>"101011011",
154=>"100100101",
155=>"100100011",
156=>"000000001",
157=>"111111111",
158=>"011111111",
159=>"000000110",
160=>"100100000",
161=>"110100111",
162=>"011011011",
163=>"000011000",
164=>"000011011",
165=>"010011010",
166=>"110101011",
167=>"000000011",
168=>"010000111",
169=>"100111011",
170=>"101100101",
171=>"010100111",
172=>"111000001",
173=>"000000000",
174=>"010010111",
175=>"000000000",
176=>"101000001",
177=>"001011110",
178=>"110000100",
179=>"000000000",
180=>"101000000",
181=>"111011111",
182=>"111001100",
183=>"100110111",
184=>"100001000",
185=>"011011011",
186=>"000010110",
187=>"001011110",
188=>"111011010",
189=>"011001000",
190=>"011001001",
191=>"000000000",
192=>"100000100",
193=>"011011011",
194=>"011011100",
195=>"001011011",
196=>"011011000",
197=>"100100000",
198=>"111000010",
199=>"011011111",
200=>"100111111",
201=>"000011000",
202=>"100001101",
203=>"100100100",
204=>"111100100",
205=>"101111111",
206=>"000100100",
207=>"100100011",
208=>"110000000",
209=>"101101111",
210=>"111100011",
211=>"010100111",
212=>"011100000",
213=>"010001101",
214=>"111010000",
215=>"011011000",
216=>"000011011",
217=>"011000100",
218=>"001001001",
219=>"000000011",
220=>"001101111",
221=>"100110100",
222=>"110011111",
223=>"111100111",
224=>"000011111",
225=>"000000001",
226=>"111001100",
227=>"100110000",
228=>"100000100",
229=>"111011001",
230=>"111111000",
231=>"000000001",
232=>"010000101",
233=>"100000011",
234=>"100001111",
235=>"111111111",
236=>"100100000",
237=>"100100000",
238=>"010110000",
239=>"001100101",
240=>"110100010",
241=>"110000100",
242=>"000000000",
243=>"010111010",
244=>"010110111",
245=>"000000000",
246=>"000000000",
247=>"111100100",
248=>"011100111",
249=>"011000000",
250=>"110110011",
251=>"100100101",
252=>"111111111",
253=>"000100100",
254=>"001100100",
255=>"101100000",
256=>"010011100",
257=>"110111111",
258=>"000000111",
259=>"111111101",
260=>"011001001",
261=>"011000111",
262=>"010010000",
263=>"111010111",
264=>"001001101",
265=>"000000111",
266=>"111011000",
267=>"111011000",
268=>"110010000",
269=>"001001000",
270=>"111011000",
271=>"000111111",
272=>"101000000",
273=>"000111011",
274=>"001000111",
275=>"000110001",
276=>"010110100",
277=>"111011011",
278=>"001000000",
279=>"110011100",
280=>"000011000",
281=>"000000010",
282=>"101101100",
283=>"010111111",
284=>"000001000",
285=>"111001000",
286=>"110100111",
287=>"111111000",
288=>"000000100",
289=>"010011100",
290=>"000110000",
291=>"000000000",
292=>"111001000",
293=>"000000000",
294=>"111111110",
295=>"000000111",
296=>"100100111",
297=>"100000000",
298=>"010000000",
299=>"000010000",
300=>"111111000",
301=>"000000000",
302=>"010010100",
303=>"110010100",
304=>"100100100",
305=>"001011000",
306=>"000111111",
307=>"111111010",
308=>"010111000",
309=>"110110011",
310=>"011011000",
311=>"010111011",
312=>"000000111",
313=>"100111011",
314=>"100100000",
315=>"000101000",
316=>"010011000",
317=>"011011111",
318=>"000000000",
319=>"110000001",
320=>"000111111",
321=>"111000101",
322=>"000000111",
323=>"110100111",
324=>"101010010",
325=>"000010011",
326=>"110110000",
327=>"001000101",
328=>"111111110",
329=>"101100000",
330=>"001111000",
331=>"111111000",
332=>"000000000",
333=>"110111111",
334=>"100100110",
335=>"000000011",
336=>"111101000",
337=>"000111111",
338=>"110011111",
339=>"001000010",
340=>"111110000",
341=>"110110010",
342=>"110100000",
343=>"110011101",
344=>"100111011",
345=>"011001000",
346=>"011000000",
347=>"100100000",
348=>"000010000",
349=>"001101000",
350=>"100100111",
351=>"101001001",
352=>"000000000",
353=>"010101111",
354=>"000111111",
355=>"111001000",
356=>"111101001",
357=>"101100010",
358=>"110111000",
359=>"000000001",
360=>"010011000",
361=>"000111111",
362=>"100100111",
363=>"111110100",
364=>"000111111",
365=>"111111011",
366=>"111111000",
367=>"000111010",
368=>"111010000",
369=>"110000110",
370=>"110110000",
371=>"010011000",
372=>"000000000",
373=>"000000111",
374=>"010111000",
375=>"000000111",
376=>"000000000",
377=>"010011010",
378=>"011111111",
379=>"001000111",
380=>"011110110",
381=>"100001011",
382=>"111111100",
383=>"111001001",
384=>"110000011",
385=>"110000010",
386=>"000100100",
387=>"110111111",
388=>"010000111",
389=>"000001010",
390=>"100100000",
391=>"010111011",
392=>"101101000",
393=>"111111000",
394=>"000000001",
395=>"000000111",
396=>"010101100",
397=>"111001000",
398=>"010000011",
399=>"101001010",
400=>"111100000",
401=>"000100000",
402=>"111111000",
403=>"111111110",
404=>"111110010",
405=>"000101111",
406=>"000010111",
407=>"111000000",
408=>"001000100",
409=>"111011000",
410=>"111111111",
411=>"000000111",
412=>"010111001",
413=>"111000000",
414=>"010000000",
415=>"101000111",
416=>"001011110",
417=>"010010011",
418=>"101010110",
419=>"000111111",
420=>"100111111",
421=>"010111110",
422=>"010000001",
423=>"111011000",
424=>"000001111",
425=>"111000000",
426=>"111101111",
427=>"001100100",
428=>"000000111",
429=>"000000010",
430=>"111011001",
431=>"011000101",
432=>"000000111",
433=>"111111111",
434=>"111111000",
435=>"100111000",
436=>"111111000",
437=>"011100000",
438=>"010100110",
439=>"111011000",
440=>"110111000",
441=>"011011011",
442=>"010111100",
443=>"111111100",
444=>"000011010",
445=>"111000001",
446=>"000001111",
447=>"010111000",
448=>"101100100",
449=>"010111000",
450=>"000000000",
451=>"111111100",
452=>"000000000",
453=>"110100000",
454=>"001011111",
455=>"111111110",
456=>"101000111",
457=>"000001001",
458=>"000010110",
459=>"111111011",
460=>"111100000",
461=>"010011001",
462=>"111000000",
463=>"010010111",
464=>"111000000",
465=>"010001000",
466=>"010010111",
467=>"000000000",
468=>"000000111",
469=>"111111000",
470=>"100000100",
471=>"010000000",
472=>"000000000",
473=>"011111111",
474=>"100100001",
475=>"000000000",
476=>"010000000",
477=>"111000100",
478=>"111111000",
479=>"101101101",
480=>"000001111",
481=>"111001111",
482=>"000000000",
483=>"111111000",
484=>"001001000",
485=>"111111000",
486=>"011000111",
487=>"010110000",
488=>"000000000",
489=>"000000000",
490=>"111111000",
491=>"101101111",
492=>"111011010",
493=>"000100010",
494=>"011011001",
495=>"010101000",
496=>"010000000",
497=>"011001000",
498=>"010111111",
499=>"111000000",
500=>"000001001",
501=>"111001000",
502=>"000101000",
503=>"000101101",
504=>"110111111",
505=>"000010000",
506=>"000111100",
507=>"111101000",
508=>"000000010",
509=>"111010011",
510=>"101101001",
511=>"000000111",
512=>"101000100",
513=>"010000000",
514=>"110110100",
515=>"000111101",
516=>"000101111",
517=>"111111111",
518=>"111011000",
519=>"010111001",
520=>"001000001",
521=>"000110110",
522=>"000000000",
523=>"001000000",
524=>"000000000",
525=>"000000000",
526=>"100000000",
527=>"011001111",
528=>"000000000",
529=>"010111110",
530=>"111100000",
531=>"000000000",
532=>"111101111",
533=>"001101111",
534=>"111011001",
535=>"110111010",
536=>"001001001",
537=>"010111111",
538=>"000000100",
539=>"000010110",
540=>"000010000",
541=>"111000000",
542=>"000001111",
543=>"111011000",
544=>"011111011",
545=>"000000111",
546=>"111001101",
547=>"101101000",
548=>"010000000",
549=>"000001100",
550=>"111001000",
551=>"000111000",
552=>"101111111",
553=>"000000111",
554=>"110000000",
555=>"000111000",
556=>"111111000",
557=>"000101000",
558=>"011010101",
559=>"100000111",
560=>"111000000",
561=>"001000000",
562=>"000000011",
563=>"001111111",
564=>"110000001",
565=>"100001101",
566=>"000000000",
567=>"001000001",
568=>"000001000",
569=>"000101111",
570=>"110111111",
571=>"111001111",
572=>"000000001",
573=>"111111111",
574=>"000000000",
575=>"001001001",
576=>"000010011",
577=>"000000010",
578=>"111111111",
579=>"010000000",
580=>"000000000",
581=>"110000111",
582=>"111111110",
583=>"001100111",
584=>"011111000",
585=>"001000000",
586=>"000100111",
587=>"000000011",
588=>"101100111",
589=>"110000010",
590=>"010000010",
591=>"111001010",
592=>"000011000",
593=>"111111111",
594=>"101000111",
595=>"000100000",
596=>"110010000",
597=>"000000000",
598=>"100100110",
599=>"011000000",
600=>"111001001",
601=>"111100000",
602=>"111110000",
603=>"100101111",
604=>"001000101",
605=>"010100000",
606=>"110111110",
607=>"000000000",
608=>"001001111",
609=>"111111101",
610=>"001101000",
611=>"111111001",
612=>"000000000",
613=>"111111100",
614=>"111000000",
615=>"111010000",
616=>"011001000",
617=>"101111101",
618=>"010111111",
619=>"111111111",
620=>"101000100",
621=>"111111111",
622=>"111000000",
623=>"000111111",
624=>"100000000",
625=>"010000000",
626=>"000000000",
627=>"001000000",
628=>"000111010",
629=>"000000110",
630=>"000111111",
631=>"000000001",
632=>"110111010",
633=>"101111000",
634=>"100000000",
635=>"000001000",
636=>"001001001",
637=>"110010010",
638=>"110110000",
639=>"111010000",
640=>"111111100",
641=>"000111111",
642=>"000111111",
643=>"111111111",
644=>"000000110",
645=>"110110010",
646=>"110100000",
647=>"100100001",
648=>"000001000",
649=>"110001001",
650=>"111101011",
651=>"001011111",
652=>"000111100",
653=>"111111011",
654=>"000000000",
655=>"001000000",
656=>"110100010",
657=>"111111000",
658=>"111111010",
659=>"111101011",
660=>"000100000",
661=>"000111111",
662=>"111101000",
663=>"010010000",
664=>"101000000",
665=>"000100010",
666=>"101000000",
667=>"010111111",
668=>"000000110",
669=>"000000011",
670=>"001101111",
671=>"111000000",
672=>"111111001",
673=>"111111111",
674=>"000000000",
675=>"111100000",
676=>"101000111",
677=>"110001011",
678=>"011000100",
679=>"000100111",
680=>"010101001",
681=>"000001110",
682=>"001100000",
683=>"000000010",
684=>"111111011",
685=>"000000000",
686=>"110100000",
687=>"111111111",
688=>"111111111",
689=>"001100000",
690=>"111011111",
691=>"110000000",
692=>"011000000",
693=>"001000110",
694=>"111100100",
695=>"001111100",
696=>"000000000",
697=>"000001001",
698=>"100100111",
699=>"000101111",
700=>"111010110",
701=>"000111110",
702=>"000000100",
703=>"100000000",
704=>"011111001",
705=>"000110010",
706=>"111011000",
707=>"001001000",
708=>"000000000",
709=>"111000100",
710=>"111111111",
711=>"100111000",
712=>"110001000",
713=>"110111111",
714=>"010000001",
715=>"111111000",
716=>"111011000",
717=>"111000001",
718=>"101000000",
719=>"000111011",
720=>"011110000",
721=>"010000000",
722=>"000000001",
723=>"010111111",
724=>"000010010",
725=>"000111000",
726=>"000000000",
727=>"111101001",
728=>"010000000",
729=>"000000000",
730=>"110111111",
731=>"111111111",
732=>"000000000",
733=>"001111111",
734=>"110000010",
735=>"000001111",
736=>"010111000",
737=>"010110000",
738=>"000110110",
739=>"011111000",
740=>"101010000",
741=>"000101111",
742=>"000000000",
743=>"000111000",
744=>"110110111",
745=>"001000000",
746=>"000000000",
747=>"001010111",
748=>"000000111",
749=>"111111110",
750=>"010110111",
751=>"000000111",
752=>"001000000",
753=>"101101001",
754=>"111111101",
755=>"110010010",
756=>"001001001",
757=>"111111011",
758=>"010010111",
759=>"110111010",
760=>"000111000",
761=>"111111111",
762=>"111111111",
763=>"011000000",
764=>"011000000",
765=>"111000000",
766=>"001000001",
767=>"111011000",
768=>"110011001",
769=>"000000011",
770=>"101000111",
771=>"110101101",
772=>"010111110",
773=>"000000101",
774=>"101000101",
775=>"010000000",
776=>"000000000",
777=>"011010000",
778=>"000111110",
779=>"100011111",
780=>"000000000",
781=>"000111110",
782=>"011011010",
783=>"011110100",
784=>"000010111",
785=>"010110110",
786=>"010001100",
787=>"000111111",
788=>"111100011",
789=>"111000000",
790=>"000000100",
791=>"010010010",
792=>"001000100",
793=>"111111101",
794=>"000000100",
795=>"000100010",
796=>"101001000",
797=>"111000111",
798=>"111110001",
799=>"000000100",
800=>"111001101",
801=>"010010101",
802=>"101101000",
803=>"111000110",
804=>"100100000",
805=>"110110100",
806=>"101000001",
807=>"000110111",
808=>"111000111",
809=>"000001000",
810=>"000111000",
811=>"000000100",
812=>"000011011",
813=>"010111111",
814=>"000101110",
815=>"110110110",
816=>"001000001",
817=>"001101111",
818=>"111000001",
819=>"110000100",
820=>"101111111",
821=>"101111110",
822=>"001011110",
823=>"101000001",
824=>"000001111",
825=>"111001000",
826=>"001000000",
827=>"000000101",
828=>"110100100",
829=>"000111001",
830=>"000000101",
831=>"001001110",
832=>"111111101",
833=>"111111000",
834=>"000100010",
835=>"110000011",
836=>"111111011",
837=>"111111110",
838=>"000000100",
839=>"111011001",
840=>"110010011",
841=>"111111101",
842=>"000001111",
843=>"100000001",
844=>"000000000",
845=>"011001000",
846=>"100100110",
847=>"000011101",
848=>"111111110",
849=>"010000000",
850=>"000000000",
851=>"000101100",
852=>"000000111",
853=>"010111010",
854=>"010100111",
855=>"101111111",
856=>"111100100",
857=>"011101100",
858=>"001001001",
859=>"111111110",
860=>"001000101",
861=>"010001001",
862=>"101000001",
863=>"001000100",
864=>"001000000",
865=>"101000101",
866=>"111111011",
867=>"101100100",
868=>"110110100",
869=>"000111010",
870=>"110111000",
871=>"000000110",
872=>"111111100",
873=>"111110000",
874=>"111000000",
875=>"111000000",
876=>"111001000",
877=>"110110010",
878=>"000010000",
879=>"010001111",
880=>"100100000",
881=>"010000000",
882=>"101110111",
883=>"111001100",
884=>"000101111",
885=>"000000000",
886=>"000111111",
887=>"101101000",
888=>"000100100",
889=>"010011100",
890=>"000000000",
891=>"001101100",
892=>"100110011",
893=>"110100001",
894=>"000000101",
895=>"000010000",
896=>"010010101",
897=>"010101000",
898=>"000000000",
899=>"011011111",
900=>"010111100",
901=>"111000000",
902=>"011011000",
903=>"001010001",
904=>"011001001",
905=>"111000110",
906=>"111000000",
907=>"111111111",
908=>"111001001",
909=>"100000101",
910=>"000000111",
911=>"010000000",
912=>"111100100",
913=>"110100000",
914=>"111110000",
915=>"010000000",
916=>"000111111",
917=>"100100001",
918=>"010111110",
919=>"111100000",
920=>"111111111",
921=>"111111110",
922=>"001111000",
923=>"000000111",
924=>"000000000",
925=>"111111011",
926=>"111100111",
927=>"001101000",
928=>"000101110",
929=>"111101111",
930=>"111001111",
931=>"000010011",
932=>"000001111",
933=>"111011011",
934=>"111001111",
935=>"001111110",
936=>"000000111",
937=>"000010111",
938=>"000000111",
939=>"010111000",
940=>"000000100",
941=>"010010000",
942=>"110100110",
943=>"110000110",
944=>"111001100",
945=>"001011001",
946=>"101101101",
947=>"111101010",
948=>"100100111",
949=>"101101110",
950=>"000010011",
951=>"110110010",
952=>"001111010",
953=>"000110000",
954=>"010010001",
955=>"111110111",
956=>"110010100",
957=>"111111111",
958=>"000110010",
959=>"110111001",
960=>"001000001",
961=>"011000000",
962=>"011011010",
963=>"011011001",
964=>"110111000",
965=>"001111011",
966=>"111000000",
967=>"111111111",
968=>"000111111",
969=>"010000000",
970=>"111110010",
971=>"100000111",
972=>"111100100",
973=>"001011110",
974=>"100000000",
975=>"000000111",
976=>"000010000",
977=>"000000010",
978=>"101010111",
979=>"011111111",
980=>"000000111",
981=>"011100100",
982=>"101000111",
983=>"111000000",
984=>"101001111",
985=>"111000000",
986=>"010001110",
987=>"100100000",
988=>"010101010",
989=>"001000001",
990=>"111010011",
991=>"000001111",
992=>"110000000",
993=>"111000001",
994=>"010000001",
995=>"000001000",
996=>"011000000",
997=>"000000000",
998=>"111111111",
999=>"010000000",
1000=>"000001111",
1001=>"000010111",
1002=>"011111011",
1003=>"111111101",
1004=>"000000000",
1005=>"100000000",
1006=>"000000000",
1007=>"000000000",
1008=>"000010111",
1009=>"100100100",
1010=>"001000111",
1011=>"000011011",
1012=>"010111101",
1013=>"101000000",
1014=>"010000100",
1015=>"110010000",
1016=>"111111000",
1017=>"010111111",
1018=>"111101111",
1019=>"000001010",
1020=>"001001101",
1021=>"000000000",
1022=>"010001101",
1023=>"110000000",
1024=>"011010100",
1025=>"100000110",
1026=>"001000100",
1027=>"000000011",
1028=>"000111110",
1029=>"110010000",
1030=>"110010011",
1031=>"111000100",
1032=>"100101101",
1033=>"000000000",
1034=>"111001100",
1035=>"100100100",
1036=>"011000000",
1037=>"000100001",
1038=>"000101001",
1039=>"011010001",
1040=>"100011011",
1041=>"111100100",
1042=>"000100000",
1043=>"111100100",
1044=>"111001010",
1045=>"111100100",
1046=>"000000110",
1047=>"001000110",
1048=>"100100100",
1049=>"000000011",
1050=>"100100100",
1051=>"100100111",
1052=>"000000001",
1053=>"100100000",
1054=>"111110110",
1055=>"111100101",
1056=>"111011000",
1057=>"100111100",
1058=>"000011001",
1059=>"000011000",
1060=>"000011000",
1061=>"100100110",
1062=>"000000101",
1063=>"100000011",
1064=>"011111101",
1065=>"111011101",
1066=>"011001000",
1067=>"000100100",
1068=>"011011111",
1069=>"011000011",
1070=>"111100111",
1071=>"100000000",
1072=>"000000000",
1073=>"001001011",
1074=>"011110101",
1075=>"100100100",
1076=>"000001000",
1077=>"111011001",
1078=>"000100100",
1079=>"111000010",
1080=>"111010000",
1081=>"111100001",
1082=>"000001000",
1083=>"010000000",
1084=>"011101010",
1085=>"010111000",
1086=>"100100100",
1087=>"110111101",
1088=>"011011000",
1089=>"110100010",
1090=>"011010010",
1091=>"001111111",
1092=>"111110000",
1093=>"111111101",
1094=>"110110000",
1095=>"111100100",
1096=>"000110111",
1097=>"001000000",
1098=>"000100111",
1099=>"011111101",
1100=>"100110000",
1101=>"101100010",
1102=>"000011101",
1103=>"111100110",
1104=>"100000000",
1105=>"011111111",
1106=>"110000011",
1107=>"101000101",
1108=>"101100100",
1109=>"001010110",
1110=>"001001000",
1111=>"001000001",
1112=>"111100100",
1113=>"000000001",
1114=>"001110110",
1115=>"000111011",
1116=>"000100010",
1117=>"000000001",
1118=>"111111111",
1119=>"100111111",
1120=>"010111000",
1121=>"000111111",
1122=>"100100101",
1123=>"000000100",
1124=>"111101100",
1125=>"100100011",
1126=>"011101000",
1127=>"000000000",
1128=>"011011000",
1129=>"000101000",
1130=>"100001100",
1131=>"011100001",
1132=>"011011000",
1133=>"011000111",
1134=>"000010011",
1135=>"101100110",
1136=>"011011011",
1137=>"101001111",
1138=>"000000010",
1139=>"011011000",
1140=>"000011110",
1141=>"100100101",
1142=>"101100010",
1143=>"000000111",
1144=>"011000111",
1145=>"011100011",
1146=>"000011011",
1147=>"110000000",
1148=>"110011100",
1149=>"010000000",
1150=>"000000101",
1151=>"001111011",
1152=>"001011000",
1153=>"110111000",
1154=>"000100000",
1155=>"000100000",
1156=>"110000100",
1157=>"111000000",
1158=>"000001011",
1159=>"100000000",
1160=>"000010111",
1161=>"001000011",
1162=>"001101001",
1163=>"100000000",
1164=>"000100000",
1165=>"000000011",
1166=>"100100010",
1167=>"101000010",
1168=>"100111110",
1169=>"101100101",
1170=>"100100110",
1171=>"101001111",
1172=>"100000010",
1173=>"010000100",
1174=>"100111111",
1175=>"000011011",
1176=>"011111011",
1177=>"101100110",
1178=>"000111111",
1179=>"000000001",
1180=>"000000111",
1181=>"000100000",
1182=>"111011111",
1183=>"000000000",
1184=>"000100100",
1185=>"100000000",
1186=>"000100111",
1187=>"011100010",
1188=>"110100011",
1189=>"101000110",
1190=>"000011011",
1191=>"111100100",
1192=>"111100111",
1193=>"010110100",
1194=>"011111110",
1195=>"100100100",
1196=>"000011000",
1197=>"100100110",
1198=>"100001001",
1199=>"011010110",
1200=>"011011000",
1201=>"100100100",
1202=>"111111111",
1203=>"000000111",
1204=>"011001001",
1205=>"000100000",
1206=>"011011001",
1207=>"101000011",
1208=>"110110001",
1209=>"100000111",
1210=>"011100111",
1211=>"111010101",
1212=>"011011000",
1213=>"010111111",
1214=>"001001011",
1215=>"011000100",
1216=>"101000001",
1217=>"100100000",
1218=>"100100000",
1219=>"001000000",
1220=>"000011000",
1221=>"000110100",
1222=>"111110000",
1223=>"100011011",
1224=>"111100001",
1225=>"111111000",
1226=>"111101110",
1227=>"001101001",
1228=>"111110110",
1229=>"000011001",
1230=>"100001001",
1231=>"011111000",
1232=>"111001000",
1233=>"000110001",
1234=>"100011011",
1235=>"000000001",
1236=>"001111000",
1237=>"111001001",
1238=>"111100111",
1239=>"100111011",
1240=>"011011111",
1241=>"111100000",
1242=>"000100010",
1243=>"000000001",
1244=>"110011001",
1245=>"011000100",
1246=>"111011000",
1247=>"111101110",
1248=>"000100000",
1249=>"100100100",
1250=>"001001001",
1251=>"010100000",
1252=>"000100110",
1253=>"011111000",
1254=>"100100111",
1255=>"000110110",
1256=>"000000000",
1257=>"100011010",
1258=>"111010111",
1259=>"010011011",
1260=>"000111110",
1261=>"011011011",
1262=>"000100000",
1263=>"000000010",
1264=>"001111000",
1265=>"110011110",
1266=>"011011111",
1267=>"100100110",
1268=>"001111111",
1269=>"000000011",
1270=>"000000000",
1271=>"111101111",
1272=>"001000010",
1273=>"111011100",
1274=>"010000000",
1275=>"111111111",
1276=>"100100000",
1277=>"011000000",
1278=>"000111011",
1279=>"111100001",
1280=>"101111111",
1281=>"010010000",
1282=>"011000101",
1283=>"000000000",
1284=>"000000000",
1285=>"101101101",
1286=>"111101101",
1287=>"010110001",
1288=>"011110100",
1289=>"111000111",
1290=>"111101101",
1291=>"111000000",
1292=>"000000110",
1293=>"000011111",
1294=>"111010010",
1295=>"111011000",
1296=>"000000000",
1297=>"000101111",
1298=>"001000111",
1299=>"010010000",
1300=>"101101111",
1301=>"100111000",
1302=>"001011010",
1303=>"000000011",
1304=>"101000000",
1305=>"000111111",
1306=>"101101000",
1307=>"010111111",
1308=>"010000000",
1309=>"111110000",
1310=>"000111111",
1311=>"110010000",
1312=>"010010000",
1313=>"101010000",
1314=>"101000111",
1315=>"000000100",
1316=>"000100000",
1317=>"111110000",
1318=>"010110010",
1319=>"111111000",
1320=>"111111010",
1321=>"000001000",
1322=>"000000110",
1323=>"110000000",
1324=>"111000000",
1325=>"010101000",
1326=>"111101101",
1327=>"000010111",
1328=>"101101111",
1329=>"110001101",
1330=>"101101000",
1331=>"101000000",
1332=>"011001100",
1333=>"101101010",
1334=>"011001111",
1335=>"000000000",
1336=>"001000101",
1337=>"101101111",
1338=>"101101000",
1339=>"110100111",
1340=>"000110100",
1341=>"111110011",
1342=>"001100000",
1343=>"001100111",
1344=>"011011100",
1345=>"000100001",
1346=>"000101001",
1347=>"000000001",
1348=>"011000000",
1349=>"000001101",
1350=>"010110000",
1351=>"000001010",
1352=>"011111000",
1353=>"101001001",
1354=>"100101000",
1355=>"101001101",
1356=>"000000000",
1357=>"101000000",
1358=>"000101101",
1359=>"111011110",
1360=>"000010000",
1361=>"111010010",
1362=>"000000000",
1363=>"110001000",
1364=>"000010111",
1365=>"011010000",
1366=>"011011011",
1367=>"101101101",
1368=>"011111111",
1369=>"000001010",
1370=>"100011001",
1371=>"001011000",
1372=>"101101000",
1373=>"011001110",
1374=>"000111111",
1375=>"000000101",
1376=>"000001001",
1377=>"101111000",
1378=>"101000111",
1379=>"001111111",
1380=>"000000101",
1381=>"110011000",
1382=>"011011000",
1383=>"010010000",
1384=>"001101111",
1385=>"101101001",
1386=>"111111101",
1387=>"110111000",
1388=>"111101000",
1389=>"111101101",
1390=>"000000100",
1391=>"010010010",
1392=>"000100000",
1393=>"100101011",
1394=>"111101001",
1395=>"001000000",
1396=>"001101000",
1397=>"000001000",
1398=>"000011110",
1399=>"000000101",
1400=>"000111110",
1401=>"111011010",
1402=>"010100110",
1403=>"111000101",
1404=>"100110110",
1405=>"011110010",
1406=>"111010101",
1407=>"001000100",
1408=>"010100111",
1409=>"111111111",
1410=>"111000101",
1411=>"011010000",
1412=>"001010000",
1413=>"010111101",
1414=>"011110100",
1415=>"000011000",
1416=>"101011010",
1417=>"110101001",
1418=>"000000100",
1419=>"001010011",
1420=>"000110111",
1421=>"111001001",
1422=>"010101111",
1423=>"101000000",
1424=>"011111011",
1425=>"101101010",
1426=>"100000100",
1427=>"101011011",
1428=>"000000000",
1429=>"101100111",
1430=>"111101111",
1431=>"101111011",
1432=>"111000000",
1433=>"010010000",
1434=>"000010010",
1435=>"110000100",
1436=>"101000000",
1437=>"011010110",
1438=>"100100110",
1439=>"111101111",
1440=>"010000100",
1441=>"111110000",
1442=>"011101101",
1443=>"000111011",
1444=>"110110001",
1445=>"000110000",
1446=>"010101011",
1447=>"110001000",
1448=>"011100100",
1449=>"000011111",
1450=>"101101000",
1451=>"000100101",
1452=>"011110111",
1453=>"000000011",
1454=>"011011001",
1455=>"101001001",
1456=>"010100111",
1457=>"001111000",
1458=>"001101101",
1459=>"000011111",
1460=>"111111010",
1461=>"111100101",
1462=>"100111011",
1463=>"011000000",
1464=>"001011111",
1465=>"000010000",
1466=>"010101000",
1467=>"000000110",
1468=>"110110001",
1469=>"111111101",
1470=>"110111111",
1471=>"101100100",
1472=>"110111000",
1473=>"110000001",
1474=>"000101010",
1475=>"100100001",
1476=>"111000100",
1477=>"110001000",
1478=>"110111100",
1479=>"000010111",
1480=>"111100100",
1481=>"010010111",
1482=>"101000101",
1483=>"000110001",
1484=>"000010000",
1485=>"001011111",
1486=>"011010111",
1487=>"111011000",
1488=>"110110101",
1489=>"011000100",
1490=>"000111111",
1491=>"111010100",
1492=>"000110000",
1493=>"101100100",
1494=>"001000101",
1495=>"000111001",
1496=>"110100000",
1497=>"111100100",
1498=>"110001000",
1499=>"101000000",
1500=>"000000000",
1501=>"001000101",
1502=>"101101111",
1503=>"000010000",
1504=>"010011000",
1505=>"000101100",
1506=>"010111000",
1507=>"110111011",
1508=>"000010000",
1509=>"100010111",
1510=>"100000100",
1511=>"010100101",
1512=>"110101000",
1513=>"100000111",
1514=>"111101100",
1515=>"101001111",
1516=>"010010010",
1517=>"111110000",
1518=>"100101010",
1519=>"101101111",
1520=>"011101111",
1521=>"100100000",
1522=>"100000010",
1523=>"111100000",
1524=>"000000110",
1525=>"101000100",
1526=>"000000111",
1527=>"010111110",
1528=>"010111111",
1529=>"101101000",
1530=>"100000110",
1531=>"010001000",
1532=>"000111011",
1533=>"011000101",
1534=>"111100100",
1535=>"010100000",
1536=>"011001000",
1537=>"000010001",
1538=>"000111000",
1539=>"000111111",
1540=>"101101011",
1541=>"110101000",
1542=>"111101011",
1543=>"000001111",
1544=>"111101000",
1545=>"111111111",
1546=>"000000000",
1547=>"101111111",
1548=>"101001111",
1549=>"111110000",
1550=>"000010011",
1551=>"101000000",
1552=>"000000011",
1553=>"000000000",
1554=>"000000111",
1555=>"101111111",
1556=>"000110111",
1557=>"111110100",
1558=>"001000001",
1559=>"001110000",
1560=>"000100111",
1561=>"001010000",
1562=>"000001000",
1563=>"000011111",
1564=>"000110000",
1565=>"001000001",
1566=>"111101000",
1567=>"000101111",
1568=>"000000000",
1569=>"111111111",
1570=>"000000110",
1571=>"111101000",
1572=>"100111010",
1573=>"110111100",
1574=>"010000000",
1575=>"111111111",
1576=>"000111111",
1577=>"100100000",
1578=>"111010000",
1579=>"000000000",
1580=>"111111001",
1581=>"000111111",
1582=>"111000000",
1583=>"000000000",
1584=>"111000000",
1585=>"100110010",
1586=>"000001010",
1587=>"001000000",
1588=>"000000000",
1589=>"110010000",
1590=>"100100100",
1591=>"010110111",
1592=>"111111111",
1593=>"000010111",
1594=>"110100100",
1595=>"000000000",
1596=>"110111111",
1597=>"101111001",
1598=>"111001100",
1599=>"111111111",
1600=>"001000000",
1601=>"110001110",
1602=>"110110110",
1603=>"111111000",
1604=>"111111110",
1605=>"100000010",
1606=>"111111111",
1607=>"111111111",
1608=>"111111111",
1609=>"000000001",
1610=>"011111011",
1611=>"000000000",
1612=>"111111000",
1613=>"111001011",
1614=>"111011110",
1615=>"100010111",
1616=>"000010011",
1617=>"111111110",
1618=>"111000101",
1619=>"011011010",
1620=>"000010000",
1621=>"111110110",
1622=>"111101100",
1623=>"100000111",
1624=>"111110000",
1625=>"100100100",
1626=>"111011010",
1627=>"111100101",
1628=>"010110111",
1629=>"001001001",
1630=>"010111111",
1631=>"111111001",
1632=>"111000000",
1633=>"000001001",
1634=>"111011000",
1635=>"000000100",
1636=>"000101101",
1637=>"001101000",
1638=>"001001001",
1639=>"110010011",
1640=>"011110110",
1641=>"000100000",
1642=>"110110111",
1643=>"111000001",
1644=>"011001000",
1645=>"000000000",
1646=>"110010001",
1647=>"000001101",
1648=>"101001000",
1649=>"010000101",
1650=>"011001000",
1651=>"101001101",
1652=>"000001000",
1653=>"000000000",
1654=>"111111111",
1655=>"111111001",
1656=>"000000000",
1657=>"001100010",
1658=>"000101000",
1659=>"000101100",
1660=>"000110111",
1661=>"110100000",
1662=>"000000000",
1663=>"011000000",
1664=>"101111000",
1665=>"111101000",
1666=>"111111000",
1667=>"001101010",
1668=>"111011100",
1669=>"000011101",
1670=>"111111011",
1671=>"110110011",
1672=>"001101011",
1673=>"000000111",
1674=>"000000000",
1675=>"000000000",
1676=>"111110000",
1677=>"000000111",
1678=>"001111111",
1679=>"101000100",
1680=>"001001001",
1681=>"100110100",
1682=>"111000111",
1683=>"000001000",
1684=>"101010111",
1685=>"100010111",
1686=>"010111011",
1687=>"110101101",
1688=>"111000100",
1689=>"010000111",
1690=>"111111000",
1691=>"000000010",
1692=>"001001001",
1693=>"111110111",
1694=>"111001111",
1695=>"011000010",
1696=>"110111111",
1697=>"000000000",
1698=>"011111000",
1699=>"000111001",
1700=>"010000000",
1701=>"010010010",
1702=>"000000000",
1703=>"010110010",
1704=>"011000011",
1705=>"100100110",
1706=>"111111000",
1707=>"000100100",
1708=>"001101110",
1709=>"111011101",
1710=>"100000000",
1711=>"111111111",
1712=>"101111011",
1713=>"101001001",
1714=>"000000100",
1715=>"001110110",
1716=>"100100010",
1717=>"000000000",
1718=>"110100000",
1719=>"100010010",
1720=>"011111111",
1721=>"110111110",
1722=>"111001001",
1723=>"000000111",
1724=>"000000000",
1725=>"111111101",
1726=>"111101000",
1727=>"000000001",
1728=>"000000000",
1729=>"000000000",
1730=>"110111101",
1731=>"101001000",
1732=>"000111011",
1733=>"000111111",
1734=>"100000011",
1735=>"110110010",
1736=>"111001011",
1737=>"101111100",
1738=>"001101000",
1739=>"101111111",
1740=>"011011110",
1741=>"000011111",
1742=>"000000000",
1743=>"111100110",
1744=>"110111001",
1745=>"011001011",
1746=>"101110111",
1747=>"111011111",
1748=>"110011101",
1749=>"010100101",
1750=>"110111001",
1751=>"111001111",
1752=>"000000000",
1753=>"000001111",
1754=>"001010010",
1755=>"000000000",
1756=>"011000010",
1757=>"000101110",
1758=>"000000010",
1759=>"111111111",
1760=>"001011111",
1761=>"000000000",
1762=>"111111111",
1763=>"000100110",
1764=>"010111111",
1765=>"011110010",
1766=>"111001000",
1767=>"011001000",
1768=>"011011000",
1769=>"010000100",
1770=>"000000000",
1771=>"000000001",
1772=>"101111111",
1773=>"101000000",
1774=>"100111000",
1775=>"111101101",
1776=>"001111000",
1777=>"000111011",
1778=>"001000011",
1779=>"011011010",
1780=>"110110100",
1781=>"000000000",
1782=>"011000001",
1783=>"011001001",
1784=>"111110111",
1785=>"001011000",
1786=>"001101101",
1787=>"001111111",
1788=>"000111111",
1789=>"101000000",
1790=>"100100111",
1791=>"001001011",
1792=>"110001000",
1793=>"010001000",
1794=>"000011011",
1795=>"010111111",
1796=>"111111111",
1797=>"111010111",
1798=>"111011000",
1799=>"000000000",
1800=>"000010000",
1801=>"000010011",
1802=>"110111110",
1803=>"111111011",
1804=>"000000010",
1805=>"000100011",
1806=>"111111100",
1807=>"000001101",
1808=>"000000000",
1809=>"111000000",
1810=>"111111000",
1811=>"111111111",
1812=>"111111010",
1813=>"111000000",
1814=>"111110011",
1815=>"111111110",
1816=>"010000001",
1817=>"111111111",
1818=>"001000010",
1819=>"000000001",
1820=>"100011011",
1821=>"111101101",
1822=>"011010110",
1823=>"000000100",
1824=>"110110111",
1825=>"000000000",
1826=>"001000001",
1827=>"110110111",
1828=>"001001000",
1829=>"111010000",
1830=>"111100111",
1831=>"000000000",
1832=>"111111010",
1833=>"000000010",
1834=>"000001101",
1835=>"101111111",
1836=>"001001001",
1837=>"111111011",
1838=>"000101001",
1839=>"100011000",
1840=>"000000000",
1841=>"011111111",
1842=>"000000111",
1843=>"111000111",
1844=>"000100011",
1845=>"000000000",
1846=>"001101001",
1847=>"111000100",
1848=>"111110010",
1849=>"001100000",
1850=>"001000000",
1851=>"000000010",
1852=>"001000001",
1853=>"111100100",
1854=>"000000110",
1855=>"011110111",
1856=>"110110010",
1857=>"000001100",
1858=>"000001000",
1859=>"110001110",
1860=>"000000000",
1861=>"111000100",
1862=>"000011010",
1863=>"001001111",
1864=>"000000101",
1865=>"000000010",
1866=>"111000100",
1867=>"011000001",
1868=>"100000011",
1869=>"010111101",
1870=>"000001100",
1871=>"000100011",
1872=>"100000100",
1873=>"110000000",
1874=>"000010001",
1875=>"000000000",
1876=>"000001000",
1877=>"000000010",
1878=>"111011011",
1879=>"000001011",
1880=>"111111110",
1881=>"001010000",
1882=>"110101111",
1883=>"000000000",
1884=>"000000001",
1885=>"101100100",
1886=>"000000000",
1887=>"111110010",
1888=>"000000011",
1889=>"000000000",
1890=>"000111001",
1891=>"101111111",
1892=>"101111101",
1893=>"000001000",
1894=>"000011111",
1895=>"000100100",
1896=>"001011011",
1897=>"101000111",
1898=>"111111010",
1899=>"000010111",
1900=>"111111110",
1901=>"111111000",
1902=>"111011001",
1903=>"000000100",
1904=>"100001100",
1905=>"001101000",
1906=>"110111010",
1907=>"000110111",
1908=>"000110000",
1909=>"110010001",
1910=>"111000000",
1911=>"000000000",
1912=>"000000111",
1913=>"000000000",
1914=>"111111111",
1915=>"000011001",
1916=>"111011011",
1917=>"010010010",
1918=>"011110000",
1919=>"000000000",
1920=>"000001000",
1921=>"010110000",
1922=>"111111111",
1923=>"000001111",
1924=>"000000000",
1925=>"101000101",
1926=>"110011111",
1927=>"001010011",
1928=>"011111011",
1929=>"000001010",
1930=>"111111111",
1931=>"111111101",
1932=>"000110111",
1933=>"110001111",
1934=>"101111111",
1935=>"010000011",
1936=>"111010110",
1937=>"000110111",
1938=>"000000000",
1939=>"110110011",
1940=>"111010011",
1941=>"000011000",
1942=>"000000000",
1943=>"000000000",
1944=>"000000000",
1945=>"011011111",
1946=>"000000000",
1947=>"000111011",
1948=>"111111110",
1949=>"000000000",
1950=>"000011101",
1951=>"000000000",
1952=>"001000010",
1953=>"111110111",
1954=>"000000000",
1955=>"011011111",
1956=>"110111001",
1957=>"110010000",
1958=>"000000000",
1959=>"000111011",
1960=>"111010000",
1961=>"000000001",
1962=>"000000000",
1963=>"110000001",
1964=>"111111111",
1965=>"101010000",
1966=>"111111000",
1967=>"001101111",
1968=>"001001100",
1969=>"000000011",
1970=>"100111111",
1971=>"011011111",
1972=>"111111111",
1973=>"000000011",
1974=>"010010000",
1975=>"110011011",
1976=>"000000000",
1977=>"100100111",
1978=>"010000000",
1979=>"000110110",
1980=>"111110100",
1981=>"111111111",
1982=>"111111100",
1983=>"000000000",
1984=>"000010000",
1985=>"000100111",
1986=>"001010010",
1987=>"111111111",
1988=>"000001001",
1989=>"111110100",
1990=>"000000001",
1991=>"000000000",
1992=>"111111001",
1993=>"000000011",
1994=>"000010010",
1995=>"001001101",
1996=>"000111111",
1997=>"110111000",
1998=>"000000000",
1999=>"101111110",
2000=>"100110100",
2001=>"110111110",
2002=>"000000001",
2003=>"010000100",
2004=>"000000000",
2005=>"000000001",
2006=>"000000000",
2007=>"011010100",
2008=>"010110000",
2009=>"000000000",
2010=>"001000100",
2011=>"101111111",
2012=>"000100110",
2013=>"000000000",
2014=>"000000000",
2015=>"000000111",
2016=>"100000011",
2017=>"111111110",
2018=>"000011010",
2019=>"011001111",
2020=>"000000011",
2021=>"111111111",
2022=>"100110101",
2023=>"010110110",
2024=>"111111111",
2025=>"110100111",
2026=>"111111111",
2027=>"000000000",
2028=>"000000000",
2029=>"000000001",
2030=>"111110000",
2031=>"110000000",
2032=>"100000000",
2033=>"001001001",
2034=>"000000000",
2035=>"110111110",
2036=>"000000110",
2037=>"000000000",
2038=>"111110110",
2039=>"000000101",
2040=>"000000000",
2041=>"111100100",
2042=>"111110111",
2043=>"011111101",
2044=>"111111111",
2045=>"000001001",
2046=>"111110100",
2047=>"000000000",
2048=>"001011111",
2049=>"010000000",
2050=>"000100000",
2051=>"001000011",
2052=>"100100111",
2053=>"000111011",
2054=>"000000000",
2055=>"111000000",
2056=>"000000110",
2057=>"000000000",
2058=>"001001000",
2059=>"000000000",
2060=>"000000101",
2061=>"111111111",
2062=>"000100100",
2063=>"011100000",
2064=>"101001000",
2065=>"010000000",
2066=>"010111100",
2067=>"011000000",
2068=>"000000111",
2069=>"000000100",
2070=>"111101000",
2071=>"111111001",
2072=>"000000000",
2073=>"101011111",
2074=>"000000111",
2075=>"111001000",
2076=>"111010010",
2077=>"011001000",
2078=>"000100111",
2079=>"001001110",
2080=>"011000010",
2081=>"111000111",
2082=>"000011111",
2083=>"000000000",
2084=>"000111111",
2085=>"010111110",
2086=>"000000111",
2087=>"111111101",
2088=>"100111111",
2089=>"100000101",
2090=>"111111000",
2091=>"110111010",
2092=>"000000110",
2093=>"110001000",
2094=>"110110111",
2095=>"111111111",
2096=>"000000110",
2097=>"110100110",
2098=>"000000010",
2099=>"111011010",
2100=>"010001000",
2101=>"111001011",
2102=>"110110100",
2103=>"000001000",
2104=>"011110111",
2105=>"101001001",
2106=>"111000000",
2107=>"110000000",
2108=>"000000010",
2109=>"010001011",
2110=>"000000010",
2111=>"111011110",
2112=>"000000010",
2113=>"101111000",
2114=>"000110110",
2115=>"110011011",
2116=>"111000000",
2117=>"001001001",
2118=>"111001001",
2119=>"100110011",
2120=>"010001001",
2121=>"000110111",
2122=>"111001001",
2123=>"111000000",
2124=>"000110111",
2125=>"010100100",
2126=>"011011111",
2127=>"110000000",
2128=>"001000111",
2129=>"110111101",
2130=>"000001001",
2131=>"000000011",
2132=>"001000000",
2133=>"111110100",
2134=>"000011011",
2135=>"111001010",
2136=>"011001011",
2137=>"010100100",
2138=>"111101000",
2139=>"111111100",
2140=>"000110110",
2141=>"000000001",
2142=>"110111111",
2143=>"110100110",
2144=>"000000000",
2145=>"000000100",
2146=>"010111001",
2147=>"111111000",
2148=>"101100110",
2149=>"110101100",
2150=>"100111110",
2151=>"000111110",
2152=>"011111001",
2153=>"111110000",
2154=>"111111001",
2155=>"000100011",
2156=>"000000110",
2157=>"111000000",
2158=>"111000101",
2159=>"101000000",
2160=>"100100011",
2161=>"111011100",
2162=>"011011000",
2163=>"000001000",
2164=>"001111000",
2165=>"000000001",
2166=>"000000000",
2167=>"000111111",
2168=>"101101000",
2169=>"111100000",
2170=>"111011011",
2171=>"000110011",
2172=>"000000000",
2173=>"000000010",
2174=>"110111111",
2175=>"000110110",
2176=>"111001000",
2177=>"001000000",
2178=>"011111111",
2179=>"111010001",
2180=>"101000111",
2181=>"111111011",
2182=>"110111111",
2183=>"000000110",
2184=>"011000111",
2185=>"111000000",
2186=>"010000000",
2187=>"000110111",
2188=>"000010111",
2189=>"001000110",
2190=>"111111110",
2191=>"100000000",
2192=>"111011011",
2193=>"101101111",
2194=>"000100000",
2195=>"011000110",
2196=>"000000110",
2197=>"111001000",
2198=>"110101000",
2199=>"000000001",
2200=>"111001001",
2201=>"010111110",
2202=>"000110110",
2203=>"100001001",
2204=>"111000000",
2205=>"111110110",
2206=>"100110000",
2207=>"001001000",
2208=>"100100011",
2209=>"110001101",
2210=>"000110111",
2211=>"111000001",
2212=>"000000000",
2213=>"000001111",
2214=>"000000110",
2215=>"000110110",
2216=>"111110110",
2217=>"000000000",
2218=>"101001000",
2219=>"000000000",
2220=>"111111010",
2221=>"000010111",
2222=>"011101101",
2223=>"011111011",
2224=>"010110101",
2225=>"000001011",
2226=>"000101000",
2227=>"000011010",
2228=>"000110111",
2229=>"111101000",
2230=>"010111111",
2231=>"101010110",
2232=>"000000010",
2233=>"000000011",
2234=>"001010111",
2235=>"111001001",
2236=>"100111010",
2237=>"000110111",
2238=>"001011001",
2239=>"110001000",
2240=>"000101101",
2241=>"001001000",
2242=>"001001001",
2243=>"000000011",
2244=>"111110111",
2245=>"000000001",
2246=>"110100000",
2247=>"011000000",
2248=>"110001010",
2249=>"111101111",
2250=>"000000011",
2251=>"111001000",
2252=>"100110110",
2253=>"000000011",
2254=>"111101001",
2255=>"111011000",
2256=>"010000001",
2257=>"000000000",
2258=>"111000011",
2259=>"010000000",
2260=>"000000011",
2261=>"001001100",
2262=>"000000100",
2263=>"000001001",
2264=>"111111001",
2265=>"000000000",
2266=>"111001000",
2267=>"010000001",
2268=>"111011011",
2269=>"100001111",
2270=>"111111010",
2271=>"101001100",
2272=>"111000100",
2273=>"011111110",
2274=>"111001001",
2275=>"000000001",
2276=>"000000000",
2277=>"111001001",
2278=>"000000010",
2279=>"001101001",
2280=>"000000010",
2281=>"000001101",
2282=>"100001000",
2283=>"000111111",
2284=>"000000111",
2285=>"110001001",
2286=>"000000100",
2287=>"000000001",
2288=>"000000000",
2289=>"001010011",
2290=>"111001101",
2291=>"111011111",
2292=>"100100111",
2293=>"111100000",
2294=>"000000010",
2295=>"111111110",
2296=>"111111001",
2297=>"110111111",
2298=>"111000000",
2299=>"000000111",
2300=>"111000000",
2301=>"100000110",
2302=>"011001001",
2303=>"111101001",
2304=>"001100111",
2305=>"100000010",
2306=>"000010111",
2307=>"111111000",
2308=>"100100110",
2309=>"110111101",
2310=>"101011000",
2311=>"111101111",
2312=>"101101111",
2313=>"100100101",
2314=>"000111100",
2315=>"111100101",
2316=>"101100000",
2317=>"101000000",
2318=>"000101101",
2319=>"011110000",
2320=>"111101000",
2321=>"010000000",
2322=>"111101000",
2323=>"101111100",
2324=>"000110111",
2325=>"101100111",
2326=>"110011001",
2327=>"000110111",
2328=>"000101100",
2329=>"010000010",
2330=>"111111101",
2331=>"011011110",
2332=>"101001111",
2333=>"111111010",
2334=>"101100111",
2335=>"111000000",
2336=>"101110001",
2337=>"010101111",
2338=>"000011101",
2339=>"000000111",
2340=>"110100001",
2341=>"100100110",
2342=>"000111110",
2343=>"100100101",
2344=>"111101001",
2345=>"011111111",
2346=>"111111110",
2347=>"010000010",
2348=>"110110110",
2349=>"111100111",
2350=>"100011111",
2351=>"000100101",
2352=>"000000100",
2353=>"001000000",
2354=>"000100101",
2355=>"000000000",
2356=>"101011101",
2357=>"101001001",
2358=>"000001100",
2359=>"000001101",
2360=>"111111101",
2361=>"101101100",
2362=>"011111000",
2363=>"000000001",
2364=>"100100101",
2365=>"111111101",
2366=>"001000000",
2367=>"001000100",
2368=>"101101111",
2369=>"110100100",
2370=>"100001000",
2371=>"111101111",
2372=>"011111000",
2373=>"000111001",
2374=>"101111101",
2375=>"111110010",
2376=>"100100111",
2377=>"111010111",
2378=>"111101110",
2379=>"101101000",
2380=>"100101101",
2381=>"111100100",
2382=>"011101000",
2383=>"000000100",
2384=>"000000000",
2385=>"011000000",
2386=>"011111111",
2387=>"001000011",
2388=>"000100101",
2389=>"100101110",
2390=>"111100000",
2391=>"000101111",
2392=>"000000011",
2393=>"011001000",
2394=>"011011011",
2395=>"001001000",
2396=>"001101101",
2397=>"010110000",
2398=>"101101111",
2399=>"111101111",
2400=>"010000110",
2401=>"110111111",
2402=>"100101101",
2403=>"110110110",
2404=>"001001000",
2405=>"011000000",
2406=>"101000011",
2407=>"000000010",
2408=>"010111011",
2409=>"000000101",
2410=>"110111101",
2411=>"100100101",
2412=>"000010110",
2413=>"100101000",
2414=>"100101001",
2415=>"010111111",
2416=>"100100100",
2417=>"000101101",
2418=>"000000001",
2419=>"100101101",
2420=>"000111010",
2421=>"010101110",
2422=>"100100000",
2423=>"001000000",
2424=>"111111111",
2425=>"010010110",
2426=>"111111101",
2427=>"101100101",
2428=>"001000000",
2429=>"000101110",
2430=>"110010010",
2431=>"111000000",
2432=>"111101100",
2433=>"000000011",
2434=>"000100111",
2435=>"111111010",
2436=>"111101111",
2437=>"111010110",
2438=>"001001101",
2439=>"010000001",
2440=>"000000100",
2441=>"011010010",
2442=>"101111011",
2443=>"000100110",
2444=>"001000001",
2445=>"111111000",
2446=>"011101111",
2447=>"110111111",
2448=>"011101000",
2449=>"111000101",
2450=>"000000000",
2451=>"000101001",
2452=>"111101011",
2453=>"101101100",
2454=>"101101001",
2455=>"100100001",
2456=>"111000101",
2457=>"011000001",
2458=>"111111001",
2459=>"111011010",
2460=>"101100000",
2461=>"111101001",
2462=>"101100001",
2463=>"110010010",
2464=>"001101101",
2465=>"101111111",
2466=>"010010010",
2467=>"000101011",
2468=>"011111011",
2469=>"100001100",
2470=>"100000100",
2471=>"000000111",
2472=>"000100000",
2473=>"001010000",
2474=>"000111111",
2475=>"000010111",
2476=>"100011010",
2477=>"010000000",
2478=>"110010110",
2479=>"111000000",
2480=>"111000110",
2481=>"000100000",
2482=>"000101000",
2483=>"010100000",
2484=>"001001111",
2485=>"111010000",
2486=>"100001000",
2487=>"110111100",
2488=>"001001100",
2489=>"101100100",
2490=>"100000000",
2491=>"010110010",
2492=>"000011011",
2493=>"101101111",
2494=>"111101001",
2495=>"000000000",
2496=>"100100001",
2497=>"010000000",
2498=>"101001101",
2499=>"001001101",
2500=>"000100000",
2501=>"100100100",
2502=>"111111011",
2503=>"001001101",
2504=>"111000001",
2505=>"101010010",
2506=>"110010001",
2507=>"100101001",
2508=>"011100100",
2509=>"100000000",
2510=>"010010101",
2511=>"000000001",
2512=>"101101001",
2513=>"011001100",
2514=>"000100011",
2515=>"111111010",
2516=>"101000100",
2517=>"000010110",
2518=>"001111011",
2519=>"000011111",
2520=>"110000000",
2521=>"101100100",
2522=>"101100011",
2523=>"100101100",
2524=>"010010011",
2525=>"101100000",
2526=>"000000000",
2527=>"101101101",
2528=>"000000101",
2529=>"111101001",
2530=>"111100000",
2531=>"111100111",
2532=>"000000000",
2533=>"001101111",
2534=>"111111000",
2535=>"110110010",
2536=>"011101101",
2537=>"011011111",
2538=>"010010000",
2539=>"000010000",
2540=>"000100111",
2541=>"000111111",
2542=>"001101101",
2543=>"000001110",
2544=>"111011110",
2545=>"001001101",
2546=>"101101100",
2547=>"110100100",
2548=>"110001111",
2549=>"010110110",
2550=>"000100100",
2551=>"000010111",
2552=>"000101001",
2553=>"010010011",
2554=>"000111011",
2555=>"111000000",
2556=>"000000111",
2557=>"100111101",
2558=>"000001001",
2559=>"101100000",
2560=>"011001100",
2561=>"000000000",
2562=>"101000111",
2563=>"011110111",
2564=>"100001001",
2565=>"110101111",
2566=>"000000110",
2567=>"001000000",
2568=>"111111101",
2569=>"010000110",
2570=>"100000100",
2571=>"000001000",
2572=>"110111011",
2573=>"111100000",
2574=>"010110100",
2575=>"000000011",
2576=>"101111001",
2577=>"111100111",
2578=>"111101011",
2579=>"000000000",
2580=>"011010100",
2581=>"111110000",
2582=>"100000000",
2583=>"101101110",
2584=>"000000111",
2585=>"000110000",
2586=>"000000001",
2587=>"011000101",
2588=>"111101111",
2589=>"001000010",
2590=>"001011000",
2591=>"111000000",
2592=>"001001001",
2593=>"000010110",
2594=>"011101110",
2595=>"001001111",
2596=>"001001001",
2597=>"001000111",
2598=>"001000000",
2599=>"000010110",
2600=>"111110000",
2601=>"111010001",
2602=>"100101100",
2603=>"110111010",
2604=>"000100111",
2605=>"010111010",
2606=>"111000000",
2607=>"110111111",
2608=>"101001011",
2609=>"101001000",
2610=>"111111111",
2611=>"101000101",
2612=>"001001001",
2613=>"101110101",
2614=>"000000101",
2615=>"010000100",
2616=>"110000000",
2617=>"000000101",
2618=>"000000000",
2619=>"101101100",
2620=>"010000000",
2621=>"000000000",
2622=>"000000001",
2623=>"010000000",
2624=>"111111111",
2625=>"000000000",
2626=>"010010100",
2627=>"111111110",
2628=>"111110000",
2629=>"111110000",
2630=>"000101111",
2631=>"100000000",
2632=>"001110000",
2633=>"111110101",
2634=>"000001111",
2635=>"110000111",
2636=>"000000101",
2637=>"000100100",
2638=>"011011000",
2639=>"000000111",
2640=>"010000000",
2641=>"001001001",
2642=>"000111100",
2643=>"010000010",
2644=>"000000000",
2645=>"100101110",
2646=>"011100010",
2647=>"000110111",
2648=>"100001000",
2649=>"100100101",
2650=>"001000000",
2651=>"001111111",
2652=>"000000000",
2653=>"000000000",
2654=>"111111111",
2655=>"111011011",
2656=>"010000000",
2657=>"110010110",
2658=>"001001001",
2659=>"100000000",
2660=>"010011011",
2661=>"000000100",
2662=>"000000111",
2663=>"111111000",
2664=>"100111111",
2665=>"110010000",
2666=>"000000101",
2667=>"110001101",
2668=>"110110000",
2669=>"001001101",
2670=>"000000111",
2671=>"000000000",
2672=>"110100100",
2673=>"001010010",
2674=>"000100000",
2675=>"110011101",
2676=>"111110000",
2677=>"010001111",
2678=>"111000000",
2679=>"010010000",
2680=>"111000111",
2681=>"000000111",
2682=>"001010000",
2683=>"111111010",
2684=>"100000100",
2685=>"000000000",
2686=>"111111101",
2687=>"011000000",
2688=>"100000000",
2689=>"000000001",
2690=>"001000000",
2691=>"111000111",
2692=>"000000110",
2693=>"111100000",
2694=>"000000100",
2695=>"000001000",
2696=>"001011000",
2697=>"111000000",
2698=>"000000111",
2699=>"010010000",
2700=>"110110000",
2701=>"111001100",
2702=>"011111101",
2703=>"000100101",
2704=>"100100000",
2705=>"000000000",
2706=>"000101101",
2707=>"101000000",
2708=>"000010111",
2709=>"011010010",
2710=>"001101111",
2711=>"111011111",
2712=>"000001000",
2713=>"000000101",
2714=>"011010111",
2715=>"000010010",
2716=>"100100100",
2717=>"010011000",
2718=>"000000111",
2719=>"101001111",
2720=>"101001010",
2721=>"101010101",
2722=>"111111110",
2723=>"000000111",
2724=>"000000000",
2725=>"111000000",
2726=>"111110000",
2727=>"111101101",
2728=>"001000100",
2729=>"010001000",
2730=>"101011111",
2731=>"110000000",
2732=>"111000110",
2733=>"010010001",
2734=>"100000101",
2735=>"111111010",
2736=>"100110111",
2737=>"010110100",
2738=>"000010000",
2739=>"000110111",
2740=>"111011011",
2741=>"111111010",
2742=>"111111111",
2743=>"111111000",
2744=>"101000100",
2745=>"000101111",
2746=>"010101001",
2747=>"000010010",
2748=>"111111111",
2749=>"010110000",
2750=>"111100100",
2751=>"011010001",
2752=>"101000010",
2753=>"010010000",
2754=>"010111000",
2755=>"001000000",
2756=>"000000100",
2757=>"001001100",
2758=>"000011011",
2759=>"000100111",
2760=>"101001100",
2761=>"010000101",
2762=>"111111111",
2763=>"011001000",
2764=>"000010000",
2765=>"000000001",
2766=>"111100100",
2767=>"111101111",
2768=>"000101111",
2769=>"110110100",
2770=>"101111111",
2771=>"000000011",
2772=>"000000000",
2773=>"000110000",
2774=>"000000100",
2775=>"000011000",
2776=>"000101000",
2777=>"100111011",
2778=>"001011001",
2779=>"000000110",
2780=>"011000101",
2781=>"110010011",
2782=>"010100111",
2783=>"111000010",
2784=>"111000101",
2785=>"110010101",
2786=>"000000110",
2787=>"101111111",
2788=>"011110111",
2789=>"010110000",
2790=>"100100000",
2791=>"000011011",
2792=>"111111110",
2793=>"010000111",
2794=>"101000001",
2795=>"110110100",
2796=>"111111101",
2797=>"110000101",
2798=>"000000000",
2799=>"010000000",
2800=>"111001000",
2801=>"100100000",
2802=>"011101111",
2803=>"000100010",
2804=>"110110011",
2805=>"000000100",
2806=>"000000010",
2807=>"001111111",
2808=>"000001111",
2809=>"111110110",
2810=>"101111001",
2811=>"101111011",
2812=>"100111111",
2813=>"111110000",
2814=>"000100000",
2815=>"000001111",
2816=>"101101101",
2817=>"000000001",
2818=>"001001111",
2819=>"101010000",
2820=>"100100111",
2821=>"010010110",
2822=>"001101101",
2823=>"000010101",
2824=>"010010000",
2825=>"011111001",
2826=>"100000001",
2827=>"000011111",
2828=>"001101111",
2829=>"111111000",
2830=>"000000100",
2831=>"101000000",
2832=>"000010000",
2833=>"111010010",
2834=>"011100000",
2835=>"110100000",
2836=>"111111111",
2837=>"000110100",
2838=>"011001000",
2839=>"000011101",
2840=>"010000000",
2841=>"111000000",
2842=>"111000000",
2843=>"011000000",
2844=>"000001111",
2845=>"111001001",
2846=>"010001000",
2847=>"111001000",
2848=>"110110000",
2849=>"010000101",
2850=>"111111111",
2851=>"000111011",
2852=>"110111100",
2853=>"011101101",
2854=>"011000000",
2855=>"001111111",
2856=>"110011001",
2857=>"010001000",
2858=>"000011011",
2859=>"111111010",
2860=>"101100101",
2861=>"010110001",
2862=>"111111011",
2863=>"100010100",
2864=>"010001100",
2865=>"011001111",
2866=>"111111100",
2867=>"000101000",
2868=>"000000101",
2869=>"100001111",
2870=>"001101111",
2871=>"010011000",
2872=>"100010011",
2873=>"000000011",
2874=>"000000000",
2875=>"111111000",
2876=>"000101011",
2877=>"011001001",
2878=>"101111111",
2879=>"011011000",
2880=>"111000000",
2881=>"101111011",
2882=>"000000001",
2883=>"011001001",
2884=>"000001001",
2885=>"010011111",
2886=>"101111000",
2887=>"001111100",
2888=>"001111011",
2889=>"110100000",
2890=>"101000100",
2891=>"110011000",
2892=>"111111000",
2893=>"101100001",
2894=>"110110011",
2895=>"000001011",
2896=>"000101111",
2897=>"111111110",
2898=>"010111001",
2899=>"011001000",
2900=>"101001000",
2901=>"111110101",
2902=>"011011001",
2903=>"001111111",
2904=>"000100111",
2905=>"101111001",
2906=>"011010011",
2907=>"011010001",
2908=>"000000100",
2909=>"000000100",
2910=>"111111000",
2911=>"110000000",
2912=>"000000101",
2913=>"010000001",
2914=>"001000111",
2915=>"111111110",
2916=>"100101011",
2917=>"100010010",
2918=>"110110000",
2919=>"110000000",
2920=>"110000000",
2921=>"000000000",
2922=>"101111101",
2923=>"000001001",
2924=>"111111000",
2925=>"001100110",
2926=>"000000000",
2927=>"001111010",
2928=>"100100000",
2929=>"001000111",
2930=>"001100111",
2931=>"000101111",
2932=>"111010000",
2933=>"000000000",
2934=>"000100111",
2935=>"001100000",
2936=>"000000100",
2937=>"111110010",
2938=>"110110111",
2939=>"111111101",
2940=>"101000000",
2941=>"110000100",
2942=>"110110010",
2943=>"111000000",
2944=>"110101000",
2945=>"101101011",
2946=>"010010000",
2947=>"001111011",
2948=>"110001010",
2949=>"111111000",
2950=>"000011011",
2951=>"001000111",
2952=>"011011000",
2953=>"111101111",
2954=>"000010000",
2955=>"101111110",
2956=>"010000000",
2957=>"100010010",
2958=>"110110000",
2959=>"000001100",
2960=>"011011010",
2961=>"111100111",
2962=>"110000000",
2963=>"101000000",
2964=>"001001100",
2965=>"000000011",
2966=>"000101111",
2967=>"001011000",
2968=>"001001101",
2969=>"010111111",
2970=>"101100101",
2971=>"110000000",
2972=>"000000000",
2973=>"010000000",
2974=>"000110111",
2975=>"000101111",
2976=>"001001011",
2977=>"111111111",
2978=>"101000100",
2979=>"001101001",
2980=>"010000000",
2981=>"100100110",
2982=>"111111001",
2983=>"000000111",
2984=>"001111111",
2985=>"000010001",
2986=>"000000110",
2987=>"100000010",
2988=>"000000011",
2989=>"110111111",
2990=>"100101111",
2991=>"111111010",
2992=>"111011000",
2993=>"000001010",
2994=>"111111101",
2995=>"100000001",
2996=>"110100000",
2997=>"001000100",
2998=>"001111011",
2999=>"000001011",
3000=>"010100111",
3001=>"100001101",
3002=>"001010100",
3003=>"110010100",
3004=>"110101011",
3005=>"111110000",
3006=>"110110001",
3007=>"000000111",
3008=>"000100110",
3009=>"000000000",
3010=>"111111101",
3011=>"100110111",
3012=>"000101100",
3013=>"100010011",
3014=>"001010111",
3015=>"000110000",
3016=>"000111011",
3017=>"000110011",
3018=>"111111101",
3019=>"011000000",
3020=>"011010000",
3021=>"001100000",
3022=>"110111111",
3023=>"111010000",
3024=>"011110000",
3025=>"111110010",
3026=>"101111011",
3027=>"110000000",
3028=>"010000000",
3029=>"000000000",
3030=>"000001111",
3031=>"111011000",
3032=>"000101111",
3033=>"001111100",
3034=>"110110100",
3035=>"001100111",
3036=>"110011001",
3037=>"000111101",
3038=>"000000000",
3039=>"110000001",
3040=>"001101101",
3041=>"001111111",
3042=>"000101111",
3043=>"100111111",
3044=>"000000000",
3045=>"101111000",
3046=>"111000001",
3047=>"010111011",
3048=>"011000001",
3049=>"000000110",
3050=>"001100100",
3051=>"000001010",
3052=>"000000111",
3053=>"010110010",
3054=>"000001011",
3055=>"011011000",
3056=>"110110000",
3057=>"001101100",
3058=>"001111001",
3059=>"110000000",
3060=>"001110010",
3061=>"000000111",
3062=>"000000111",
3063=>"000000000",
3064=>"000110111",
3065=>"001111000",
3066=>"111110000",
3067=>"001000010",
3068=>"000101011",
3069=>"000000000",
3070=>"011111100",
3071=>"101101111",
3072=>"101100100",
3073=>"111011110",
3074=>"100100110",
3075=>"010011000",
3076=>"011110001",
3077=>"011011000",
3078=>"100110111",
3079=>"100100100",
3080=>"011011001",
3081=>"100100000",
3082=>"100100110",
3083=>"000000001",
3084=>"100110111",
3085=>"011001001",
3086=>"110110110",
3087=>"100100100",
3088=>"001010001",
3089=>"100110111",
3090=>"110110110",
3091=>"010000000",
3092=>"110110011",
3093=>"001011000",
3094=>"111001111",
3095=>"000110010",
3096=>"100100111",
3097=>"001000110",
3098=>"011011001",
3099=>"000010110",
3100=>"100111111",
3101=>"110110111",
3102=>"001110110",
3103=>"111011001",
3104=>"011000000",
3105=>"011111100",
3106=>"110111000",
3107=>"011001000",
3108=>"100100010",
3109=>"000011001",
3110=>"011011000",
3111=>"000100100",
3112=>"001000000",
3113=>"011011011",
3114=>"000000110",
3115=>"111100001",
3116=>"011110111",
3117=>"110111111",
3118=>"011111101",
3119=>"000100100",
3120=>"110111000",
3121=>"000000000",
3122=>"111011001",
3123=>"110100100",
3124=>"100100111",
3125=>"000000100",
3126=>"001100110",
3127=>"100100011",
3128=>"011101111",
3129=>"100100111",
3130=>"000000000",
3131=>"110111100",
3132=>"001001000",
3133=>"111111010",
3134=>"100100110",
3135=>"001001000",
3136=>"100000111",
3137=>"000111101",
3138=>"011001001",
3139=>"101101000",
3140=>"011011000",
3141=>"111011000",
3142=>"100110011",
3143=>"000000110",
3144=>"011011011",
3145=>"110000111",
3146=>"100110111",
3147=>"100100111",
3148=>"001011011",
3149=>"110111101",
3150=>"001001010",
3151=>"110111110",
3152=>"100100110",
3153=>"110111000",
3154=>"011100011",
3155=>"000000000",
3156=>"100100100",
3157=>"010100111",
3158=>"001000000",
3159=>"100100111",
3160=>"111111011",
3161=>"011111011",
3162=>"111110110",
3163=>"001101100",
3164=>"000000000",
3165=>"100100000",
3166=>"001101111",
3167=>"000010010",
3168=>"011011000",
3169=>"001011101",
3170=>"100110010",
3171=>"100110011",
3172=>"011001100",
3173=>"110110101",
3174=>"011100110",
3175=>"100100110",
3176=>"011011000",
3177=>"011110100",
3178=>"001110011",
3179=>"011110000",
3180=>"001011100",
3181=>"000000101",
3182=>"000000001",
3183=>"101011011",
3184=>"110101100",
3185=>"000101001",
3186=>"100010011",
3187=>"001000000",
3188=>"011111000",
3189=>"100100011",
3190=>"011001011",
3191=>"101111110",
3192=>"000001011",
3193=>"011011011",
3194=>"110111000",
3195=>"011110011",
3196=>"011001001",
3197=>"011011001",
3198=>"110100100",
3199=>"100010011",
3200=>"011111010",
3201=>"110110010",
3202=>"001000000",
3203=>"011000111",
3204=>"100101000",
3205=>"000100001",
3206=>"101001101",
3207=>"000100100",
3208=>"111010010",
3209=>"100100101",
3210=>"100100100",
3211=>"000100100",
3212=>"011011000",
3213=>"000100111",
3214=>"000110100",
3215=>"100100010",
3216=>"111110000",
3217=>"010111110",
3218=>"000111111",
3219=>"110110000",
3220=>"010011000",
3221=>"101101111",
3222=>"100100111",
3223=>"011001000",
3224=>"001101110",
3225=>"110001000",
3226=>"100110111",
3227=>"000100111",
3228=>"110110000",
3229=>"000100111",
3230=>"000100100",
3231=>"100110111",
3232=>"000011111",
3233=>"100001001",
3234=>"000110110",
3235=>"100101111",
3236=>"011010000",
3237=>"001011010",
3238=>"111001001",
3239=>"011110100",
3240=>"000110111",
3241=>"011001001",
3242=>"011011001",
3243=>"111110110",
3244=>"011000000",
3245=>"001011011",
3246=>"000110110",
3247=>"111010111",
3248=>"111111111",
3249=>"100100000",
3250=>"000111001",
3251=>"000000000",
3252=>"011001010",
3253=>"111001001",
3254=>"011010000",
3255=>"001100100",
3256=>"100100011",
3257=>"111000010",
3258=>"011000000",
3259=>"010001101",
3260=>"010100100",
3261=>"011011011",
3262=>"011011001",
3263=>"110110011",
3264=>"100100111",
3265=>"100110110",
3266=>"000001101",
3267=>"110100110",
3268=>"100100110",
3269=>"110000001",
3270=>"100010010",
3271=>"001001001",
3272=>"101000000",
3273=>"111000000",
3274=>"101100011",
3275=>"111001001",
3276=>"100110111",
3277=>"000000110",
3278=>"100110110",
3279=>"011001001",
3280=>"100100100",
3281=>"111111101",
3282=>"100110011",
3283=>"011011011",
3284=>"000100111",
3285=>"011011001",
3286=>"111110110",
3287=>"100001111",
3288=>"100110111",
3289=>"000000001",
3290=>"111111001",
3291=>"100100111",
3292=>"110110010",
3293=>"011001001",
3294=>"011001001",
3295=>"111111111",
3296=>"000001011",
3297=>"100100111",
3298=>"010100101",
3299=>"011000000",
3300=>"000000000",
3301=>"000110011",
3302=>"001001001",
3303=>"000010111",
3304=>"001000001",
3305=>"011101101",
3306=>"100000011",
3307=>"011011000",
3308=>"001001000",
3309=>"001001001",
3310=>"010111000",
3311=>"000011000",
3312=>"011011000",
3313=>"110110111",
3314=>"001111010",
3315=>"111100111",
3316=>"011011011",
3317=>"110111110",
3318=>"100000000",
3319=>"000001101",
3320=>"100100111",
3321=>"110110000",
3322=>"110110000",
3323=>"110000000",
3324=>"100011111",
3325=>"100100110",
3326=>"000010000",
3327=>"100100111",
3328=>"010100100",
3329=>"000000011",
3330=>"101101001",
3331=>"100110111",
3332=>"000000010",
3333=>"000000010",
3334=>"110000010",
3335=>"000111111",
3336=>"000110110",
3337=>"000010110",
3338=>"010010000",
3339=>"001000000",
3340=>"000000110",
3341=>"000000000",
3342=>"011011101",
3343=>"001110111",
3344=>"000000110",
3345=>"000000000",
3346=>"100001001",
3347=>"110111000",
3348=>"111111110",
3349=>"000000011",
3350=>"111111111",
3351=>"101110100",
3352=>"001010001",
3353=>"000000000",
3354=>"100101101",
3355=>"101101111",
3356=>"101000011",
3357=>"000001111",
3358=>"110000100",
3359=>"000000101",
3360=>"000000000",
3361=>"000101110",
3362=>"000101111",
3363=>"011110111",
3364=>"010110000",
3365=>"111000101",
3366=>"000010000",
3367=>"111000000",
3368=>"001111111",
3369=>"000010111",
3370=>"000000000",
3371=>"111100111",
3372=>"011011000",
3373=>"000110111",
3374=>"110000000",
3375=>"001001111",
3376=>"010001000",
3377=>"001011011",
3378=>"111111111",
3379=>"000100101",
3380=>"110000000",
3381=>"111110000",
3382=>"110000000",
3383=>"000000011",
3384=>"111111111",
3385=>"111000000",
3386=>"000000000",
3387=>"101111111",
3388=>"110111000",
3389=>"111111110",
3390=>"101000001",
3391=>"111100100",
3392=>"001001101",
3393=>"111011111",
3394=>"001111010",
3395=>"011100010",
3396=>"111011000",
3397=>"000000110",
3398=>"110000000",
3399=>"101000000",
3400=>"001001011",
3401=>"111000000",
3402=>"000001010",
3403=>"011110010",
3404=>"010001001",
3405=>"001011000",
3406=>"100110010",
3407=>"110111110",
3408=>"010001001",
3409=>"110001011",
3410=>"010111000",
3411=>"101100000",
3412=>"111000101",
3413=>"000001000",
3414=>"110111100",
3415=>"111000001",
3416=>"001000000",
3417=>"011011010",
3418=>"110111110",
3419=>"011001110",
3420=>"000000011",
3421=>"000001011",
3422=>"111000010",
3423=>"101001011",
3424=>"010111110",
3425=>"100001111",
3426=>"011010000",
3427=>"000001111",
3428=>"100111000",
3429=>"000100110",
3430=>"111001110",
3431=>"010000111",
3432=>"001000000",
3433=>"010000000",
3434=>"111000111",
3435=>"001000000",
3436=>"010001111",
3437=>"111010010",
3438=>"000000011",
3439=>"011011111",
3440=>"111111001",
3441=>"001111111",
3442=>"011000000",
3443=>"000000000",
3444=>"101111111",
3445=>"001101000",
3446=>"100000010",
3447=>"011001111",
3448=>"001000000",
3449=>"101111111",
3450=>"111100000",
3451=>"010010111",
3452=>"100110010",
3453=>"100000100",
3454=>"000100111",
3455=>"000000101",
3456=>"111000111",
3457=>"000000110",
3458=>"110010000",
3459=>"101011111",
3460=>"000000001",
3461=>"111101111",
3462=>"110000111",
3463=>"000011010",
3464=>"011101110",
3465=>"111011111",
3466=>"000000010",
3467=>"011000110",
3468=>"000001111",
3469=>"110100001",
3470=>"101101110",
3471=>"001001110",
3472=>"110100100",
3473=>"111101101",
3474=>"000010000",
3475=>"000001101",
3476=>"111111001",
3477=>"111111001",
3478=>"111110011",
3479=>"000000011",
3480=>"111000000",
3481=>"001111111",
3482=>"111111000",
3483=>"001000011",
3484=>"111111011",
3485=>"111101100",
3486=>"011101101",
3487=>"001001000",
3488=>"101101010",
3489=>"111000101",
3490=>"101001100",
3491=>"000000001",
3492=>"111101000",
3493=>"111001000",
3494=>"100111111",
3495=>"001101000",
3496=>"101101111",
3497=>"000101101",
3498=>"100111111",
3499=>"100111000",
3500=>"000010011",
3501=>"110111101",
3502=>"111111111",
3503=>"010001111",
3504=>"111000000",
3505=>"001100001",
3506=>"101001101",
3507=>"000100111",
3508=>"100110010",
3509=>"000101110",
3510=>"000000000",
3511=>"011010000",
3512=>"001111100",
3513=>"100110011",
3514=>"010110000",
3515=>"111111001",
3516=>"010000010",
3517=>"001000000",
3518=>"100111001",
3519=>"000100001",
3520=>"110000000",
3521=>"000001101",
3522=>"111000000",
3523=>"111110010",
3524=>"111011010",
3525=>"101101010",
3526=>"010000000",
3527=>"000000000",
3528=>"100111110",
3529=>"001001111",
3530=>"000010000",
3531=>"111000101",
3532=>"011001001",
3533=>"011011010",
3534=>"111111111",
3535=>"000101111",
3536=>"111110000",
3537=>"011000110",
3538=>"000010111",
3539=>"000111111",
3540=>"011000000",
3541=>"000000100",
3542=>"111011010",
3543=>"001011111",
3544=>"000111110",
3545=>"100000101",
3546=>"111100000",
3547=>"000000101",
3548=>"101000110",
3549=>"010111111",
3550=>"000101111",
3551=>"000000100",
3552=>"000000101",
3553=>"111110000",
3554=>"000000111",
3555=>"100110111",
3556=>"000000001",
3557=>"000001111",
3558=>"111110000",
3559=>"000101111",
3560=>"110010000",
3561=>"000000000",
3562=>"101001000",
3563=>"001101000",
3564=>"000000110",
3565=>"000000000",
3566=>"000000000",
3567=>"001001011",
3568=>"000111101",
3569=>"101010010",
3570=>"110010000",
3571=>"011101110",
3572=>"010001011",
3573=>"000001011",
3574=>"000010101",
3575=>"000100100",
3576=>"010010000",
3577=>"110001111",
3578=>"101101111",
3579=>"001111111",
3580=>"111010111",
3581=>"100100111",
3582=>"111000010",
3583=>"111000010",
3584=>"010010011",
3585=>"000011001",
3586=>"111001001",
3587=>"011001110",
3588=>"001011111",
3589=>"100100000",
3590=>"111001001",
3591=>"110000110",
3592=>"000000110",
3593=>"000001001",
3594=>"111001000",
3595=>"000110111",
3596=>"000110110",
3597=>"000110110",
3598=>"100100110",
3599=>"101110011",
3600=>"000000100",
3601=>"000001100",
3602=>"110111000",
3603=>"000000000",
3604=>"000000101",
3605=>"001001001",
3606=>"010000011",
3607=>"100110101",
3608=>"011000001",
3609=>"000110111",
3610=>"000111011",
3611=>"001001111",
3612=>"110001101",
3613=>"000000101",
3614=>"111111001",
3615=>"001000000",
3616=>"000000111",
3617=>"001111111",
3618=>"001001000",
3619=>"011001001",
3620=>"011110010",
3621=>"100100100",
3622=>"111001001",
3623=>"001111110",
3624=>"001001101",
3625=>"001111111",
3626=>"111000000",
3627=>"100001000",
3628=>"000110110",
3629=>"011000111",
3630=>"000100111",
3631=>"111111000",
3632=>"000111111",
3633=>"000110100",
3634=>"001111000",
3635=>"111001101",
3636=>"010001000",
3637=>"001101110",
3638=>"000001001",
3639=>"001001001",
3640=>"011001111",
3641=>"000000111",
3642=>"110111001",
3643=>"001111111",
3644=>"010100110",
3645=>"111111000",
3646=>"000001000",
3647=>"011001000",
3648=>"001111110",
3649=>"100001110",
3650=>"110000100",
3651=>"111011000",
3652=>"011010001",
3653=>"001111000",
3654=>"000100110",
3655=>"000000010",
3656=>"001110110",
3657=>"000110110",
3658=>"111011011",
3659=>"110111100",
3660=>"000000000",
3661=>"000111101",
3662=>"010100110",
3663=>"101001000",
3664=>"011011000",
3665=>"110000101",
3666=>"000110111",
3667=>"000010011",
3668=>"111001001",
3669=>"001110001",
3670=>"101100000",
3671=>"000010000",
3672=>"000110000",
3673=>"000000100",
3674=>"111101101",
3675=>"011111111",
3676=>"010001011",
3677=>"000011010",
3678=>"111101001",
3679=>"001001001",
3680=>"000110010",
3681=>"001011011",
3682=>"100001001",
3683=>"111011101",
3684=>"000000101",
3685=>"000110010",
3686=>"001100000",
3687=>"000000001",
3688=>"000110111",
3689=>"111110000",
3690=>"001000000",
3691=>"100110110",
3692=>"101011111",
3693=>"111011110",
3694=>"110110000",
3695=>"000111111",
3696=>"111011011",
3697=>"000111111",
3698=>"010011001",
3699=>"000011111",
3700=>"000110000",
3701=>"111001011",
3702=>"111110110",
3703=>"010110100",
3704=>"111110000",
3705=>"000100000",
3706=>"000001011",
3707=>"000110110",
3708=>"011000111",
3709=>"000100100",
3710=>"001000111",
3711=>"111000000",
3712=>"000110100",
3713=>"111111111",
3714=>"011111010",
3715=>"001101000",
3716=>"000111111",
3717=>"001001000",
3718=>"100000100",
3719=>"001000010",
3720=>"000111110",
3721=>"111001101",
3722=>"000000101",
3723=>"101110010",
3724=>"010001101",
3725=>"000000110",
3726=>"111011011",
3727=>"110000001",
3728=>"011101111",
3729=>"001010001",
3730=>"110000001",
3731=>"010001000",
3732=>"000001001",
3733=>"110001001",
3734=>"001110011",
3735=>"000000010",
3736=>"000110110",
3737=>"111001001",
3738=>"111001001",
3739=>"111000001",
3740=>"000000011",
3741=>"111011001",
3742=>"001000001",
3743=>"111001011",
3744=>"001110111",
3745=>"011011111",
3746=>"000001110",
3747=>"011001000",
3748=>"001001010",
3749=>"000101100",
3750=>"101100000",
3751=>"110111001",
3752=>"000001001",
3753=>"111111111",
3754=>"111111001",
3755=>"110011001",
3756=>"000100000",
3757=>"110111111",
3758=>"011001110",
3759=>"001000100",
3760=>"101100100",
3761=>"010011111",
3762=>"110110111",
3763=>"000001011",
3764=>"000010110",
3765=>"101111000",
3766=>"000110110",
3767=>"000110110",
3768=>"100110110",
3769=>"000000101",
3770=>"001110100",
3771=>"111110110",
3772=>"111110000",
3773=>"010011011",
3774=>"100111011",
3775=>"001111110",
3776=>"001001111",
3777=>"000000000",
3778=>"111110000",
3779=>"000010001",
3780=>"111111110",
3781=>"000100010",
3782=>"000000110",
3783=>"010001000",
3784=>"001110110",
3785=>"111001001",
3786=>"001110100",
3787=>"001100110",
3788=>"000000010",
3789=>"001000110",
3790=>"111011000",
3791=>"000110000",
3792=>"111000001",
3793=>"000101111",
3794=>"000101101",
3795=>"001110110",
3796=>"111111100",
3797=>"110110100",
3798=>"111111000",
3799=>"000100001",
3800=>"000000111",
3801=>"001001001",
3802=>"001100110",
3803=>"100000000",
3804=>"001001001",
3805=>"001000001",
3806=>"000110110",
3807=>"100110001",
3808=>"110101000",
3809=>"010000001",
3810=>"101101111",
3811=>"001110110",
3812=>"000000111",
3813=>"010110110",
3814=>"011100110",
3815=>"001001101",
3816=>"000110111",
3817=>"000011111",
3818=>"110000000",
3819=>"011010110",
3820=>"111001000",
3821=>"000000110",
3822=>"010001000",
3823=>"110011101",
3824=>"101000011",
3825=>"110000010",
3826=>"000001001",
3827=>"000101100",
3828=>"000100010",
3829=>"110011001",
3830=>"010010110",
3831=>"011001001",
3832=>"001000001",
3833=>"101110110",
3834=>"000111111",
3835=>"001000010",
3836=>"100111101",
3837=>"001001000",
3838=>"000101001",
3839=>"111111100",
3840=>"111101111",
3841=>"000011111",
3842=>"000000010",
3843=>"101111111",
3844=>"000000001",
3845=>"110110000",
3846=>"001010011",
3847=>"000000011",
3848=>"001000000",
3849=>"000000000",
3850=>"111010010",
3851=>"111110000",
3852=>"010010000",
3853=>"010111011",
3854=>"100001011",
3855=>"000000100",
3856=>"111101000",
3857=>"000000000",
3858=>"110000000",
3859=>"101011011",
3860=>"111101101",
3861=>"111010000",
3862=>"000000011",
3863=>"000100000",
3864=>"000000000",
3865=>"000101101",
3866=>"110111110",
3867=>"001001100",
3868=>"000000100",
3869=>"000000000",
3870=>"110000011",
3871=>"111011000",
3872=>"111111111",
3873=>"111111111",
3874=>"101000000",
3875=>"111111101",
3876=>"100100111",
3877=>"111111111",
3878=>"111011010",
3879=>"001101001",
3880=>"000001111",
3881=>"110111111",
3882=>"000000000",
3883=>"010000011",
3884=>"111111111",
3885=>"000010000",
3886=>"111111111",
3887=>"111111111",
3888=>"111001111",
3889=>"001001001",
3890=>"101100110",
3891=>"001001111",
3892=>"011000000",
3893=>"011111100",
3894=>"001001000",
3895=>"111111000",
3896=>"111111110",
3897=>"000000000",
3898=>"000000000",
3899=>"001101111",
3900=>"011101101",
3901=>"111111110",
3902=>"000000000",
3903=>"001000010",
3904=>"101101101",
3905=>"111111111",
3906=>"101111111",
3907=>"000000100",
3908=>"000000000",
3909=>"000000000",
3910=>"100000111",
3911=>"101000010",
3912=>"111111100",
3913=>"000000110",
3914=>"000000000",
3915=>"111111101",
3916=>"011000000",
3917=>"000000000",
3918=>"001101011",
3919=>"111000110",
3920=>"000111111",
3921=>"000110010",
3922=>"111011011",
3923=>"111001100",
3924=>"000000000",
3925=>"000001100",
3926=>"111011110",
3927=>"000100100",
3928=>"111111001",
3929=>"010110011",
3930=>"100100101",
3931=>"101101111",
3932=>"111111000",
3933=>"011001011",
3934=>"000000000",
3935=>"000000001",
3936=>"100000000",
3937=>"111101000",
3938=>"100010101",
3939=>"101101100",
3940=>"110101111",
3941=>"111101000",
3942=>"100111000",
3943=>"000000000",
3944=>"000001001",
3945=>"000010110",
3946=>"010010111",
3947=>"110110111",
3948=>"111110110",
3949=>"000011111",
3950=>"011100000",
3951=>"000000111",
3952=>"111101101",
3953=>"000111111",
3954=>"101100001",
3955=>"111000001",
3956=>"010000000",
3957=>"101000011",
3958=>"000001111",
3959=>"000000110",
3960=>"000110000",
3961=>"111111111",
3962=>"100111000",
3963=>"000000001",
3964=>"100111111",
3965=>"100100100",
3966=>"000010110",
3967=>"000000001",
3968=>"001011000",
3969=>"111010010",
3970=>"111000000",
3971=>"000000000",
3972=>"110101101",
3973=>"001101101",
3974=>"101111111",
3975=>"101111100",
3976=>"111101111",
3977=>"001101110",
3978=>"100000000",
3979=>"000100101",
3980=>"000000000",
3981=>"000100111",
3982=>"111111110",
3983=>"100000101",
3984=>"010110011",
3985=>"110111111",
3986=>"001001111",
3987=>"111000010",
3988=>"001001101",
3989=>"000000101",
3990=>"110111000",
3991=>"001011111",
3992=>"111000000",
3993=>"000000000",
3994=>"111000000",
3995=>"000000000",
3996=>"010111000",
3997=>"101111111",
3998=>"111100100",
3999=>"101000000",
4000=>"000000001",
4001=>"000000011",
4002=>"000000000",
4003=>"010110110",
4004=>"010111111",
4005=>"000000000",
4006=>"010000000",
4007=>"000010010",
4008=>"000111111",
4009=>"101110111",
4010=>"010001111",
4011=>"000000101",
4012=>"110111111",
4013=>"111001101",
4014=>"010000011",
4015=>"010010000",
4016=>"000000000",
4017=>"110101101",
4018=>"000000000",
4019=>"000000001",
4020=>"000000101",
4021=>"000000000",
4022=>"101111111",
4023=>"111111111",
4024=>"111101111",
4025=>"111101101",
4026=>"111111111",
4027=>"000000110",
4028=>"111111110",
4029=>"111111111",
4030=>"100000101",
4031=>"000000000",
4032=>"000000000",
4033=>"100111110",
4034=>"101111111",
4035=>"010111111",
4036=>"000010000",
4037=>"010010100",
4038=>"000011010",
4039=>"000001100",
4040=>"101000010",
4041=>"000000000",
4042=>"111111111",
4043=>"101000111",
4044=>"000000100",
4045=>"011111111",
4046=>"000010011",
4047=>"100010110",
4048=>"000010000",
4049=>"110100110",
4050=>"111111110",
4051=>"000000000",
4052=>"101101111",
4053=>"101100110",
4054=>"110111000",
4055=>"111000001",
4056=>"000010000",
4057=>"111111111",
4058=>"000000110",
4059=>"000000000",
4060=>"000101011",
4061=>"011000000",
4062=>"000000111",
4063=>"011111111",
4064=>"000000000",
4065=>"111000101",
4066=>"000000000",
4067=>"110101110",
4068=>"000000111",
4069=>"010111010",
4070=>"111111110",
4071=>"101101100",
4072=>"110111101",
4073=>"000000100",
4074=>"011011011",
4075=>"010111000",
4076=>"000000000",
4077=>"000001111",
4078=>"000010010",
4079=>"011001101",
4080=>"000111011",
4081=>"010101000",
4082=>"111011000",
4083=>"011101000",
4084=>"111100111",
4085=>"000000100",
4086=>"000000000",
4087=>"101000000",
4088=>"000000111",
4089=>"000000000",
4090=>"000010011",
4091=>"001111001",
4092=>"000000100",
4093=>"100110101",
4094=>"000000000",
4095=>"000010010",
4096=>"010011000",
4097=>"000000000",
4098=>"100100101",
4099=>"011000000",
4100=>"001011011",
4101=>"001000000",
4102=>"010011000",
4103=>"000011010",
4104=>"110111111",
4105=>"000000000",
4106=>"111000011",
4107=>"000000010",
4108=>"010111000",
4109=>"010101000",
4110=>"011011001",
4111=>"001000000",
4112=>"010000111",
4113=>"010000111",
4114=>"000111000",
4115=>"001111111",
4116=>"010111101",
4117=>"100000100",
4118=>"001111101",
4119=>"111000011",
4120=>"001000000",
4121=>"111100100",
4122=>"000100101",
4123=>"111110000",
4124=>"111111111",
4125=>"000100100",
4126=>"011001101",
4127=>"000000000",
4128=>"000010010",
4129=>"110000000",
4130=>"111111000",
4131=>"000111011",
4132=>"001001001",
4133=>"011000000",
4134=>"000000110",
4135=>"000010000",
4136=>"100100100",
4137=>"000111000",
4138=>"101001111",
4139=>"000000100",
4140=>"001011011",
4141=>"000010110",
4142=>"011011111",
4143=>"100000100",
4144=>"000111111",
4145=>"110100001",
4146=>"111000011",
4147=>"000111111",
4148=>"010100111",
4149=>"011000000",
4150=>"110100111",
4151=>"000100110",
4152=>"100111000",
4153=>"000000011",
4154=>"111111000",
4155=>"100111111",
4156=>"110110110",
4157=>"101101000",
4158=>"000011001",
4159=>"110100111",
4160=>"010111100",
4161=>"111000000",
4162=>"001011000",
4163=>"000000000",
4164=>"000000000",
4165=>"000011000",
4166=>"000010000",
4167=>"011010100",
4168=>"000000110",
4169=>"111011011",
4170=>"010000000",
4171=>"101000000",
4172=>"000110111",
4173=>"110110110",
4174=>"011111110",
4175=>"100010001",
4176=>"000000001",
4177=>"110000000",
4178=>"000011111",
4179=>"001010110",
4180=>"011111011",
4181=>"001100110",
4182=>"110110100",
4183=>"101101001",
4184=>"100000000",
4185=>"010110100",
4186=>"100100100",
4187=>"111110110",
4188=>"000000000",
4189=>"001001001",
4190=>"111100111",
4191=>"010000000",
4192=>"000011011",
4193=>"001101000",
4194=>"111111000",
4195=>"100101101",
4196=>"000111110",
4197=>"011000000",
4198=>"110010000",
4199=>"100100111",
4200=>"101000110",
4201=>"111000100",
4202=>"010111000",
4203=>"000000000",
4204=>"000010011",
4205=>"111100011",
4206=>"000000011",
4207=>"011011000",
4208=>"101111001",
4209=>"000000000",
4210=>"011100110",
4211=>"111100010",
4212=>"011000000",
4213=>"000100111",
4214=>"000010001",
4215=>"111111110",
4216=>"111010111",
4217=>"111011000",
4218=>"111101100",
4219=>"000100000",
4220=>"100110011",
4221=>"110100101",
4222=>"111101111",
4223=>"100100011",
4224=>"001011111",
4225=>"110100100",
4226=>"100111000",
4227=>"111011000",
4228=>"000011111",
4229=>"001011111",
4230=>"111001000",
4231=>"000111000",
4232=>"110110100",
4233=>"000110110",
4234=>"011000111",
4235=>"001000100",
4236=>"101100100",
4237=>"000111110",
4238=>"011111000",
4239=>"111001000",
4240=>"001001000",
4241=>"000000000",
4242=>"100000111",
4243=>"000111111",
4244=>"000011110",
4245=>"001111001",
4246=>"000000101",
4247=>"110010000",
4248=>"000010111",
4249=>"111001111",
4250=>"000000100",
4251=>"000011101",
4252=>"000000000",
4253=>"011011010",
4254=>"110000000",
4255=>"000100010",
4256=>"100100000",
4257=>"010000111",
4258=>"111100000",
4259=>"011011011",
4260=>"100100111",
4261=>"111001000",
4262=>"010101101",
4263=>"011011011",
4264=>"010110111",
4265=>"000011111",
4266=>"100110111",
4267=>"011111000",
4268=>"111111000",
4269=>"111111001",
4270=>"110101001",
4271=>"111111010",
4272=>"100000000",
4273=>"000001000",
4274=>"010100100",
4275=>"111001100",
4276=>"111110111",
4277=>"000000111",
4278=>"011011000",
4279=>"000111001",
4280=>"001011001",
4281=>"000111011",
4282=>"010010000",
4283=>"101100011",
4284=>"100110000",
4285=>"101111011",
4286=>"011001001",
4287=>"000000011",
4288=>"101000100",
4289=>"100100111",
4290=>"000000010",
4291=>"000111100",
4292=>"111111010",
4293=>"001100011",
4294=>"010011111",
4295=>"010010100",
4296=>"100011011",
4297=>"100100000",
4298=>"010000000",
4299=>"000100110",
4300=>"111000000",
4301=>"000011010",
4302=>"111111101",
4303=>"111111100",
4304=>"000100111",
4305=>"011111011",
4306=>"100010000",
4307=>"100100010",
4308=>"010011010",
4309=>"100100010",
4310=>"000111111",
4311=>"111000001",
4312=>"110100111",
4313=>"000000111",
4314=>"110100011",
4315=>"011001000",
4316=>"110111110",
4317=>"101000111",
4318=>"001000100",
4319=>"000100010",
4320=>"111100100",
4321=>"000100100",
4322=>"011000000",
4323=>"111111110",
4324=>"011000000",
4325=>"011011100",
4326=>"000011000",
4327=>"010100100",
4328=>"000100001",
4329=>"000100111",
4330=>"111000001",
4331=>"000101000",
4332=>"010100100",
4333=>"000101000",
4334=>"010010000",
4335=>"000100111",
4336=>"111100111",
4337=>"101001010",
4338=>"000000011",
4339=>"100001111",
4340=>"010001001",
4341=>"001001010",
4342=>"000000010",
4343=>"111000000",
4344=>"000001000",
4345=>"000011111",
4346=>"100101000",
4347=>"000111111",
4348=>"100000111",
4349=>"000100110",
4350=>"101111111",
4351=>"011111000",
4352=>"000001111",
4353=>"000100101",
4354=>"000110111",
4355=>"111010000",
4356=>"011011010",
4357=>"101111001",
4358=>"001101001",
4359=>"111010111",
4360=>"000000010",
4361=>"100000000",
4362=>"101100101",
4363=>"010000000",
4364=>"000000000",
4365=>"010000000",
4366=>"011011010",
4367=>"000001011",
4368=>"111010000",
4369=>"000000111",
4370=>"000010010",
4371=>"001101000",
4372=>"000010010",
4373=>"001101111",
4374=>"100111111",
4375=>"010111111",
4376=>"000000100",
4377=>"101000110",
4378=>"000011010",
4379=>"111010000",
4380=>"000000010",
4381=>"101100000",
4382=>"001001001",
4383=>"110000000",
4384=>"000110000",
4385=>"110000111",
4386=>"000000110",
4387=>"110010000",
4388=>"111001000",
4389=>"000011110",
4390=>"110100000",
4391=>"010010001",
4392=>"010011111",
4393=>"110000011",
4394=>"000101111",
4395=>"000110110",
4396=>"011111111",
4397=>"101111010",
4398=>"101001000",
4399=>"000100110",
4400=>"110001000",
4401=>"011000010",
4402=>"010000101",
4403=>"001001101",
4404=>"110110110",
4405=>"011010010",
4406=>"000011011",
4407=>"101001000",
4408=>"000010010",
4409=>"111001000",
4410=>"000000000",
4411=>"111111001",
4412=>"111100100",
4413=>"010000100",
4414=>"000101001",
4415=>"011011111",
4416=>"111100111",
4417=>"100000110",
4418=>"101001000",
4419=>"001001111",
4420=>"001000000",
4421=>"000000000",
4422=>"101111100",
4423=>"001000111",
4424=>"111111001",
4425=>"000000000",
4426=>"000000000",
4427=>"101111111",
4428=>"000010010",
4429=>"111001000",
4430=>"110100000",
4431=>"001111111",
4432=>"000111111",
4433=>"100111010",
4434=>"110001101",
4435=>"001100010",
4436=>"000001001",
4437=>"100000110",
4438=>"011010000",
4439=>"000101111",
4440=>"001001101",
4441=>"111000000",
4442=>"101101111",
4443=>"111110011",
4444=>"001001111",
4445=>"001110000",
4446=>"110000000",
4447=>"100001110",
4448=>"101111000",
4449=>"011111010",
4450=>"000111110",
4451=>"011011111",
4452=>"110000000",
4453=>"011000000",
4454=>"111001000",
4455=>"000101010",
4456=>"111001000",
4457=>"000011101",
4458=>"111010011",
4459=>"000010100",
4460=>"110010010",
4461=>"110000111",
4462=>"000000110",
4463=>"111110000",
4464=>"111000110",
4465=>"111010000",
4466=>"000111011",
4467=>"111000000",
4468=>"111110100",
4469=>"000111000",
4470=>"111000000",
4471=>"100111110",
4472=>"000111111",
4473=>"000101000",
4474=>"110010001",
4475=>"111001111",
4476=>"110110000",
4477=>"100001000",
4478=>"101111011",
4479=>"000001111",
4480=>"111111000",
4481=>"100000000",
4482=>"111101000",
4483=>"111010001",
4484=>"000000000",
4485=>"010001111",
4486=>"001011011",
4487=>"101000000",
4488=>"011000011",
4489=>"110101001",
4490=>"000010001",
4491=>"110000001",
4492=>"000100100",
4493=>"000001111",
4494=>"101011110",
4495=>"001000000",
4496=>"000110100",
4497=>"010111000",
4498=>"111111001",
4499=>"000101101",
4500=>"111000001",
4501=>"000001111",
4502=>"010011101",
4503=>"011000000",
4504=>"001000000",
4505=>"000000111",
4506=>"001000010",
4507=>"000101111",
4508=>"101000000",
4509=>"010010101",
4510=>"111111111",
4511=>"001000001",
4512=>"111111110",
4513=>"001001111",
4514=>"000000010",
4515=>"000111111",
4516=>"000000000",
4517=>"100000111",
4518=>"110000000",
4519=>"010010010",
4520=>"000111111",
4521=>"111000011",
4522=>"000000111",
4523=>"000101111",
4524=>"000000000",
4525=>"000100000",
4526=>"001010011",
4527=>"111110001",
4528=>"010001001",
4529=>"000011001",
4530=>"000000000",
4531=>"011000111",
4532=>"101110011",
4533=>"011111111",
4534=>"111010000",
4535=>"010000000",
4536=>"111001001",
4537=>"111000000",
4538=>"110100010",
4539=>"110000111",
4540=>"110000000",
4541=>"010111111",
4542=>"011001011",
4543=>"000000000",
4544=>"101111100",
4545=>"000100111",
4546=>"010001000",
4547=>"001000000",
4548=>"010000000",
4549=>"001011001",
4550=>"010000000",
4551=>"000111001",
4552=>"111010000",
4553=>"111101110",
4554=>"000010100",
4555=>"111010000",
4556=>"100100100",
4557=>"101010000",
4558=>"101111010",
4559=>"110111111",
4560=>"011010000",
4561=>"110010001",
4562=>"110010000",
4563=>"110001010",
4564=>"000100111",
4565=>"110111100",
4566=>"000111101",
4567=>"111000011",
4568=>"111001000",
4569=>"111010011",
4570=>"111011111",
4571=>"001000111",
4572=>"011111111",
4573=>"000000011",
4574=>"000000111",
4575=>"111001000",
4576=>"000111110",
4577=>"001001011",
4578=>"010100101",
4579=>"010100111",
4580=>"001101111",
4581=>"011000000",
4582=>"111011101",
4583=>"111011101",
4584=>"111000000",
4585=>"000110011",
4586=>"100111111",
4587=>"001111111",
4588=>"000000010",
4589=>"110000000",
4590=>"000000000",
4591=>"101111001",
4592=>"110000000",
4593=>"000110110",
4594=>"000111000",
4595=>"100011110",
4596=>"111100001",
4597=>"001001111",
4598=>"000001010",
4599=>"100000011",
4600=>"101110111",
4601=>"111000000",
4602=>"111101010",
4603=>"111000000",
4604=>"000111111",
4605=>"000000100",
4606=>"110100110",
4607=>"000100110",
4608=>"001011011",
4609=>"001100011",
4610=>"000001101",
4611=>"000000000",
4612=>"011001001",
4613=>"000000110",
4614=>"000000101",
4615=>"110110011",
4616=>"111000010",
4617=>"101100111",
4618=>"101101100",
4619=>"000000101",
4620=>"100010110",
4621=>"001000110",
4622=>"000010000",
4623=>"000000011",
4624=>"001000000",
4625=>"111111111",
4626=>"100100111",
4627=>"000000010",
4628=>"010000000",
4629=>"000010000",
4630=>"110000000",
4631=>"101000111",
4632=>"110100010",
4633=>"001101111",
4634=>"000010110",
4635=>"110100000",
4636=>"100111111",
4637=>"111111011",
4638=>"000000000",
4639=>"101010111",
4640=>"101101010",
4641=>"111011000",
4642=>"111111111",
4643=>"100000000",
4644=>"011011111",
4645=>"000101011",
4646=>"111110000",
4647=>"111111111",
4648=>"110100100",
4649=>"111110111",
4650=>"001000101",
4651=>"000010000",
4652=>"101111111",
4653=>"000000001",
4654=>"000000101",
4655=>"011111010",
4656=>"001001000",
4657=>"011000001",
4658=>"000000000",
4659=>"111111100",
4660=>"000000100",
4661=>"111000000",
4662=>"110110011",
4663=>"110000000",
4664=>"111111010",
4665=>"000000110",
4666=>"000100000",
4667=>"110011000",
4668=>"010100000",
4669=>"110111011",
4670=>"001000100",
4671=>"110110110",
4672=>"101000101",
4673=>"000110111",
4674=>"000000000",
4675=>"111001110",
4676=>"000110010",
4677=>"010000000",
4678=>"000000000",
4679=>"000000011",
4680=>"110011111",
4681=>"000000010",
4682=>"101000111",
4683=>"001000110",
4684=>"111110111",
4685=>"110000010",
4686=>"110010100",
4687=>"101010111",
4688=>"001111001",
4689=>"011001000",
4690=>"000000011",
4691=>"011000001",
4692=>"001111111",
4693=>"100111111",
4694=>"000001111",
4695=>"000000101",
4696=>"000001000",
4697=>"111110011",
4698=>"000011001",
4699=>"100000110",
4700=>"101101110",
4701=>"001011011",
4702=>"010110111",
4703=>"110100111",
4704=>"110110110",
4705=>"001000100",
4706=>"111111101",
4707=>"011011100",
4708=>"010010000",
4709=>"111111111",
4710=>"001001101",
4711=>"111110000",
4712=>"000110111",
4713=>"000001000",
4714=>"011000111",
4715=>"000000100",
4716=>"111110110",
4717=>"000001001",
4718=>"001101000",
4719=>"110101100",
4720=>"011100001",
4721=>"000001101",
4722=>"101110111",
4723=>"011010001",
4724=>"000000000",
4725=>"000000010",
4726=>"111110111",
4727=>"111110010",
4728=>"110101101",
4729=>"111101010",
4730=>"101000110",
4731=>"101100010",
4732=>"001000100",
4733=>"100100100",
4734=>"111111100",
4735=>"000000001",
4736=>"110011110",
4737=>"000011001",
4738=>"000000000",
4739=>"111101000",
4740=>"000010101",
4741=>"111111110",
4742=>"000110110",
4743=>"011000001",
4744=>"000011000",
4745=>"011011110",
4746=>"100000100",
4747=>"010000000",
4748=>"010010011",
4749=>"001000000",
4750=>"010000000",
4751=>"000000001",
4752=>"001001100",
4753=>"010111110",
4754=>"001011111",
4755=>"001000000",
4756=>"111001000",
4757=>"001100000",
4758=>"101000111",
4759=>"111111000",
4760=>"101000000",
4761=>"000000001",
4762=>"000000111",
4763=>"000000101",
4764=>"000000101",
4765=>"110110010",
4766=>"010001000",
4767=>"000000111",
4768=>"110101011",
4769=>"111101001",
4770=>"111000111",
4771=>"101101111",
4772=>"010011111",
4773=>"111010000",
4774=>"110110000",
4775=>"001101111",
4776=>"000011111",
4777=>"111110111",
4778=>"000000101",
4779=>"000000100",
4780=>"111111011",
4781=>"000011101",
4782=>"111101111",
4783=>"010110111",
4784=>"000111111",
4785=>"011011101",
4786=>"000110100",
4787=>"111011000",
4788=>"111010001",
4789=>"110000010",
4790=>"111111111",
4791=>"000111111",
4792=>"010000001",
4793=>"101100000",
4794=>"111000000",
4795=>"000001010",
4796=>"001001000",
4797=>"111111111",
4798=>"111100000",
4799=>"111111000",
4800=>"000000101",
4801=>"000000000",
4802=>"001111110",
4803=>"100010110",
4804=>"010110011",
4805=>"010110111",
4806=>"000001011",
4807=>"000001111",
4808=>"101001111",
4809=>"110010000",
4810=>"111111110",
4811=>"010010000",
4812=>"111000010",
4813=>"100000001",
4814=>"001000100",
4815=>"111111000",
4816=>"111011111",
4817=>"100100100",
4818=>"001101111",
4819=>"000101111",
4820=>"101111010",
4821=>"100111111",
4822=>"000001111",
4823=>"001111011",
4824=>"101111111",
4825=>"110000000",
4826=>"111111111",
4827=>"001001101",
4828=>"011111010",
4829=>"011000000",
4830=>"001111000",
4831=>"001101111",
4832=>"000000000",
4833=>"000000100",
4834=>"010000000",
4835=>"101101101",
4836=>"101111111",
4837=>"111110110",
4838=>"111000000",
4839=>"111101110",
4840=>"111011111",
4841=>"111111010",
4842=>"001001101",
4843=>"000000101",
4844=>"110010000",
4845=>"001001110",
4846=>"000000000",
4847=>"101100000",
4848=>"000000010",
4849=>"001000111",
4850=>"000000000",
4851=>"101000100",
4852=>"101100101",
4853=>"000100110",
4854=>"000000000",
4855=>"000110110",
4856=>"101001101",
4857=>"101111110",
4858=>"100100000",
4859=>"101101111",
4860=>"000000111",
4861=>"000111001",
4862=>"100100100",
4863=>"000110010",
4864=>"000100010",
4865=>"000000101",
4866=>"000000001",
4867=>"001111011",
4868=>"001000110",
4869=>"111111111",
4870=>"101100111",
4871=>"111111111",
4872=>"110111111",
4873=>"000000000",
4874=>"111111100",
4875=>"010111000",
4876=>"000000000",
4877=>"000010010",
4878=>"001100101",
4879=>"000101101",
4880=>"111101110",
4881=>"000000111",
4882=>"000000010",
4883=>"111110010",
4884=>"111111111",
4885=>"010010110",
4886=>"001000101",
4887=>"111001001",
4888=>"000111010",
4889=>"000000100",
4890=>"001111110",
4891=>"010110110",
4892=>"100100000",
4893=>"111111111",
4894=>"001101001",
4895=>"000000010",
4896=>"100001111",
4897=>"111001000",
4898=>"001100000",
4899=>"000000000",
4900=>"000000100",
4901=>"000000101",
4902=>"001001110",
4903=>"000001010",
4904=>"000011111",
4905=>"110100011",
4906=>"011000101",
4907=>"010000111",
4908=>"111111100",
4909=>"111011000",
4910=>"100100110",
4911=>"010010010",
4912=>"000000010",
4913=>"011101011",
4914=>"000001010",
4915=>"100111111",
4916=>"101101111",
4917=>"011111111",
4918=>"001000101",
4919=>"000000000",
4920=>"110000111",
4921=>"000000000",
4922=>"101011011",
4923=>"000101000",
4924=>"100111101",
4925=>"111011111",
4926=>"001000111",
4927=>"110111111",
4928=>"000111100",
4929=>"101000000",
4930=>"000000000",
4931=>"101000110",
4932=>"000001101",
4933=>"000000010",
4934=>"000101111",
4935=>"101000110",
4936=>"011111111",
4937=>"101101111",
4938=>"000000111",
4939=>"111101011",
4940=>"000111111",
4941=>"001001001",
4942=>"100010000",
4943=>"111101001",
4944=>"000000101",
4945=>"011001000",
4946=>"110000000",
4947=>"000000001",
4948=>"000000000",
4949=>"011011011",
4950=>"001011010",
4951=>"000000000",
4952=>"101111101",
4953=>"001000101",
4954=>"111011011",
4955=>"000101000",
4956=>"000000001",
4957=>"000000111",
4958=>"111111111",
4959=>"000000101",
4960=>"101111111",
4961=>"111111111",
4962=>"000000000",
4963=>"111111110",
4964=>"000000000",
4965=>"111111100",
4966=>"111111010",
4967=>"000111111",
4968=>"101111111",
4969=>"111111010",
4970=>"000001111",
4971=>"111111110",
4972=>"111000001",
4973=>"111111111",
4974=>"000000111",
4975=>"101111111",
4976=>"111110010",
4977=>"101101000",
4978=>"001001111",
4979=>"110111000",
4980=>"000000011",
4981=>"000000110",
4982=>"111000010",
4983=>"000101010",
4984=>"010111111",
4985=>"101000110",
4986=>"110000001",
4987=>"111110010",
4988=>"000001001",
4989=>"100000000",
4990=>"110000111",
4991=>"000000111",
4992=>"001000000",
4993=>"111000000",
4994=>"110111111",
4995=>"000000000",
4996=>"111100000",
4997=>"111111111",
4998=>"100001111",
4999=>"000000000",
5000=>"100101101",
5001=>"101100000",
5002=>"000001111",
5003=>"000000000",
5004=>"000111111",
5005=>"110111000",
5006=>"000000010",
5007=>"001000100",
5008=>"111000000",
5009=>"111000000",
5010=>"111001111",
5011=>"111100101",
5012=>"010111000",
5013=>"000000100",
5014=>"001101111",
5015=>"100001010",
5016=>"111111011",
5017=>"101110001",
5018=>"011111101",
5019=>"010110110",
5020=>"111001000",
5021=>"110111111",
5022=>"000000011",
5023=>"000000000",
5024=>"110100100",
5025=>"000101111",
5026=>"000000100",
5027=>"001001000",
5028=>"101011100",
5029=>"000000000",
5030=>"000111011",
5031=>"000000100",
5032=>"111010101",
5033=>"000001111",
5034=>"111111010",
5035=>"111000001",
5036=>"001111111",
5037=>"000000100",
5038=>"011100111",
5039=>"111011100",
5040=>"101111000",
5041=>"100000101",
5042=>"000001011",
5043=>"000000011",
5044=>"111110111",
5045=>"001001000",
5046=>"000000000",
5047=>"101001000",
5048=>"011100011",
5049=>"111101001",
5050=>"110000011",
5051=>"000111111",
5052=>"111111010",
5053=>"111000111",
5054=>"111111110",
5055=>"001001011",
5056=>"000000000",
5057=>"111111000",
5058=>"111110011",
5059=>"000000010",
5060=>"010001000",
5061=>"111011111",
5062=>"110110100",
5063=>"111011000",
5064=>"100001010",
5065=>"000001000",
5066=>"000001101",
5067=>"111111100",
5068=>"100111111",
5069=>"000100100",
5070=>"000001111",
5071=>"000110111",
5072=>"010111010",
5073=>"100000001",
5074=>"000000111",
5075=>"000000000",
5076=>"000000000",
5077=>"001000110",
5078=>"000000000",
5079=>"101000010",
5080=>"000001000",
5081=>"010010100",
5082=>"010001001",
5083=>"111110000",
5084=>"010001100",
5085=>"110010111",
5086=>"000000000",
5087=>"111111000",
5088=>"000001000",
5089=>"001000101",
5090=>"010111111",
5091=>"110011011",
5092=>"000000110",
5093=>"111111111",
5094=>"111001000",
5095=>"000011011",
5096=>"010010010",
5097=>"100000000",
5098=>"111111101",
5099=>"000000000",
5100=>"011000100",
5101=>"001100110",
5102=>"000000000",
5103=>"000001000",
5104=>"111111010",
5105=>"111100110",
5106=>"010000000",
5107=>"110011111",
5108=>"100000110",
5109=>"100110011",
5110=>"010000000",
5111=>"010101111",
5112=>"000000001",
5113=>"011101001",
5114=>"101000111",
5115=>"000110010",
5116=>"010111010",
5117=>"100110100",
5118=>"000001010",
5119=>"111000000",
5120=>"000011000",
5121=>"111111111",
5122=>"000010000",
5123=>"111101111",
5124=>"000000000",
5125=>"111110000",
5126=>"000111011",
5127=>"000111111",
5128=>"000000111",
5129=>"001000011",
5130=>"111111011",
5131=>"111111011",
5132=>"000000101",
5133=>"101011001",
5134=>"001001000",
5135=>"001000111",
5136=>"001000111",
5137=>"111110111",
5138=>"110110000",
5139=>"000000000",
5140=>"110111100",
5141=>"000110000",
5142=>"000000011",
5143=>"111101001",
5144=>"000000001",
5145=>"000000110",
5146=>"010010000",
5147=>"010000000",
5148=>"011001000",
5149=>"000010000",
5150=>"110000000",
5151=>"000111000",
5152=>"111000001",
5153=>"111111111",
5154=>"001111000",
5155=>"000101010",
5156=>"000000000",
5157=>"000011000",
5158=>"111001011",
5159=>"000000000",
5160=>"000001111",
5161=>"111010000",
5162=>"111000000",
5163=>"110001011",
5164=>"000001000",
5165=>"101011000",
5166=>"111111111",
5167=>"101111101",
5168=>"101111000",
5169=>"000000001",
5170=>"111111011",
5171=>"111110111",
5172=>"110111111",
5173=>"101001101",
5174=>"110111111",
5175=>"100111111",
5176=>"111100001",
5177=>"000000101",
5178=>"010011010",
5179=>"001100111",
5180=>"110111111",
5181=>"111111000",
5182=>"000000000",
5183=>"000000000",
5184=>"000111111",
5185=>"000000000",
5186=>"010111110",
5187=>"000000110",
5188=>"011011000",
5189=>"010000000",
5190=>"000111111",
5191=>"111111001",
5192=>"000000000",
5193=>"011111111",
5194=>"000000100",
5195=>"001000101",
5196=>"111000010",
5197=>"000000001",
5198=>"000000000",
5199=>"010110000",
5200=>"111111111",
5201=>"000000000",
5202=>"010011111",
5203=>"101000000",
5204=>"110110001",
5205=>"111111011",
5206=>"000000000",
5207=>"110111010",
5208=>"001000000",
5209=>"000000001",
5210=>"000000000",
5211=>"000000000",
5212=>"000000111",
5213=>"000000000",
5214=>"111110000",
5215=>"100100011",
5216=>"111111111",
5217=>"101111100",
5218=>"000000111",
5219=>"000000000",
5220=>"000100101",
5221=>"000000111",
5222=>"010111101",
5223=>"100001000",
5224=>"100111101",
5225=>"011100111",
5226=>"111111101",
5227=>"111111111",
5228=>"010111111",
5229=>"111111000",
5230=>"111000000",
5231=>"001010100",
5232=>"000000000",
5233=>"010111000",
5234=>"011101110",
5235=>"111010000",
5236=>"111111000",
5237=>"000000100",
5238=>"110000110",
5239=>"111000000",
5240=>"111101001",
5241=>"111111000",
5242=>"111001101",
5243=>"000000000",
5244=>"101111111",
5245=>"000000000",
5246=>"101111000",
5247=>"000000111",
5248=>"111111000",
5249=>"111000010",
5250=>"101100111",
5251=>"101111100",
5252=>"111111000",
5253=>"111111000",
5254=>"111110010",
5255=>"000000100",
5256=>"000000000",
5257=>"110111001",
5258=>"001111000",
5259=>"110000011",
5260=>"101000100",
5261=>"000011111",
5262=>"000000000",
5263=>"101000010",
5264=>"000000000",
5265=>"000000100",
5266=>"101000111",
5267=>"000000001",
5268=>"000000000",
5269=>"111000110",
5270=>"000111111",
5271=>"000000000",
5272=>"101000110",
5273=>"110111110",
5274=>"101111110",
5275=>"111111111",
5276=>"000001001",
5277=>"111010001",
5278=>"111111111",
5279=>"000000111",
5280=>"100101000",
5281=>"000111100",
5282=>"001111000",
5283=>"100111000",
5284=>"101100000",
5285=>"000000000",
5286=>"000000000",
5287=>"001111000",
5288=>"111111000",
5289=>"111111000",
5290=>"101000111",
5291=>"000000100",
5292=>"111101000",
5293=>"000000000",
5294=>"001101100",
5295=>"001111111",
5296=>"001111111",
5297=>"000000001",
5298=>"000000011",
5299=>"001000000",
5300=>"000000000",
5301=>"000110100",
5302=>"011111000",
5303=>"110001000",
5304=>"111111111",
5305=>"000000001",
5306=>"000111000",
5307=>"111111111",
5308=>"111111001",
5309=>"110000110",
5310=>"000000000",
5311=>"011111111",
5312=>"000000000",
5313=>"000000100",
5314=>"111111000",
5315=>"110001101",
5316=>"000111000",
5317=>"001011000",
5318=>"111110111",
5319=>"000000110",
5320=>"000000001",
5321=>"110010000",
5322=>"011001110",
5323=>"011000101",
5324=>"001001001",
5325=>"100111111",
5326=>"000000111",
5327=>"111111000",
5328=>"000000000",
5329=>"000000000",
5330=>"111111111",
5331=>"111100000",
5332=>"101000101",
5333=>"000000001",
5334=>"111111011",
5335=>"111111101",
5336=>"001101101",
5337=>"011111101",
5338=>"000001001",
5339=>"111000001",
5340=>"111001000",
5341=>"111111001",
5342=>"101101110",
5343=>"100111111",
5344=>"000000110",
5345=>"101100111",
5346=>"000000001",
5347=>"001000000",
5348=>"001000010",
5349=>"111111000",
5350=>"000000000",
5351=>"000000001",
5352=>"111111110",
5353=>"000000111",
5354=>"111111110",
5355=>"010110011",
5356=>"111110010",
5357=>"000000000",
5358=>"010000000",
5359=>"000000001",
5360=>"111111000",
5361=>"000000000",
5362=>"110111000",
5363=>"000000000",
5364=>"000000000",
5365=>"111111101",
5366=>"111111000",
5367=>"101011000",
5368=>"000001111",
5369=>"101111111",
5370=>"111111111",
5371=>"001101001",
5372=>"000000111",
5373=>"111111001",
5374=>"000000000",
5375=>"000110110",
5376=>"101100110",
5377=>"111111000",
5378=>"000010000",
5379=>"000000000",
5380=>"000011111",
5381=>"000000001",
5382=>"010111111",
5383=>"010110100",
5384=>"101001000",
5385=>"010000000",
5386=>"010111111",
5387=>"000000000",
5388=>"100000000",
5389=>"101100101",
5390=>"000000000",
5391=>"000000000",
5392=>"000000010",
5393=>"111111001",
5394=>"110111000",
5395=>"111011000",
5396=>"110111111",
5397=>"111101111",
5398=>"111111010",
5399=>"000010100",
5400=>"111111000",
5401=>"111000111",
5402=>"111100000",
5403=>"111111000",
5404=>"000000001",
5405=>"000001101",
5406=>"101111111",
5407=>"000000100",
5408=>"010011111",
5409=>"000000100",
5410=>"101111110",
5411=>"111101111",
5412=>"110110100",
5413=>"000001011",
5414=>"110000100",
5415=>"000001111",
5416=>"000000110",
5417=>"111100111",
5418=>"010001111",
5419=>"000000000",
5420=>"111111111",
5421=>"111100000",
5422=>"110111011",
5423=>"011111101",
5424=>"001011010",
5425=>"010110110",
5426=>"111101111",
5427=>"001011111",
5428=>"111111111",
5429=>"111111111",
5430=>"110000000",
5431=>"101010010",
5432=>"000111111",
5433=>"000000100",
5434=>"000000000",
5435=>"010010000",
5436=>"000000001",
5437=>"111010111",
5438=>"001000000",
5439=>"111111110",
5440=>"000010010",
5441=>"000011111",
5442=>"000001111",
5443=>"000010000",
5444=>"100000100",
5445=>"000001111",
5446=>"111000000",
5447=>"001001101",
5448=>"011100010",
5449=>"100100010",
5450=>"000000000",
5451=>"000000010",
5452=>"110101001",
5453=>"011110010",
5454=>"110111011",
5455=>"001001011",
5456=>"100111111",
5457=>"111000010",
5458=>"100000000",
5459=>"000010000",
5460=>"001000000",
5461=>"000110111",
5462=>"000110011",
5463=>"000000100",
5464=>"001001011",
5465=>"000001111",
5466=>"000111100",
5467=>"111111011",
5468=>"100000100",
5469=>"110110000",
5470=>"010111110",
5471=>"011001000",
5472=>"111111111",
5473=>"001101100",
5474=>"001000000",
5475=>"011111111",
5476=>"010011110",
5477=>"000000110",
5478=>"101100100",
5479=>"010011111",
5480=>"111110011",
5481=>"000010000",
5482=>"000000000",
5483=>"000000111",
5484=>"101000101",
5485=>"010111111",
5486=>"001000001",
5487=>"010000000",
5488=>"011111111",
5489=>"000000000",
5490=>"111000100",
5491=>"000111010",
5492=>"000000100",
5493=>"000000011",
5494=>"100000000",
5495=>"010000000",
5496=>"000100000",
5497=>"111111111",
5498=>"011011010",
5499=>"101100000",
5500=>"011001000",
5501=>"001011110",
5502=>"001110110",
5503=>"100000011",
5504=>"001111001",
5505=>"011011011",
5506=>"010111111",
5507=>"000011100",
5508=>"000000111",
5509=>"111110111",
5510=>"000100110",
5511=>"100100100",
5512=>"111111111",
5513=>"001101000",
5514=>"000111000",
5515=>"000010010",
5516=>"100110011",
5517=>"111010001",
5518=>"000000100",
5519=>"000000000",
5520=>"011000111",
5521=>"101010110",
5522=>"010011011",
5523=>"100001000",
5524=>"111000000",
5525=>"110000100",
5526=>"111111111",
5527=>"111100111",
5528=>"111111111",
5529=>"111000000",
5530=>"111111000",
5531=>"001000001",
5532=>"100000100",
5533=>"110111111",
5534=>"111111001",
5535=>"111000000",
5536=>"111010010",
5537=>"111111111",
5538=>"111000110",
5539=>"001011000",
5540=>"000010011",
5541=>"111011000",
5542=>"000010010",
5543=>"000011111",
5544=>"111111110",
5545=>"010010001",
5546=>"101000000",
5547=>"101100000",
5548=>"000110111",
5549=>"100000000",
5550=>"101001110",
5551=>"001111000",
5552=>"111000100",
5553=>"000100101",
5554=>"000000000",
5555=>"111100000",
5556=>"111101011",
5557=>"000110011",
5558=>"000000011",
5559=>"000101111",
5560=>"000100000",
5561=>"000000000",
5562=>"111101000",
5563=>"010000100",
5564=>"000100100",
5565=>"000010010",
5566=>"110100000",
5567=>"111111111",
5568=>"000000000",
5569=>"000000000",
5570=>"000011000",
5571=>"110111111",
5572=>"000000111",
5573=>"010111110",
5574=>"111011111",
5575=>"000100111",
5576=>"000000000",
5577=>"000100000",
5578=>"000010001",
5579=>"111000111",
5580=>"011000000",
5581=>"110100100",
5582=>"000111111",
5583=>"111011011",
5584=>"011111111",
5585=>"011101111",
5586=>"001000100",
5587=>"001111111",
5588=>"101000101",
5589=>"101111110",
5590=>"000000000",
5591=>"001000000",
5592=>"000110111",
5593=>"101111101",
5594=>"111011111",
5595=>"000111111",
5596=>"000111010",
5597=>"010111111",
5598=>"101001111",
5599=>"000000010",
5600=>"101000000",
5601=>"000011000",
5602=>"011111110",
5603=>"111111000",
5604=>"111000100",
5605=>"000011000",
5606=>"011011001",
5607=>"101000100",
5608=>"111101010",
5609=>"111101111",
5610=>"111111110",
5611=>"111100000",
5612=>"000001001",
5613=>"111111111",
5614=>"111000000",
5615=>"000000111",
5616=>"000010110",
5617=>"010111111",
5618=>"011001000",
5619=>"001011001",
5620=>"011011011",
5621=>"111111111",
5622=>"000010111",
5623=>"000000000",
5624=>"000000111",
5625=>"000000100",
5626=>"000000000",
5627=>"010000000",
5628=>"101100101",
5629=>"000000000",
5630=>"111111011",
5631=>"000011011",
5632=>"011110100",
5633=>"000100000",
5634=>"000000110",
5635=>"110010101",
5636=>"100100000",
5637=>"000000000",
5638=>"111101000",
5639=>"000001010",
5640=>"110010010",
5641=>"010110000",
5642=>"100010011",
5643=>"010000001",
5644=>"000000000",
5645=>"010111011",
5646=>"111111111",
5647=>"000101101",
5648=>"001000000",
5649=>"101000110",
5650=>"111000110",
5651=>"001000000",
5652=>"000100101",
5653=>"111111110",
5654=>"000110100",
5655=>"101101110",
5656=>"000000000",
5657=>"111111111",
5658=>"111111111",
5659=>"110110100",
5660=>"111111111",
5661=>"000000000",
5662=>"000001001",
5663=>"000000101",
5664=>"000001000",
5665=>"010101111",
5666=>"000111011",
5667=>"011111111",
5668=>"001111101",
5669=>"000000011",
5670=>"000111111",
5671=>"111001011",
5672=>"010010000",
5673=>"000111111",
5674=>"111111111",
5675=>"110001110",
5676=>"001011100",
5677=>"000000101",
5678=>"011000101",
5679=>"100000001",
5680=>"000000100",
5681=>"001111111",
5682=>"000011110",
5683=>"001011010",
5684=>"100000000",
5685=>"000000111",
5686=>"010110100",
5687=>"000010000",
5688=>"011001010",
5689=>"100000001",
5690=>"000000000",
5691=>"000100001",
5692=>"110011110",
5693=>"111111111",
5694=>"000111000",
5695=>"000100110",
5696=>"000000000",
5697=>"000000100",
5698=>"111111111",
5699=>"000000000",
5700=>"000000001",
5701=>"101001101",
5702=>"100111000",
5703=>"100101111",
5704=>"101101110",
5705=>"010000000",
5706=>"000000000",
5707=>"000000010",
5708=>"111111111",
5709=>"001111001",
5710=>"011011011",
5711=>"101111011",
5712=>"101111111",
5713=>"000011110",
5714=>"000101011",
5715=>"001000100",
5716=>"000000000",
5717=>"000001100",
5718=>"101111011",
5719=>"010111110",
5720=>"110110110",
5721=>"100110110",
5722=>"100101101",
5723=>"110100000",
5724=>"001100110",
5725=>"001001001",
5726=>"011001100",
5727=>"010000000",
5728=>"110010010",
5729=>"110000001",
5730=>"010111011",
5731=>"111101101",
5732=>"111110110",
5733=>"010101011",
5734=>"010010010",
5735=>"011111010",
5736=>"100001001",
5737=>"101000000",
5738=>"001001000",
5739=>"111110101",
5740=>"111111111",
5741=>"111111110",
5742=>"100100100",
5743=>"111010010",
5744=>"000111001",
5745=>"100000011",
5746=>"000111001",
5747=>"001001001",
5748=>"001001001",
5749=>"000000000",
5750=>"000100010",
5751=>"111010001",
5752=>"001101110",
5753=>"111001000",
5754=>"111001111",
5755=>"000000110",
5756=>"100111001",
5757=>"000000000",
5758=>"000000010",
5759=>"000000000",
5760=>"101111111",
5761=>"000100110",
5762=>"010000000",
5763=>"111111011",
5764=>"101001001",
5765=>"001100100",
5766=>"001000000",
5767=>"000100111",
5768=>"001011100",
5769=>"000000000",
5770=>"111000000",
5771=>"011000110",
5772=>"110000000",
5773=>"000000000",
5774=>"101000111",
5775=>"000001000",
5776=>"100011111",
5777=>"000001101",
5778=>"001101110",
5779=>"111100010",
5780=>"000000000",
5781=>"000010010",
5782=>"010111111",
5783=>"011010001",
5784=>"110110110",
5785=>"000001000",
5786=>"010000010",
5787=>"000000110",
5788=>"010000000",
5789=>"001010010",
5790=>"001000000",
5791=>"011010000",
5792=>"100111111",
5793=>"101100000",
5794=>"111101111",
5795=>"110110110",
5796=>"001000000",
5797=>"011011001",
5798=>"011111111",
5799=>"011011111",
5800=>"000000100",
5801=>"000000111",
5802=>"100000111",
5803=>"000001000",
5804=>"011101001",
5805=>"111111111",
5806=>"100101001",
5807=>"111111111",
5808=>"000000010",
5809=>"011011010",
5810=>"101100100",
5811=>"100011110",
5812=>"100000100",
5813=>"111110111",
5814=>"100111010",
5815=>"000100111",
5816=>"011110111",
5817=>"100000001",
5818=>"111010011",
5819=>"111010000",
5820=>"111111111",
5821=>"010111110",
5822=>"110011011",
5823=>"100111111",
5824=>"000010111",
5825=>"000000000",
5826=>"101101100",
5827=>"001100111",
5828=>"010001110",
5829=>"110100111",
5830=>"110110000",
5831=>"000000000",
5832=>"001111111",
5833=>"000000000",
5834=>"111111001",
5835=>"001000010",
5836=>"011000000",
5837=>"001110110",
5838=>"000000000",
5839=>"110000000",
5840=>"000000111",
5841=>"110110110",
5842=>"110000110",
5843=>"001001001",
5844=>"001001000",
5845=>"100100100",
5846=>"111011011",
5847=>"000000111",
5848=>"111101111",
5849=>"011011111",
5850=>"010111110",
5851=>"000000000",
5852=>"000100001",
5853=>"000011110",
5854=>"100001010",
5855=>"011010000",
5856=>"110111010",
5857=>"100100000",
5858=>"011100111",
5859=>"111111110",
5860=>"101000010",
5861=>"000000000",
5862=>"111110000",
5863=>"011111001",
5864=>"000101100",
5865=>"100000000",
5866=>"010010110",
5867=>"011000101",
5868=>"010010010",
5869=>"000101101",
5870=>"100010010",
5871=>"101100111",
5872=>"000000111",
5873=>"011111111",
5874=>"011010000",
5875=>"011010000",
5876=>"110011000",
5877=>"101101001",
5878=>"100100001",
5879=>"000101101",
5880=>"000000111",
5881=>"000000111",
5882=>"000100100",
5883=>"111001000",
5884=>"101000000",
5885=>"001000000",
5886=>"101111111",
5887=>"001001101",
5888=>"000001000",
5889=>"000011001",
5890=>"110100101",
5891=>"010011101",
5892=>"000001000",
5893=>"110110010",
5894=>"001011111",
5895=>"110110111",
5896=>"110100100",
5897=>"100100000",
5898=>"000110100",
5899=>"000011000",
5900=>"001001011",
5901=>"101111111",
5902=>"000101001",
5903=>"011010111",
5904=>"100100010",
5905=>"100110100",
5906=>"110001100",
5907=>"000000100",
5908=>"010000101",
5909=>"110111011",
5910=>"111011000",
5911=>"100111000",
5912=>"100000000",
5913=>"111001011",
5914=>"010001110",
5915=>"000100100",
5916=>"001101101",
5917=>"100110111",
5918=>"010110111",
5919=>"100000000",
5920=>"000110000",
5921=>"011001001",
5922=>"000011101",
5923=>"010110011",
5924=>"000100000",
5925=>"001011001",
5926=>"100100110",
5927=>"011001011",
5928=>"100100000",
5929=>"010001011",
5930=>"111111011",
5931=>"100001010",
5932=>"000000001",
5933=>"111111110",
5934=>"111001011",
5935=>"101100110",
5936=>"110100100",
5937=>"101111111",
5938=>"011000011",
5939=>"011001111",
5940=>"010110100",
5941=>"000001001",
5942=>"110110100",
5943=>"010000010",
5944=>"001000111",
5945=>"011001001",
5946=>"001001001",
5947=>"100101100",
5948=>"011011011",
5949=>"001011001",
5950=>"001000001",
5951=>"110111000",
5952=>"111001001",
5953=>"000111100",
5954=>"011011111",
5955=>"011100000",
5956=>"011011011",
5957=>"010010001",
5958=>"011111000",
5959=>"100111011",
5960=>"011001001",
5961=>"101100010",
5962=>"010010110",
5963=>"001011011",
5964=>"101001001",
5965=>"000001011",
5966=>"001100101",
5967=>"001001011",
5968=>"001001011",
5969=>"101000000",
5970=>"011001011",
5971=>"011001000",
5972=>"100100100",
5973=>"001000000",
5974=>"110110010",
5975=>"100100100",
5976=>"101000000",
5977=>"001011111",
5978=>"011011011",
5979=>"111111101",
5980=>"111110000",
5981=>"011111010",
5982=>"011011111",
5983=>"100100110",
5984=>"011011011",
5985=>"001111001",
5986=>"001001111",
5987=>"000000000",
5988=>"000001000",
5989=>"001000100",
5990=>"011111001",
5991=>"100100100",
5992=>"110110110",
5993=>"100110110",
5994=>"111111011",
5995=>"010001011",
5996=>"100000010",
5997=>"001111100",
5998=>"001011111",
5999=>"001011111",
6000=>"100100101",
6001=>"000011111",
6002=>"110110100",
6003=>"010000100",
6004=>"011111000",
6005=>"010000011",
6006=>"001000000",
6007=>"111001111",
6008=>"110111110",
6009=>"000000110",
6010=>"110010010",
6011=>"000000000",
6012=>"011001000",
6013=>"100000000",
6014=>"100100000",
6015=>"100100000",
6016=>"011001110",
6017=>"110110000",
6018=>"110100100",
6019=>"011010111",
6020=>"110000111",
6021=>"100110100",
6022=>"011001111",
6023=>"001011001",
6024=>"101111100",
6025=>"011010011",
6026=>"100110000",
6027=>"001000110",
6028=>"100100100",
6029=>"000010111",
6030=>"100010000",
6031=>"001000001",
6032=>"111101000",
6033=>"110100110",
6034=>"100110100",
6035=>"011011011",
6036=>"001001011",
6037=>"110100110",
6038=>"011001111",
6039=>"000001000",
6040=>"010000000",
6041=>"111001111",
6042=>"110110000",
6043=>"110100100",
6044=>"001001001",
6045=>"110100000",
6046=>"010010000",
6047=>"011001001",
6048=>"011111111",
6049=>"100111100",
6050=>"010000001",
6051=>"000011000",
6052=>"000111011",
6053=>"000000000",
6054=>"010000010",
6055=>"011000011",
6056=>"100100110",
6057=>"010000000",
6058=>"111101001",
6059=>"000000011",
6060=>"011001000",
6061=>"001100000",
6062=>"111011001",
6063=>"001001110",
6064=>"000001110",
6065=>"010001001",
6066=>"110010100",
6067=>"000000100",
6068=>"000111000",
6069=>"011011111",
6070=>"011001011",
6071=>"000001011",
6072=>"000000001",
6073=>"011001001",
6074=>"111001000",
6075=>"000100110",
6076=>"001000100",
6077=>"110100000",
6078=>"100100000",
6079=>"110000110",
6080=>"011001011",
6081=>"000001000",
6082=>"000000000",
6083=>"111101100",
6084=>"001011011",
6085=>"000011011",
6086=>"100001101",
6087=>"111001011",
6088=>"111110110",
6089=>"111000000",
6090=>"001001010",
6091=>"110111111",
6092=>"100100100",
6093=>"001000001",
6094=>"100100000",
6095=>"001110101",
6096=>"100100110",
6097=>"101101101",
6098=>"001001011",
6099=>"000000100",
6100=>"000001011",
6101=>"001011000",
6102=>"011001001",
6103=>"110110100",
6104=>"000000100",
6105=>"000100000",
6106=>"001000101",
6107=>"100110110",
6108=>"111100000",
6109=>"011110110",
6110=>"000000011",
6111=>"110000011",
6112=>"000000011",
6113=>"011000001",
6114=>"100100000",
6115=>"001101101",
6116=>"000100100",
6117=>"011011100",
6118=>"001001001",
6119=>"100101111",
6120=>"111100011",
6121=>"110110100",
6122=>"000110000",
6123=>"111001011",
6124=>"011000000",
6125=>"011101011",
6126=>"000110000",
6127=>"001000100",
6128=>"110110111",
6129=>"011011001",
6130=>"011011011",
6131=>"100000000",
6132=>"110111000",
6133=>"000010010",
6134=>"000001100",
6135=>"000001011",
6136=>"011001101",
6137=>"011110110",
6138=>"000000000",
6139=>"110000001",
6140=>"011011011",
6141=>"100110000",
6142=>"111111001",
6143=>"011001111",
6144=>"011001000",
6145=>"100011001",
6146=>"111100100",
6147=>"000011011",
6148=>"111111111",
6149=>"011011000",
6150=>"001000000",
6151=>"011010010",
6152=>"000100011",
6153=>"000000100",
6154=>"001001000",
6155=>"001011011",
6156=>"100100110",
6157=>"000011011",
6158=>"111001001",
6159=>"100100000",
6160=>"011011011",
6161=>"100000000",
6162=>"000011000",
6163=>"011001011",
6164=>"111011100",
6165=>"111100100",
6166=>"110111110",
6167=>"111110000",
6168=>"000000100",
6169=>"111000110",
6170=>"000100100",
6171=>"000001111",
6172=>"111100100",
6173=>"011101110",
6174=>"011111000",
6175=>"110100100",
6176=>"011001011",
6177=>"100111100",
6178=>"000000100",
6179=>"001000100",
6180=>"101111100",
6181=>"001011010",
6182=>"000010111",
6183=>"000011010",
6184=>"111011000",
6185=>"000000000",
6186=>"000011000",
6187=>"100000000",
6188=>"100101111",
6189=>"011001001",
6190=>"111011100",
6191=>"011001000",
6192=>"000000011",
6193=>"001001001",
6194=>"101100000",
6195=>"110110011",
6196=>"011011100",
6197=>"111100111",
6198=>"110011000",
6199=>"110100100",
6200=>"000100111",
6201=>"100100100",
6202=>"000100010",
6203=>"010100000",
6204=>"000110110",
6205=>"000100100",
6206=>"000000000",
6207=>"000011011",
6208=>"101100001",
6209=>"111111000",
6210=>"111100000",
6211=>"011011010",
6212=>"000100100",
6213=>"100000001",
6214=>"110000011",
6215=>"111101000",
6216=>"100001000",
6217=>"010011001",
6218=>"111111111",
6219=>"100100100",
6220=>"111100000",
6221=>"001001100",
6222=>"000111111",
6223=>"101110100",
6224=>"101111101",
6225=>"011100000",
6226=>"101001000",
6227=>"011001000",
6228=>"100100000",
6229=>"000100111",
6230=>"100001000",
6231=>"011011011",
6232=>"110111010",
6233=>"000000000",
6234=>"110000000",
6235=>"011011011",
6236=>"100100100",
6237=>"001000101",
6238=>"111100000",
6239=>"011011001",
6240=>"000011000",
6241=>"000011011",
6242=>"110000100",
6243=>"010110110",
6244=>"000011110",
6245=>"001111010",
6246=>"000011000",
6247=>"100100000",
6248=>"010011011",
6249=>"000001110",
6250=>"000011011",
6251=>"110110000",
6252=>"000101111",
6253=>"101101000",
6254=>"110100000",
6255=>"111111011",
6256=>"000111000",
6257=>"010011001",
6258=>"001100100",
6259=>"000000110",
6260=>"111000011",
6261=>"010000001",
6262=>"011011011",
6263=>"111001000",
6264=>"001001010",
6265=>"000000000",
6266=>"000100111",
6267=>"100100101",
6268=>"111110011",
6269=>"000010000",
6270=>"100100000",
6271=>"011011001",
6272=>"100000000",
6273=>"010110100",
6274=>"011011011",
6275=>"000001001",
6276=>"011011010",
6277=>"001011001",
6278=>"011001100",
6279=>"000011000",
6280=>"000111111",
6281=>"001001000",
6282=>"000001001",
6283=>"110000000",
6284=>"111101111",
6285=>"100100100",
6286=>"100000111",
6287=>"000000101",
6288=>"111100001",
6289=>"111110110",
6290=>"010000011",
6291=>"111111111",
6292=>"000011011",
6293=>"011001011",
6294=>"100100100",
6295=>"110100000",
6296=>"010011000",
6297=>"100111011",
6298=>"111100000",
6299=>"001011000",
6300=>"100100000",
6301=>"000011011",
6302=>"000000010",
6303=>"100100100",
6304=>"111110011",
6305=>"111110001",
6306=>"100100000",
6307=>"010101100",
6308=>"111010100",
6309=>"110101000",
6310=>"001000011",
6311=>"000000000",
6312=>"000000111",
6313=>"000011011",
6314=>"111100100",
6315=>"110000100",
6316=>"110111101",
6317=>"101001000",
6318=>"111000010",
6319=>"001011111",
6320=>"000001000",
6321=>"010011100",
6322=>"100101010",
6323=>"000000000",
6324=>"011000011",
6325=>"111111111",
6326=>"011010010",
6327=>"001011000",
6328=>"100111000",
6329=>"010111100",
6330=>"000011000",
6331=>"000101111",
6332=>"000111000",
6333=>"011011011",
6334=>"010011000",
6335=>"000000000",
6336=>"101000000",
6337=>"110000000",
6338=>"111011011",
6339=>"010011000",
6340=>"000100010",
6341=>"100101100",
6342=>"011000001",
6343=>"111100111",
6344=>"000111011",
6345=>"010100100",
6346=>"100011011",
6347=>"000011011",
6348=>"000011010",
6349=>"100001011",
6350=>"101000100",
6351=>"000011011",
6352=>"000001000",
6353=>"100110010",
6354=>"111010100",
6355=>"111100000",
6356=>"000011111",
6357=>"111110111",
6358=>"111100100",
6359=>"111001001",
6360=>"111110111",
6361=>"000000010",
6362=>"111100111",
6363=>"100000001",
6364=>"110111110",
6365=>"011001011",
6366=>"000100101",
6367=>"011011011",
6368=>"111100101",
6369=>"100100100",
6370=>"000011000",
6371=>"110111111",
6372=>"001000000",
6373=>"000000010",
6374=>"100001000",
6375=>"101100011",
6376=>"011111001",
6377=>"011011111",
6378=>"010011000",
6379=>"100000001",
6380=>"110111111",
6381=>"011010010",
6382=>"000000000",
6383=>"110000000",
6384=>"011011000",
6385=>"010110000",
6386=>"000000000",
6387=>"010111000",
6388=>"011110101",
6389=>"100000101",
6390=>"000000000",
6391=>"000100100",
6392=>"000110110",
6393=>"111011000",
6394=>"011100100",
6395=>"110111011",
6396=>"100100010",
6397=>"000011011",
6398=>"100001000",
6399=>"100000100",
6400=>"100111011",
6401=>"011001110",
6402=>"100100100",
6403=>"110100010",
6404=>"000011010",
6405=>"001001000",
6406=>"000001001",
6407=>"001111110",
6408=>"010110100",
6409=>"001000000",
6410=>"101111100",
6411=>"111110010",
6412=>"100100011",
6413=>"000000000",
6414=>"000100011",
6415=>"011000000",
6416=>"001100100",
6417=>"001100100",
6418=>"000100100",
6419=>"001101110",
6420=>"000011011",
6421=>"100111000",
6422=>"101101100",
6423=>"001101100",
6424=>"011000000",
6425=>"110111000",
6426=>"110010000",
6427=>"101101000",
6428=>"011000001",
6429=>"111100000",
6430=>"011010110",
6431=>"100000001",
6432=>"101110010",
6433=>"000100010",
6434=>"000010010",
6435=>"000010111",
6436=>"110011001",
6437=>"111001000",
6438=>"100000001",
6439=>"011111110",
6440=>"010111111",
6441=>"001000000",
6442=>"001100010",
6443=>"110111100",
6444=>"000000011",
6445=>"101001100",
6446=>"011011011",
6447=>"011110010",
6448=>"011111100",
6449=>"100110001",
6450=>"011010110",
6451=>"010100100",
6452=>"000011011",
6453=>"101011010",
6454=>"001000111",
6455=>"000110011",
6456=>"000010000",
6457=>"100100100",
6458=>"000001000",
6459=>"001100100",
6460=>"110100000",
6461=>"110000011",
6462=>"111110100",
6463=>"100111010",
6464=>"001100100",
6465=>"011011100",
6466=>"011011100",
6467=>"100111101",
6468=>"000100001",
6469=>"001011010",
6470=>"101111111",
6471=>"010100000",
6472=>"111000111",
6473=>"000111111",
6474=>"111011111",
6475=>"001011011",
6476=>"000001111",
6477=>"100010000",
6478=>"100100011",
6479=>"011110110",
6480=>"110111000",
6481=>"001000101",
6482=>"011101001",
6483=>"101111000",
6484=>"011011101",
6485=>"111110001",
6486=>"000011001",
6487=>"001100000",
6488=>"001011011",
6489=>"000000001",
6490=>"111000000",
6491=>"100101001",
6492=>"001001111",
6493=>"000001000",
6494=>"111011110",
6495=>"010010110",
6496=>"110111111",
6497=>"110010011",
6498=>"101101111",
6499=>"100101101",
6500=>"100000000",
6501=>"100000011",
6502=>"010010001",
6503=>"001011110",
6504=>"100100001",
6505=>"011011101",
6506=>"001010000",
6507=>"010010010",
6508=>"000110011",
6509=>"011001000",
6510=>"111100001",
6511=>"001011100",
6512=>"011101001",
6513=>"001110100",
6514=>"000111100",
6515=>"000110011",
6516=>"011100111",
6517=>"000000000",
6518=>"111100100",
6519=>"000011111",
6520=>"011011100",
6521=>"100111100",
6522=>"001100111",
6523=>"100000000",
6524=>"110100000",
6525=>"010000110",
6526=>"010010000",
6527=>"100111001",
6528=>"001000100",
6529=>"000100000",
6530=>"001011110",
6531=>"111100001",
6532=>"110000100",
6533=>"101111111",
6534=>"001011011",
6535=>"000100011",
6536=>"101100001",
6537=>"011000001",
6538=>"011111111",
6539=>"010010101",
6540=>"110110001",
6541=>"100110010",
6542=>"001100000",
6543=>"010000000",
6544=>"000011001",
6545=>"000010010",
6546=>"000000001",
6547=>"010110110",
6548=>"000100000",
6549=>"001100100",
6550=>"000111100",
6551=>"100000001",
6552=>"000001000",
6553=>"100111110",
6554=>"100101101",
6555=>"100100111",
6556=>"110110111",
6557=>"001011111",
6558=>"011001111",
6559=>"110101111",
6560=>"100011011",
6561=>"001110010",
6562=>"100111111",
6563=>"100010110",
6564=>"111111100",
6565=>"111001001",
6566=>"010011000",
6567=>"010110111",
6568=>"001001100",
6569=>"011010110",
6570=>"111100100",
6571=>"000110100",
6572=>"111000001",
6573=>"111101110",
6574=>"001000000",
6575=>"100110011",
6576=>"010000110",
6577=>"110110000",
6578=>"100000001",
6579=>"110100000",
6580=>"111000001",
6581=>"100111001",
6582=>"000000011",
6583=>"011011011",
6584=>"100111111",
6585=>"110100000",
6586=>"001011001",
6587=>"000000001",
6588=>"010001001",
6589=>"101001100",
6590=>"111001011",
6591=>"000100110",
6592=>"000001000",
6593=>"000000100",
6594=>"011011111",
6595=>"110111001",
6596=>"011011010",
6597=>"111010001",
6598=>"001000110",
6599=>"001100001",
6600=>"100010000",
6601=>"001011100",
6602=>"000100110",
6603=>"011011011",
6604=>"100100000",
6605=>"000110111",
6606=>"100000000",
6607=>"100100110",
6608=>"111100001",
6609=>"101101011",
6610=>"001000100",
6611=>"100000001",
6612=>"101001111",
6613=>"000111111",
6614=>"010011111",
6615=>"011001110",
6616=>"011011111",
6617=>"011000010",
6618=>"101100011",
6619=>"111101101",
6620=>"010100111",
6621=>"111001111",
6622=>"001000001",
6623=>"011111111",
6624=>"100001011",
6625=>"100100011",
6626=>"001100011",
6627=>"110010001",
6628=>"000000000",
6629=>"101011111",
6630=>"011111100",
6631=>"100110011",
6632=>"101110111",
6633=>"011001100",
6634=>"011011001",
6635=>"001101101",
6636=>"000000010",
6637=>"010010000",
6638=>"100000100",
6639=>"000100000",
6640=>"000000010",
6641=>"000000011",
6642=>"011010110",
6643=>"000010111",
6644=>"010010000",
6645=>"010000001",
6646=>"000000001",
6647=>"001110110",
6648=>"001100100",
6649=>"010010110",
6650=>"100000001",
6651=>"100101001",
6652=>"111111111",
6653=>"001001101",
6654=>"000001011",
6655=>"010011111",
6656=>"100000111",
6657=>"111111101",
6658=>"111100100",
6659=>"111011000",
6660=>"111100100",
6661=>"111101001",
6662=>"000000000",
6663=>"111001101",
6664=>"111111111",
6665=>"000000001",
6666=>"111111001",
6667=>"000000100",
6668=>"000000000",
6669=>"000010111",
6670=>"000000101",
6671=>"000110000",
6672=>"000110100",
6673=>"111000111",
6674=>"111101101",
6675=>"001111000",
6676=>"100000000",
6677=>"111111101",
6678=>"011011100",
6679=>"111111111",
6680=>"000000001",
6681=>"000000000",
6682=>"111100111",
6683=>"010010001",
6684=>"111011010",
6685=>"000000001",
6686=>"110111111",
6687=>"010000010",
6688=>"000000000",
6689=>"000000000",
6690=>"111111011",
6691=>"111111101",
6692=>"000000010",
6693=>"110001010",
6694=>"110000000",
6695=>"000010110",
6696=>"100010000",
6697=>"000001010",
6698=>"000000000",
6699=>"000000000",
6700=>"100000000",
6701=>"111111100",
6702=>"000001111",
6703=>"101111111",
6704=>"000111111",
6705=>"111110101",
6706=>"000000000",
6707=>"000001001",
6708=>"110000000",
6709=>"111010111",
6710=>"010000001",
6711=>"101101111",
6712=>"101000000",
6713=>"000000111",
6714=>"100101100",
6715=>"011111111",
6716=>"101100001",
6717=>"111111111",
6718=>"010111011",
6719=>"011111011",
6720=>"110110000",
6721=>"010101101",
6722=>"001000000",
6723=>"111101100",
6724=>"000000000",
6725=>"101101111",
6726=>"000000000",
6727=>"000001111",
6728=>"000011111",
6729=>"010000000",
6730=>"000000101",
6731=>"111111001",
6732=>"111000101",
6733=>"010110100",
6734=>"010011111",
6735=>"111100101",
6736=>"000101101",
6737=>"111111101",
6738=>"010110010",
6739=>"001000000",
6740=>"111111010",
6741=>"000100100",
6742=>"010010100",
6743=>"100100011",
6744=>"001001010",
6745=>"000000000",
6746=>"000111010",
6747=>"001001001",
6748=>"010111111",
6749=>"110110000",
6750=>"000000111",
6751=>"110001011",
6752=>"000000000",
6753=>"110111011",
6754=>"110110100",
6755=>"110111101",
6756=>"001000000",
6757=>"010011011",
6758=>"000000111",
6759=>"000000001",
6760=>"000111000",
6761=>"010011010",
6762=>"011110111",
6763=>"000000111",
6764=>"101001101",
6765=>"111111111",
6766=>"000000101",
6767=>"110010000",
6768=>"010110111",
6769=>"100010100",
6770=>"011000010",
6771=>"000000011",
6772=>"000110111",
6773=>"000000100",
6774=>"111000000",
6775=>"100000010",
6776=>"101010010",
6777=>"001000011",
6778=>"000011000",
6779=>"101111110",
6780=>"011001001",
6781=>"001001011",
6782=>"000000000",
6783=>"111111111",
6784=>"000100100",
6785=>"000011000",
6786=>"011111110",
6787=>"000001001",
6788=>"000100000",
6789=>"111111110",
6790=>"110101100",
6791=>"000000000",
6792=>"010111011",
6793=>"001000000",
6794=>"111010011",
6795=>"000101111",
6796=>"000111111",
6797=>"111111010",
6798=>"111010110",
6799=>"000111000",
6800=>"000100100",
6801=>"111011000",
6802=>"000001111",
6803=>"000011000",
6804=>"100000000",
6805=>"111000000",
6806=>"111111010",
6807=>"110110100",
6808=>"010011000",
6809=>"101111101",
6810=>"110111000",
6811=>"011010000",
6812=>"001000000",
6813=>"110111010",
6814=>"010010000",
6815=>"111001001",
6816=>"011001001",
6817=>"111010111",
6818=>"000000111",
6819=>"101011111",
6820=>"000111011",
6821=>"110100100",
6822=>"000000100",
6823=>"000100101",
6824=>"111110110",
6825=>"111111101",
6826=>"111111111",
6827=>"111000000",
6828=>"111101001",
6829=>"000111101",
6830=>"110100111",
6831=>"100011111",
6832=>"001101000",
6833=>"100110110",
6834=>"011011001",
6835=>"100100000",
6836=>"111101011",
6837=>"111101101",
6838=>"000000000",
6839=>"011011000",
6840=>"101001101",
6841=>"000000000",
6842=>"001010000",
6843=>"010000110",
6844=>"001100000",
6845=>"101000010",
6846=>"011111010",
6847=>"000000000",
6848=>"100100110",
6849=>"010111111",
6850=>"000000000",
6851=>"011001001",
6852=>"001001101",
6853=>"000010101",
6854=>"001000000",
6855=>"000000111",
6856=>"001101101",
6857=>"101000100",
6858=>"000001000",
6859=>"000001100",
6860=>"011010011",
6861=>"110100100",
6862=>"000111010",
6863=>"100101110",
6864=>"111000111",
6865=>"001011010",
6866=>"000000000",
6867=>"101000010",
6868=>"011110000",
6869=>"001011010",
6870=>"000000001",
6871=>"111111000",
6872=>"011111111",
6873=>"000010001",
6874=>"101100100",
6875=>"111111011",
6876=>"100110000",
6877=>"101100101",
6878=>"000000000",
6879=>"110110000",
6880=>"001000000",
6881=>"000111111",
6882=>"000000110",
6883=>"111111111",
6884=>"000000111",
6885=>"001000000",
6886=>"001111110",
6887=>"010011111",
6888=>"011111010",
6889=>"000000000",
6890=>"011111100",
6891=>"111101111",
6892=>"100000000",
6893=>"000010100",
6894=>"101001000",
6895=>"111111111",
6896=>"111111000",
6897=>"000000100",
6898=>"100100111",
6899=>"100000000",
6900=>"001011001",
6901=>"100111110",
6902=>"101101101",
6903=>"000010011",
6904=>"000000000",
6905=>"000111111",
6906=>"000000000",
6907=>"100000000",
6908=>"110111010",
6909=>"011111111",
6910=>"011011011",
6911=>"000101111",
6912=>"101001001",
6913=>"011010100",
6914=>"111000001",
6915=>"000111000",
6916=>"111111111",
6917=>"001111101",
6918=>"110111110",
6919=>"011010111",
6920=>"000000111",
6921=>"011111110",
6922=>"011000000",
6923=>"010000000",
6924=>"001000100",
6925=>"001110001",
6926=>"000000100",
6927=>"100001001",
6928=>"101100100",
6929=>"111001011",
6930=>"100000000",
6931=>"110001100",
6932=>"110011011",
6933=>"110011111",
6934=>"101101001",
6935=>"001111111",
6936=>"111010111",
6937=>"000100100",
6938=>"111111100",
6939=>"110011000",
6940=>"111011001",
6941=>"111010000",
6942=>"011011000",
6943=>"100000000",
6944=>"111011011",
6945=>"111111100",
6946=>"110111111",
6947=>"111111100",
6948=>"000101011",
6949=>"111000000",
6950=>"001001111",
6951=>"011100110",
6952=>"110000011",
6953=>"110111000",
6954=>"001001101",
6955=>"100011110",
6956=>"100101011",
6957=>"111000010",
6958=>"111111011",
6959=>"010111000",
6960=>"100111001",
6961=>"001000110",
6962=>"101100111",
6963=>"101111100",
6964=>"011001000",
6965=>"001011010",
6966=>"001011001",
6967=>"000101111",
6968=>"110111101",
6969=>"000001001",
6970=>"100010011",
6971=>"111011101",
6972=>"100100000",
6973=>"000001001",
6974=>"100000000",
6975=>"010000110",
6976=>"110100100",
6977=>"000011001",
6978=>"101111111",
6979=>"001001011",
6980=>"000000000",
6981=>"110100000",
6982=>"011001110",
6983=>"100111111",
6984=>"110111111",
6985=>"011111100",
6986=>"000001001",
6987=>"001010100",
6988=>"101101000",
6989=>"101101000",
6990=>"100111111",
6991=>"100000000",
6992=>"000100000",
6993=>"000100100",
6994=>"001011011",
6995=>"111011000",
6996=>"101110000",
6997=>"100000011",
6998=>"100111100",
6999=>"001001000",
7000=>"000100110",
7001=>"100010010",
7002=>"111011000",
7003=>"101100110",
7004=>"000111011",
7005=>"110010001",
7006=>"111000111",
7007=>"011001000",
7008=>"011000111",
7009=>"110100000",
7010=>"001000111",
7011=>"101111011",
7012=>"000000000",
7013=>"100110011",
7014=>"100100100",
7015=>"000010000",
7016=>"010000010",
7017=>"111001001",
7018=>"111011110",
7019=>"000110100",
7020=>"111011111",
7021=>"111011001",
7022=>"011011101",
7023=>"010110110",
7024=>"001110000",
7025=>"001000100",
7026=>"000000001",
7027=>"101100110",
7028=>"111111010",
7029=>"001011111",
7030=>"011000101",
7031=>"111011111",
7032=>"110001000",
7033=>"000111110",
7034=>"100100110",
7035=>"010011101",
7036=>"000100100",
7037=>"110000010",
7038=>"011011111",
7039=>"111011001",
7040=>"100001111",
7041=>"100000001",
7042=>"110011011",
7043=>"110111011",
7044=>"000000110",
7045=>"001101000",
7046=>"100011011",
7047=>"000100000",
7048=>"000101101",
7049=>"110100000",
7050=>"100000011",
7051=>"101111000",
7052=>"001100111",
7053=>"101011111",
7054=>"000010110",
7055=>"001010000",
7056=>"111110000",
7057=>"001011000",
7058=>"110101001",
7059=>"100110110",
7060=>"000100110",
7061=>"001001000",
7062=>"100100100",
7063=>"111001000",
7064=>"110110011",
7065=>"111001111",
7066=>"011111011",
7067=>"011000001",
7068=>"000001000",
7069=>"000100010",
7070=>"010011000",
7071=>"000000000",
7072=>"011001100",
7073=>"000001011",
7074=>"111111001",
7075=>"000100110",
7076=>"000101001",
7077=>"100100000",
7078=>"010010101",
7079=>"000000001",
7080=>"101111000",
7081=>"100000000",
7082=>"110000000",
7083=>"100001001",
7084=>"110110000",
7085=>"000010101",
7086=>"110011000",
7087=>"000100100",
7088=>"110000110",
7089=>"001111111",
7090=>"001011110",
7091=>"000100100",
7092=>"101000011",
7093=>"010011110",
7094=>"100100000",
7095=>"100000000",
7096=>"110110000",
7097=>"000110110",
7098=>"100101001",
7099=>"101111011",
7100=>"111010000",
7101=>"000001111",
7102=>"011001111",
7103=>"100100110",
7104=>"000100000",
7105=>"000000111",
7106=>"011001010",
7107=>"111111000",
7108=>"000000011",
7109=>"111100001",
7110=>"000001001",
7111=>"001010011",
7112=>"111011110",
7113=>"111000001",
7114=>"101000111",
7115=>"110000111",
7116=>"010000001",
7117=>"000110110",
7118=>"110111000",
7119=>"101100000",
7120=>"011011001",
7121=>"000100101",
7122=>"001110110",
7123=>"100000111",
7124=>"001000111",
7125=>"110111011",
7126=>"011000000",
7127=>"011011011",
7128=>"000000101",
7129=>"100000000",
7130=>"100000111",
7131=>"001001111",
7132=>"110111000",
7133=>"010000100",
7134=>"000100000",
7135=>"001100101",
7136=>"000011111",
7137=>"001001100",
7138=>"001111111",
7139=>"111111111",
7140=>"010000000",
7141=>"011111111",
7142=>"011001001",
7143=>"010101111",
7144=>"101000000",
7145=>"010000000",
7146=>"011001001",
7147=>"100001100",
7148=>"101000100",
7149=>"110110000",
7150=>"000100000",
7151=>"011001001",
7152=>"110001000",
7153=>"110001010",
7154=>"010111000",
7155=>"010001011",
7156=>"001111000",
7157=>"011001001",
7158=>"111011000",
7159=>"011110000",
7160=>"001111110",
7161=>"011001111",
7162=>"100000000",
7163=>"010110000",
7164=>"000111000",
7165=>"000010011",
7166=>"110110000",
7167=>"000000000",
7168=>"001001001",
7169=>"110000011",
7170=>"000010000",
7171=>"011101000",
7172=>"100011100",
7173=>"100000111",
7174=>"010111111",
7175=>"111111110",
7176=>"011101100",
7177=>"111110100",
7178=>"101000000",
7179=>"101000001",
7180=>"010011110",
7181=>"000000110",
7182=>"100000100",
7183=>"111111111",
7184=>"000000000",
7185=>"000000010",
7186=>"111001000",
7187=>"000101011",
7188=>"111111000",
7189=>"111101111",
7190=>"011101011",
7191=>"110111111",
7192=>"100000000",
7193=>"111111011",
7194=>"000000101",
7195=>"000000000",
7196=>"000000000",
7197=>"000000000",
7198=>"101000000",
7199=>"111001000",
7200=>"000000010",
7201=>"111010001",
7202=>"101000100",
7203=>"111101100",
7204=>"100001100",
7205=>"001000000",
7206=>"000000001",
7207=>"110001100",
7208=>"000000101",
7209=>"100000000",
7210=>"100101110",
7211=>"000000000",
7212=>"111100001",
7213=>"000001010",
7214=>"010010111",
7215=>"111111111",
7216=>"111000000",
7217=>"000000000",
7218=>"111110111",
7219=>"001010010",
7220=>"000000000",
7221=>"000000000",
7222=>"000000011",
7223=>"111111100",
7224=>"111111111",
7225=>"000000000",
7226=>"000000100",
7227=>"111000000",
7228=>"111000000",
7229=>"111111111",
7230=>"000000000",
7231=>"100100100",
7232=>"111111110",
7233=>"001000000",
7234=>"000000000",
7235=>"011011111",
7236=>"100000111",
7237=>"111001110",
7238=>"001010111",
7239=>"000000111",
7240=>"000000011",
7241=>"100000001",
7242=>"101011111",
7243=>"111111111",
7244=>"000000111",
7245=>"111100001",
7246=>"111001001",
7247=>"011000000",
7248=>"000000000",
7249=>"111111111",
7250=>"111100110",
7251=>"001000000",
7252=>"000101001",
7253=>"000100110",
7254=>"011000000",
7255=>"000000000",
7256=>"000001000",
7257=>"000100000",
7258=>"010010010",
7259=>"111011101",
7260=>"011111111",
7261=>"110000001",
7262=>"011111110",
7263=>"100100000",
7264=>"000000000",
7265=>"000100000",
7266=>"110111000",
7267=>"011011000",
7268=>"010100100",
7269=>"111011100",
7270=>"000001110",
7271=>"111110000",
7272=>"111011000",
7273=>"110000000",
7274=>"000001111",
7275=>"111001111",
7276=>"000010111",
7277=>"100000011",
7278=>"111110001",
7279=>"000001000",
7280=>"000100100",
7281=>"111001001",
7282=>"001000110",
7283=>"101000100",
7284=>"000000101",
7285=>"000000111",
7286=>"111100101",
7287=>"000010010",
7288=>"010110110",
7289=>"000000010",
7290=>"101111111",
7291=>"000111111",
7292=>"001100010",
7293=>"100100100",
7294=>"111011000",
7295=>"000001001",
7296=>"101010010",
7297=>"111000000",
7298=>"000111000",
7299=>"110110111",
7300=>"000000000",
7301=>"010101100",
7302=>"000000001",
7303=>"011001001",
7304=>"000111111",
7305=>"101000010",
7306=>"110000101",
7307=>"100000111",
7308=>"010010000",
7309=>"100000000",
7310=>"010111111",
7311=>"000000000",
7312=>"101111100",
7313=>"000000011",
7314=>"000000010",
7315=>"001011011",
7316=>"110000001",
7317=>"010000000",
7318=>"110111111",
7319=>"110101001",
7320=>"100001010",
7321=>"000010100",
7322=>"000100100",
7323=>"000010010",
7324=>"000001011",
7325=>"000000000",
7326=>"111000011",
7327=>"111001111",
7328=>"000100101",
7329=>"000000010",
7330=>"111111111",
7331=>"110110111",
7332=>"000000111",
7333=>"001101111",
7334=>"011010000",
7335=>"000000111",
7336=>"111000110",
7337=>"100110010",
7338=>"101000000",
7339=>"010000000",
7340=>"111110111",
7341=>"000000000",
7342=>"000100100",
7343=>"110111111",
7344=>"111111111",
7345=>"100000010",
7346=>"011011011",
7347=>"001000100",
7348=>"010001000",
7349=>"111111111",
7350=>"000000100",
7351=>"010111100",
7352=>"101100000",
7353=>"011000110",
7354=>"000000000",
7355=>"000100111",
7356=>"100000000",
7357=>"000000000",
7358=>"111111010",
7359=>"011010111",
7360=>"000111101",
7361=>"000000000",
7362=>"001111111",
7363=>"001001111",
7364=>"100000110",
7365=>"001100000",
7366=>"100000011",
7367=>"011011011",
7368=>"000000000",
7369=>"101000111",
7370=>"010000110",
7371=>"111101000",
7372=>"111000010",
7373=>"100001010",
7374=>"000000010",
7375=>"000000010",
7376=>"101101101",
7377=>"001001100",
7378=>"101000011",
7379=>"111111111",
7380=>"011111011",
7381=>"100100100",
7382=>"000000100",
7383=>"110010000",
7384=>"111111111",
7385=>"111100110",
7386=>"101111111",
7387=>"111000000",
7388=>"000001011",
7389=>"101110011",
7390=>"111101100",
7391=>"111101110",
7392=>"111010011",
7393=>"111111111",
7394=>"000001111",
7395=>"011110000",
7396=>"000000000",
7397=>"101110111",
7398=>"100110000",
7399=>"010011100",
7400=>"000000000",
7401=>"000010010",
7402=>"100000010",
7403=>"000010001",
7404=>"101000000",
7405=>"000000000",
7406=>"111000001",
7407=>"000000111",
7408=>"000001000",
7409=>"000001100",
7410=>"000001110",
7411=>"001001010",
7412=>"100000100",
7413=>"111101110",
7414=>"000000000",
7415=>"000010111",
7416=>"011011000",
7417=>"111011001",
7418=>"111111111",
7419=>"110100000",
7420=>"011001111",
7421=>"100110000",
7422=>"000000001",
7423=>"000100110",
7424=>"100000100",
7425=>"110011101",
7426=>"011010101",
7427=>"101001111",
7428=>"000100111",
7429=>"110100100",
7430=>"111000000",
7431=>"011000101",
7432=>"111001001",
7433=>"000000010",
7434=>"110110000",
7435=>"110101110",
7436=>"001000111",
7437=>"111000010",
7438=>"110101010",
7439=>"110010001",
7440=>"101101000",
7441=>"011010000",
7442=>"111110111",
7443=>"000000000",
7444=>"101101000",
7445=>"010011011",
7446=>"011011111",
7447=>"110111000",
7448=>"010000110",
7449=>"000101001",
7450=>"011000110",
7451=>"000111000",
7452=>"000100100",
7453=>"000000111",
7454=>"000000111",
7455=>"000000111",
7456=>"010000010",
7457=>"000101011",
7458=>"000000010",
7459=>"001101000",
7460=>"111111111",
7461=>"100001001",
7462=>"110110000",
7463=>"101011000",
7464=>"001001111",
7465=>"011001001",
7466=>"111001000",
7467=>"010111011",
7468=>"000111010",
7469=>"111110000",
7470=>"101111010",
7471=>"001111111",
7472=>"011010000",
7473=>"111111110",
7474=>"101001101",
7475=>"111111000",
7476=>"011010010",
7477=>"010011001",
7478=>"010011011",
7479=>"010000110",
7480=>"101000111",
7481=>"101100111",
7482=>"000000111",
7483=>"111111000",
7484=>"110111010",
7485=>"000111111",
7486=>"000000101",
7487=>"111111110",
7488=>"011000000",
7489=>"000000100",
7490=>"011010000",
7491=>"100101001",
7492=>"000000000",
7493=>"010010100",
7494=>"001001111",
7495=>"000111110",
7496=>"100101111",
7497=>"111100111",
7498=>"101100111",
7499=>"000111111",
7500=>"000100101",
7501=>"111110000",
7502=>"110010111",
7503=>"111111000",
7504=>"000000111",
7505=>"111111101",
7506=>"101001111",
7507=>"011101000",
7508=>"111110111",
7509=>"100100011",
7510=>"110110011",
7511=>"101100001",
7512=>"000100011",
7513=>"000001000",
7514=>"000000000",
7515=>"000000011",
7516=>"000000110",
7517=>"001000111",
7518=>"100111001",
7519=>"001100110",
7520=>"011101000",
7521=>"000100111",
7522=>"101000111",
7523=>"110100000",
7524=>"111000111",
7525=>"110110111",
7526=>"100000110",
7527=>"111111010",
7528=>"000000000",
7529=>"000000010",
7530=>"000000000",
7531=>"111000111",
7532=>"010111011",
7533=>"000010010",
7534=>"111100111",
7535=>"011010000",
7536=>"011110111",
7537=>"000000000",
7538=>"000010110",
7539=>"111000100",
7540=>"000000000",
7541=>"011000001",
7542=>"000000000",
7543=>"111010101",
7544=>"000000000",
7545=>"000010111",
7546=>"000000000",
7547=>"111111110",
7548=>"011101001",
7549=>"010000000",
7550=>"111111010",
7551=>"100100111",
7552=>"111101000",
7553=>"110000011",
7554=>"000000101",
7555=>"000011011",
7556=>"000000110",
7557=>"010111110",
7558=>"001000000",
7559=>"000000100",
7560=>"111011010",
7561=>"010110100",
7562=>"010000010",
7563=>"110010111",
7564=>"111011001",
7565=>"101011000",
7566=>"000000100",
7567=>"000110000",
7568=>"101111100",
7569=>"011011110",
7570=>"000000101",
7571=>"011111111",
7572=>"100000001",
7573=>"000000110",
7574=>"111101100",
7575=>"101100110",
7576=>"000001101",
7577=>"000000101",
7578=>"100100101",
7579=>"110010110",
7580=>"111100111",
7581=>"000100101",
7582=>"000000000",
7583=>"111010010",
7584=>"111001000",
7585=>"111111000",
7586=>"111111010",
7587=>"000111111",
7588=>"000000100",
7589=>"110100010",
7590=>"010011101",
7591=>"001000000",
7592=>"110111010",
7593=>"001111101",
7594=>"111100111",
7595=>"011000001",
7596=>"001101101",
7597=>"100101111",
7598=>"001000011",
7599=>"110100111",
7600=>"110101101",
7601=>"000001111",
7602=>"111100011",
7603=>"000001011",
7604=>"110110000",
7605=>"110111010",
7606=>"001100111",
7607=>"000000001",
7608=>"100110110",
7609=>"001001101",
7610=>"110010100",
7611=>"101001111",
7612=>"001000101",
7613=>"101000001",
7614=>"000100111",
7615=>"111010000",
7616=>"010010000",
7617=>"100000001",
7618=>"000000110",
7619=>"111110111",
7620=>"101001000",
7621=>"011000111",
7622=>"000100111",
7623=>"110110111",
7624=>"111101111",
7625=>"111010000",
7626=>"100000001",
7627=>"100000100",
7628=>"011000000",
7629=>"000100100",
7630=>"000000000",
7631=>"000101111",
7632=>"010000000",
7633=>"011011000",
7634=>"100101111",
7635=>"111111110",
7636=>"000000011",
7637=>"000111101",
7638=>"111000000",
7639=>"001001111",
7640=>"111111000",
7641=>"101000011",
7642=>"110110000",
7643=>"000000100",
7644=>"011011010",
7645=>"101101111",
7646=>"111111100",
7647=>"101000111",
7648=>"010111010",
7649=>"000010111",
7650=>"100000111",
7651=>"111011010",
7652=>"001000001",
7653=>"100101111",
7654=>"110000111",
7655=>"000010111",
7656=>"000000111",
7657=>"011111001",
7658=>"011010010",
7659=>"000000101",
7660=>"101101001",
7661=>"011111101",
7662=>"101001010",
7663=>"010110011",
7664=>"000010000",
7665=>"010001001",
7666=>"000000110",
7667=>"010011000",
7668=>"001000010",
7669=>"000111000",
7670=>"000100100",
7671=>"000011000",
7672=>"000000000",
7673=>"111011000",
7674=>"100000100",
7675=>"011001001",
7676=>"111111111",
7677=>"000000000",
7678=>"110010011",
7679=>"111000010",
7680=>"011001100",
7681=>"011011011",
7682=>"100100011",
7683=>"000010011",
7684=>"111011111",
7685=>"000000000",
7686=>"011011011",
7687=>"011011011",
7688=>"000000000",
7689=>"110100110",
7690=>"000001011",
7691=>"111011110",
7692=>"000100110",
7693=>"100100100",
7694=>"100000001",
7695=>"001001101",
7696=>"000001011",
7697=>"001001000",
7698=>"100100110",
7699=>"000001001",
7700=>"001011111",
7701=>"110100110",
7702=>"001001001",
7703=>"001001001",
7704=>"000000001",
7705=>"011000000",
7706=>"001010111",
7707=>"000000000",
7708=>"011111011",
7709=>"110110010",
7710=>"001011110",
7711=>"000100000",
7712=>"000001100",
7713=>"001101101",
7714=>"111101010",
7715=>"000100111",
7716=>"111110110",
7717=>"101111011",
7718=>"110010010",
7719=>"101001000",
7720=>"000110101",
7721=>"000100100",
7722=>"001001011",
7723=>"100100011",
7724=>"111110011",
7725=>"001011101",
7726=>"010000000",
7727=>"001000000",
7728=>"001001100",
7729=>"011111110",
7730=>"001000000",
7731=>"001111001",
7732=>"000000111",
7733=>"110011000",
7734=>"100000000",
7735=>"010000001",
7736=>"000110000",
7737=>"001000100",
7738=>"110110111",
7739=>"001001001",
7740=>"000000000",
7741=>"111110010",
7742=>"000100110",
7743=>"110001100",
7744=>"111101101",
7745=>"111110110",
7746=>"100100000",
7747=>"000010000",
7748=>"100100100",
7749=>"001000000",
7750=>"011001001",
7751=>"100110001",
7752=>"011010000",
7753=>"001111111",
7754=>"001000100",
7755=>"000000000",
7756=>"000001011",
7757=>"110110001",
7758=>"110010101",
7759=>"110001011",
7760=>"110000000",
7761=>"111110111",
7762=>"000100001",
7763=>"101100000",
7764=>"110001001",
7765=>"011001000",
7766=>"010110100",
7767=>"100100111",
7768=>"001001110",
7769=>"001011010",
7770=>"011011110",
7771=>"110100000",
7772=>"100011011",
7773=>"000100011",
7774=>"101101111",
7775=>"100100100",
7776=>"010010010",
7777=>"010110011",
7778=>"100100101",
7779=>"111011101",
7780=>"001010010",
7781=>"101010001",
7782=>"111011110",
7783=>"110110100",
7784=>"001111110",
7785=>"001011101",
7786=>"001101101",
7787=>"100110000",
7788=>"000111111",
7789=>"001011110",
7790=>"011000011",
7791=>"101111001",
7792=>"001010010",
7793=>"001001100",
7794=>"110100000",
7795=>"000100000",
7796=>"000100100",
7797=>"010000110",
7798=>"110110101",
7799=>"000000001",
7800=>"011011111",
7801=>"001001011",
7802=>"001001001",
7803=>"000010000",
7804=>"110100101",
7805=>"110000000",
7806=>"001001001",
7807=>"110100100",
7808=>"100001111",
7809=>"010011000",
7810=>"100001001",
7811=>"110100111",
7812=>"001001001",
7813=>"111110100",
7814=>"101101000",
7815=>"000000000",
7816=>"000010111",
7817=>"000000100",
7818=>"010001000",
7819=>"000000111",
7820=>"000010010",
7821=>"110110111",
7822=>"010011101",
7823=>"100100000",
7824=>"000100100",
7825=>"011010011",
7826=>"000001000",
7827=>"010110100",
7828=>"000001001",
7829=>"000000001",
7830=>"100011111",
7831=>"101111100",
7832=>"100111110",
7833=>"011001011",
7834=>"100111111",
7835=>"100100110",
7836=>"101110010",
7837=>"000001101",
7838=>"001011100",
7839=>"110111011",
7840=>"010010100",
7841=>"001010110",
7842=>"110100011",
7843=>"101100011",
7844=>"011001001",
7845=>"111111101",
7846=>"001001001",
7847=>"101001000",
7848=>"011001001",
7849=>"001001010",
7850=>"100100100",
7851=>"000000000",
7852=>"000000001",
7853=>"100000000",
7854=>"000000110",
7855=>"001110000",
7856=>"100100000",
7857=>"111111101",
7858=>"000011011",
7859=>"111110100",
7860=>"011011100",
7861=>"110011001",
7862=>"011110110",
7863=>"100100111",
7864=>"110011010",
7865=>"101111101",
7866=>"001101101",
7867=>"001011111",
7868=>"001010111",
7869=>"010110111",
7870=>"010110110",
7871=>"001010101",
7872=>"010110010",
7873=>"010000000",
7874=>"010111000",
7875=>"110110110",
7876=>"001001111",
7877=>"111011110",
7878=>"000001001",
7879=>"010000010",
7880=>"011011000",
7881=>"110000000",
7882=>"110110100",
7883=>"000111110",
7884=>"001000111",
7885=>"000110111",
7886=>"010000110",
7887=>"000000100",
7888=>"100100100",
7889=>"101110000",
7890=>"111010100",
7891=>"001001101",
7892=>"100100111",
7893=>"000000011",
7894=>"000100100",
7895=>"001001100",
7896=>"011011010",
7897=>"001100001",
7898=>"000000100",
7899=>"001001001",
7900=>"000100011",
7901=>"000001010",
7902=>"001000010",
7903=>"001001001",
7904=>"000100000",
7905=>"100100111",
7906=>"101011111",
7907=>"111110000",
7908=>"000000000",
7909=>"110110110",
7910=>"110010110",
7911=>"110110001",
7912=>"110101011",
7913=>"011011011",
7914=>"111101100",
7915=>"011001011",
7916=>"000100100",
7917=>"110000010",
7918=>"010110011",
7919=>"000000011",
7920=>"101000001",
7921=>"100001000",
7922=>"001001001",
7923=>"101001101",
7924=>"000011011",
7925=>"011011001",
7926=>"100000001",
7927=>"001000001",
7928=>"001001001",
7929=>"111100000",
7930=>"111110110",
7931=>"001110000",
7932=>"110000011",
7933=>"100100110",
7934=>"000000000",
7935=>"010110001",
7936=>"000000001",
7937=>"100000011",
7938=>"101010010",
7939=>"011010011",
7940=>"011101011",
7941=>"011001000",
7942=>"000000010",
7943=>"000000111",
7944=>"101101000",
7945=>"000000000",
7946=>"001001011",
7947=>"101011101",
7948=>"100000000",
7949=>"100100000",
7950=>"000101001",
7951=>"000000011",
7952=>"000000111",
7953=>"110110010",
7954=>"111011000",
7955=>"010101000",
7956=>"111010001",
7957=>"100100111",
7958=>"101111110",
7959=>"000010010",
7960=>"111000001",
7961=>"011101000",
7962=>"000011101",
7963=>"000100100",
7964=>"111000101",
7965=>"110101111",
7966=>"110111000",
7967=>"111100101",
7968=>"111000000",
7969=>"010010010",
7970=>"000000010",
7971=>"011011010",
7972=>"100100000",
7973=>"110100000",
7974=>"000101000",
7975=>"000000010",
7976=>"010111000",
7977=>"010000111",
7978=>"000000111",
7979=>"111000000",
7980=>"000001011",
7981=>"010011000",
7982=>"011101001",
7983=>"000001000",
7984=>"010110000",
7985=>"000100100",
7986=>"000010000",
7987=>"010011011",
7988=>"000100100",
7989=>"101000001",
7990=>"100110100",
7991=>"111000001",
7992=>"000011111",
7993=>"101000000",
7994=>"111000000",
7995=>"110111001",
7996=>"011101001",
7997=>"001100101",
7998=>"000000010",
7999=>"000100001",
8000=>"001111100",
8001=>"111111000",
8002=>"011111111",
8003=>"001000101",
8004=>"111001000",
8005=>"111111010",
8006=>"000100111",
8007=>"110111010",
8008=>"000100110",
8009=>"000110111",
8010=>"110000000",
8011=>"000000000",
8012=>"000110000",
8013=>"001001100",
8014=>"110001100",
8015=>"111000110",
8016=>"000000010",
8017=>"010110110",
8018=>"000111010",
8019=>"011001100",
8020=>"001111100",
8021=>"001101110",
8022=>"000011100",
8023=>"110111111",
8024=>"011001001",
8025=>"010110110",
8026=>"011011100",
8027=>"000000111",
8028=>"101001000",
8029=>"110111001",
8030=>"000111111",
8031=>"100100100",
8032=>"010000101",
8033=>"000010010",
8034=>"111111111",
8035=>"110110011",
8036=>"001000101",
8037=>"110100000",
8038=>"110110001",
8039=>"111111001",
8040=>"001101100",
8041=>"000011010",
8042=>"010111100",
8043=>"000000000",
8044=>"011010000",
8045=>"000010010",
8046=>"100000100",
8047=>"000000000",
8048=>"111001001",
8049=>"111111011",
8050=>"000001001",
8051=>"111000000",
8052=>"011011101",
8053=>"101000100",
8054=>"000000001",
8055=>"000111111",
8056=>"111110111",
8057=>"000101000",
8058=>"110000110",
8059=>"001010000",
8060=>"000110111",
8061=>"100100000",
8062=>"011110000",
8063=>"101000000",
8064=>"001100111",
8065=>"111111001",
8066=>"000111111",
8067=>"011111111",
8068=>"000001000",
8069=>"000110111",
8070=>"011011001",
8071=>"000000110",
8072=>"101100100",
8073=>"000111011",
8074=>"111010000",
8075=>"111011010",
8076=>"101000000",
8077=>"101010000",
8078=>"001111011",
8079=>"011001011",
8080=>"000001001",
8081=>"100101100",
8082=>"000110001",
8083=>"110001010",
8084=>"000000011",
8085=>"010111110",
8086=>"001100010",
8087=>"000100001",
8088=>"111010110",
8089=>"001000110",
8090=>"001111000",
8091=>"100100111",
8092=>"011111111",
8093=>"100010011",
8094=>"011111001",
8095=>"010101111",
8096=>"100100010",
8097=>"111010010",
8098=>"000101101",
8099=>"000000010",
8100=>"110111101",
8101=>"000001001",
8102=>"001100000",
8103=>"100100000",
8104=>"111111110",
8105=>"101111111",
8106=>"000000101",
8107=>"000010000",
8108=>"111111111",
8109=>"000111111",
8110=>"111001000",
8111=>"000111111",
8112=>"111111000",
8113=>"110110000",
8114=>"111101011",
8115=>"000001001",
8116=>"110110110",
8117=>"000010010",
8118=>"001101100",
8119=>"101011010",
8120=>"010100100",
8121=>"100000110",
8122=>"100101010",
8123=>"111111000",
8124=>"000000010",
8125=>"000011100",
8126=>"100110100",
8127=>"000010111",
8128=>"011000000",
8129=>"000001110",
8130=>"011111111",
8131=>"001100100",
8132=>"000010000",
8133=>"001000111",
8134=>"000110100",
8135=>"100000011",
8136=>"111111111",
8137=>"111000001",
8138=>"011000000",
8139=>"101111111",
8140=>"001000111",
8141=>"001011111",
8142=>"100100110",
8143=>"000110111",
8144=>"000011000",
8145=>"001001001",
8146=>"111111010",
8147=>"100001001",
8148=>"000101111",
8149=>"011001000",
8150=>"101000011",
8151=>"111111110",
8152=>"100101001",
8153=>"010101000",
8154=>"001001000",
8155=>"000000010",
8156=>"100101011",
8157=>"101000111",
8158=>"000110111",
8159=>"111111111",
8160=>"000101111",
8161=>"111001100",
8162=>"000001111",
8163=>"011001001",
8164=>"010100000",
8165=>"111111101",
8166=>"101111000",
8167=>"001000000",
8168=>"111000000",
8169=>"111000011",
8170=>"100110110",
8171=>"000101101",
8172=>"000000000",
8173=>"111100111",
8174=>"010000000",
8175=>"100000011",
8176=>"100101100",
8177=>"000001001",
8178=>"111011000",
8179=>"011001001",
8180=>"100100001",
8181=>"000000001",
8182=>"000000111",
8183=>"000111100",
8184=>"001001011",
8185=>"000100010",
8186=>"010111111",
8187=>"000000111",
8188=>"101111111",
8189=>"101111010",
8190=>"110110000",
8191=>"001011011",
8192=>"111111100",
8193=>"000011001",
8194=>"101000101",
8195=>"000000111",
8196=>"001001011",
8197=>"001000000",
8198=>"111111111",
8199=>"111101101",
8200=>"010011001",
8201=>"110100000",
8202=>"000000110",
8203=>"101111101",
8204=>"000011000",
8205=>"011000011",
8206=>"100010011",
8207=>"110000010",
8208=>"011000000",
8209=>"101000101",
8210=>"100000100",
8211=>"000000000",
8212=>"111111101",
8213=>"000000010",
8214=>"101001001",
8215=>"000000001",
8216=>"000000111",
8217=>"010000001",
8218=>"000010111",
8219=>"010110000",
8220=>"000000000",
8221=>"010000000",
8222=>"000100001",
8223=>"000001000",
8224=>"111000100",
8225=>"110100110",
8226=>"001000000",
8227=>"111010000",
8228=>"000000100",
8229=>"000100110",
8230=>"000000000",
8231=>"000000000",
8232=>"100110111",
8233=>"111111111",
8234=>"001000000",
8235=>"011000000",
8236=>"011011111",
8237=>"111111110",
8238=>"001000010",
8239=>"110100000",
8240=>"101001011",
8241=>"001011111",
8242=>"010101000",
8243=>"000100110",
8244=>"000001100",
8245=>"111110000",
8246=>"000100000",
8247=>"010101000",
8248=>"101101000",
8249=>"000001001",
8250=>"010000100",
8251=>"111000001",
8252=>"101100100",
8253=>"110111111",
8254=>"000010000",
8255=>"100011001",
8256=>"101010010",
8257=>"000011111",
8258=>"101111110",
8259=>"000000100",
8260=>"111101100",
8261=>"011000000",
8262=>"110111000",
8263=>"010010000",
8264=>"111000000",
8265=>"111011000",
8266=>"000000000",
8267=>"001101111",
8268=>"000101111",
8269=>"000000111",
8270=>"100101011",
8271=>"101101111",
8272=>"001000001",
8273=>"000011001",
8274=>"010011000",
8275=>"001101001",
8276=>"000011000",
8277=>"101001001",
8278=>"000101001",
8279=>"101101000",
8280=>"110001111",
8281=>"011101011",
8282=>"001111111",
8283=>"000011111",
8284=>"001000110",
8285=>"100000001",
8286=>"011111111",
8287=>"000001101",
8288=>"000111111",
8289=>"111101110",
8290=>"000111011",
8291=>"110000101",
8292=>"001111110",
8293=>"011001001",
8294=>"111110110",
8295=>"111010110",
8296=>"000010011",
8297=>"011001101",
8298=>"010010000",
8299=>"000000010",
8300=>"111000001",
8301=>"010000010",
8302=>"010000010",
8303=>"000000000",
8304=>"001111111",
8305=>"101111101",
8306=>"001001100",
8307=>"101010000",
8308=>"000111011",
8309=>"001100100",
8310=>"000101011",
8311=>"111111001",
8312=>"111000000",
8313=>"110010010",
8314=>"001000000",
8315=>"011000100",
8316=>"011000000",
8317=>"111111100",
8318=>"111010000",
8319=>"100000111",
8320=>"001000000",
8321=>"000101111",
8322=>"110000000",
8323=>"010100000",
8324=>"110010010",
8325=>"111111111",
8326=>"000001111",
8327=>"011000100",
8328=>"111111101",
8329=>"100101111",
8330=>"010100011",
8331=>"000000001",
8332=>"000101100",
8333=>"100110010",
8334=>"101111001",
8335=>"100001000",
8336=>"110111000",
8337=>"010111000",
8338=>"101111010",
8339=>"000010000",
8340=>"010011111",
8341=>"000000010",
8342=>"111101010",
8343=>"100110110",
8344=>"110011010",
8345=>"000000100",
8346=>"110110000",
8347=>"010010111",
8348=>"001000010",
8349=>"100010000",
8350=>"101011111",
8351=>"111001101",
8352=>"000100100",
8353=>"100011001",
8354=>"100000111",
8355=>"000000000",
8356=>"010000000",
8357=>"000010110",
8358=>"011010111",
8359=>"010110010",
8360=>"101000000",
8361=>"001000010",
8362=>"101010001",
8363=>"111101001",
8364=>"111111100",
8365=>"100000000",
8366=>"111111000",
8367=>"011010010",
8368=>"000000010",
8369=>"011000001",
8370=>"101101101",
8371=>"001001001",
8372=>"011011001",
8373=>"011111000",
8374=>"000110110",
8375=>"110111111",
8376=>"100011001",
8377=>"110110110",
8378=>"101111111",
8379=>"000000010",
8380=>"111111010",
8381=>"111111111",
8382=>"010111100",
8383=>"000000111",
8384=>"101000101",
8385=>"000011010",
8386=>"000111100",
8387=>"010111000",
8388=>"010111001",
8389=>"000001111",
8390=>"111000101",
8391=>"100000010",
8392=>"111000001",
8393=>"000100101",
8394=>"101000101",
8395=>"101000100",
8396=>"100010110",
8397=>"110000000",
8398=>"010111000",
8399=>"010110101",
8400=>"010111000",
8401=>"110110001",
8402=>"010000110",
8403=>"011101011",
8404=>"001110111",
8405=>"000001101",
8406=>"100000110",
8407=>"010111111",
8408=>"101001101",
8409=>"000000001",
8410=>"100000001",
8411=>"000000111",
8412=>"101111101",
8413=>"011010010",
8414=>"010110110",
8415=>"010000000",
8416=>"000100011",
8417=>"100101101",
8418=>"010111101",
8419=>"101111100",
8420=>"000000011",
8421=>"111111001",
8422=>"000011010",
8423=>"011011000",
8424=>"000000010",
8425=>"101000111",
8426=>"000000111",
8427=>"101111111",
8428=>"000001000",
8429=>"101011110",
8430=>"000111000",
8431=>"110101000",
8432=>"110111000",
8433=>"000100101",
8434=>"000000110",
8435=>"110011101",
8436=>"110110000",
8437=>"000000111",
8438=>"000000111",
8439=>"001000000",
8440=>"101000000",
8441=>"000000000",
8442=>"111111011",
8443=>"010101101",
8444=>"101100001",
8445=>"000111111",
8446=>"110111000",
8447=>"001111000",
8448=>"011011110",
8449=>"100000011",
8450=>"100000100",
8451=>"100000010",
8452=>"100011011",
8453=>"101100100",
8454=>"111110110",
8455=>"000001001",
8456=>"110100100",
8457=>"000011111",
8458=>"110111000",
8459=>"000100100",
8460=>"100000000",
8461=>"000111100",
8462=>"000111011",
8463=>"011011100",
8464=>"111000100",
8465=>"000000000",
8466=>"010100000",
8467=>"010000000",
8468=>"111000101",
8469=>"000110011",
8470=>"001110001",
8471=>"000011010",
8472=>"001100100",
8473=>"011100000",
8474=>"000011000",
8475=>"111100100",
8476=>"010111111",
8477=>"100000100",
8478=>"111011000",
8479=>"010010110",
8480=>"000011000",
8481=>"111100000",
8482=>"101101011",
8483=>"010011011",
8484=>"000110100",
8485=>"010011000",
8486=>"001010000",
8487=>"110011000",
8488=>"101000100",
8489=>"101100100",
8490=>"111100100",
8491=>"011111111",
8492=>"010011011",
8493=>"111101010",
8494=>"111100000",
8495=>"010000000",
8496=>"000110011",
8497=>"000110000",
8498=>"000010011",
8499=>"011100111",
8500=>"111100000",
8501=>"101111111",
8502=>"101111110",
8503=>"100100100",
8504=>"111001101",
8505=>"111100000",
8506=>"110100111",
8507=>"110100111",
8508=>"010011000",
8509=>"000111010",
8510=>"100000000",
8511=>"011111111",
8512=>"100110011",
8513=>"111001000",
8514=>"110110000",
8515=>"111011110",
8516=>"111101111",
8517=>"100000101",
8518=>"000000011",
8519=>"110011111",
8520=>"001000100",
8521=>"011011010",
8522=>"111111111",
8523=>"100011111",
8524=>"000100000",
8525=>"100101110",
8526=>"111101000",
8527=>"111101111",
8528=>"110111111",
8529=>"111100000",
8530=>"101000100",
8531=>"011001010",
8532=>"111100100",
8533=>"100110100",
8534=>"001011000",
8535=>"001011011",
8536=>"011010100",
8537=>"100100100",
8538=>"110011011",
8539=>"011011001",
8540=>"000011100",
8541=>"000101001",
8542=>"101100101",
8543=>"000100111",
8544=>"011100000",
8545=>"000000110",
8546=>"011011010",
8547=>"001000000",
8548=>"100111100",
8549=>"110100111",
8550=>"010111011",
8551=>"110011011",
8552=>"000111111",
8553=>"000000100",
8554=>"011011011",
8555=>"111111011",
8556=>"111111110",
8557=>"000000100",
8558=>"000000011",
8559=>"111111000",
8560=>"100111100",
8561=>"110000000",
8562=>"010000000",
8563=>"001011001",
8564=>"111111111",
8565=>"100000110",
8566=>"000111011",
8567=>"011000011",
8568=>"111101111",
8569=>"000000011",
8570=>"101100101",
8571=>"000100100",
8572=>"000110011",
8573=>"001110100",
8574=>"011011011",
8575=>"000011011",
8576=>"000100111",
8577=>"000011011",
8578=>"111111011",
8579=>"011110000",
8580=>"110100100",
8581=>"111100111",
8582=>"010001110",
8583=>"100110010",
8584=>"000111000",
8585=>"000111100",
8586=>"111100011",
8587=>"011011011",
8588=>"100000111",
8589=>"111111111",
8590=>"011101001",
8591=>"100001001",
8592=>"100110011",
8593=>"010000110",
8594=>"111000000",
8595=>"100000000",
8596=>"011011001",
8597=>"111000100",
8598=>"111100110",
8599=>"000001000",
8600=>"011011010",
8601=>"000010011",
8602=>"010010010",
8603=>"011000001",
8604=>"110100100",
8605=>"111100100",
8606=>"111000111",
8607=>"000100100",
8608=>"100100100",
8609=>"000100000",
8610=>"110100100",
8611=>"100000111",
8612=>"111011011",
8613=>"000100010",
8614=>"101111111",
8615=>"111100110",
8616=>"100010000",
8617=>"010100100",
8618=>"100100111",
8619=>"100100100",
8620=>"101000101",
8621=>"011100100",
8622=>"110111110",
8623=>"111000000",
8624=>"000100100",
8625=>"000011001",
8626=>"000101100",
8627=>"000010010",
8628=>"011101001",
8629=>"111111111",
8630=>"111100100",
8631=>"011011001",
8632=>"101110100",
8633=>"000011011",
8634=>"010111111",
8635=>"011011001",
8636=>"000100100",
8637=>"011011011",
8638=>"011110111",
8639=>"100000100",
8640=>"110000000",
8641=>"011010000",
8642=>"000111111",
8643=>"011111110",
8644=>"000000001",
8645=>"111001001",
8646=>"110111101",
8647=>"000011010",
8648=>"101100100",
8649=>"011011100",
8650=>"001100111",
8651=>"010111111",
8652=>"110100100",
8653=>"100011111",
8654=>"000000010",
8655=>"100111011",
8656=>"111011000",
8657=>"011101011",
8658=>"110110100",
8659=>"011000011",
8660=>"011011000",
8661=>"000000110",
8662=>"111100000",
8663=>"100001111",
8664=>"011001001",
8665=>"000100000",
8666=>"011011001",
8667=>"101000100",
8668=>"111001001",
8669=>"110101000",
8670=>"111100100",
8671=>"011110100",
8672=>"000000000",
8673=>"101100111",
8674=>"101000000",
8675=>"100110100",
8676=>"000000000",
8677=>"100000000",
8678=>"111100000",
8679=>"010011001",
8680=>"011010000",
8681=>"000000011",
8682=>"011011000",
8683=>"000111011",
8684=>"011110100",
8685=>"000000100",
8686=>"001000000",
8687=>"011001010",
8688=>"110100100",
8689=>"100000100",
8690=>"000010011",
8691=>"010100111",
8692=>"111110000",
8693=>"101010111",
8694=>"000100000",
8695=>"111100110",
8696=>"000000000",
8697=>"111101000",
8698=>"100000000",
8699=>"101111100",
8700=>"010110110",
8701=>"000000000",
8702=>"001110111",
8703=>"111111011",
8704=>"001011101",
8705=>"111100000",
8706=>"101100100",
8707=>"110011010",
8708=>"010011001",
8709=>"011010000",
8710=>"100100100",
8711=>"000010011",
8712=>"000011010",
8713=>"000000010",
8714=>"110100101",
8715=>"000100000",
8716=>"111100111",
8717=>"100100000",
8718=>"101011011",
8719=>"000000100",
8720=>"010011011",
8721=>"110100011",
8722=>"111100100",
8723=>"000000011",
8724=>"101011100",
8725=>"110111000",
8726=>"001110110",
8727=>"111111000",
8728=>"101000000",
8729=>"000111011",
8730=>"001011000",
8731=>"011000001",
8732=>"100100100",
8733=>"111001001",
8734=>"000010000",
8735=>"100100100",
8736=>"110011011",
8737=>"001011100",
8738=>"000011100",
8739=>"011100000",
8740=>"001001011",
8741=>"100101000",
8742=>"000011011",
8743=>"110010100",
8744=>"101011101",
8745=>"010011111",
8746=>"000010010",
8747=>"001011010",
8748=>"000001001",
8749=>"101110001",
8750=>"011011011",
8751=>"011111001",
8752=>"100101111",
8753=>"011011010",
8754=>"000110111",
8755=>"000100111",
8756=>"111100000",
8757=>"001011000",
8758=>"110110001",
8759=>"001100000",
8760=>"000100011",
8761=>"111100101",
8762=>"100100111",
8763=>"000000100",
8764=>"000000100",
8765=>"011111000",
8766=>"000000000",
8767=>"000011010",
8768=>"100000101",
8769=>"001011111",
8770=>"111011110",
8771=>"000011001",
8772=>"111111011",
8773=>"100000100",
8774=>"100100000",
8775=>"000011100",
8776=>"110101111",
8777=>"000100111",
8778=>"101100100",
8779=>"000000100",
8780=>"000011011",
8781=>"000101100",
8782=>"000011101",
8783=>"100100001",
8784=>"101011000",
8785=>"011111111",
8786=>"100000100",
8787=>"011001000",
8788=>"111100000",
8789=>"000100110",
8790=>"100100111",
8791=>"101000000",
8792=>"011000111",
8793=>"000100101",
8794=>"100100100",
8795=>"000011000",
8796=>"000000000",
8797=>"000001001",
8798=>"111111100",
8799=>"100110001",
8800=>"000011011",
8801=>"000010110",
8802=>"111000001",
8803=>"001000100",
8804=>"000000001",
8805=>"111111111",
8806=>"110011111",
8807=>"100011001",
8808=>"000011101",
8809=>"101100111",
8810=>"000111110",
8811=>"101111110",
8812=>"000011011",
8813=>"100100111",
8814=>"000111011",
8815=>"111100111",
8816=>"100101001",
8817=>"010011111",
8818=>"001101110",
8819=>"111111001",
8820=>"011111000",
8821=>"100000010",
8822=>"000000011",
8823=>"000011010",
8824=>"100100111",
8825=>"011010010",
8826=>"001000101",
8827=>"011000101",
8828=>"011000001",
8829=>"000110000",
8830=>"110011110",
8831=>"100011111",
8832=>"000000000",
8833=>"010010010",
8834=>"001011011",
8835=>"101111111",
8836=>"000110000",
8837=>"000011001",
8838=>"001001001",
8839=>"000100101",
8840=>"000111111",
8841=>"011101101",
8842=>"111101111",
8843=>"011011000",
8844=>"000011011",
8845=>"000110111",
8846=>"111000101",
8847=>"101001001",
8848=>"000000100",
8849=>"100110011",
8850=>"110000000",
8851=>"100111100",
8852=>"000010100",
8853=>"000000000",
8854=>"111101101",
8855=>"001011011",
8856=>"011000000",
8857=>"000011011",
8858=>"111100100",
8859=>"010111100",
8860=>"011100101",
8861=>"000000000",
8862=>"001010100",
8863=>"000000000",
8864=>"000100100",
8865=>"110100110",
8866=>"000011001",
8867=>"011111011",
8868=>"011011001",
8869=>"100111010",
8870=>"110011000",
8871=>"000100101",
8872=>"111000111",
8873=>"000011001",
8874=>"110100100",
8875=>"100100100",
8876=>"101111111",
8877=>"000000000",
8878=>"001011101",
8879=>"111111010",
8880=>"000010100",
8881=>"110101101",
8882=>"000001000",
8883=>"011000000",
8884=>"000111010",
8885=>"000100100",
8886=>"000000111",
8887=>"010001101",
8888=>"111000001",
8889=>"100010000",
8890=>"000010100",
8891=>"011111011",
8892=>"101000100",
8893=>"001111111",
8894=>"011111001",
8895=>"000000011",
8896=>"000100000",
8897=>"011000000",
8898=>"000011011",
8899=>"010010010",
8900=>"000100100",
8901=>"000110100",
8902=>"000011011",
8903=>"000100111",
8904=>"011000100",
8905=>"011111011",
8906=>"001101111",
8907=>"011000000",
8908=>"100101101",
8909=>"110101000",
8910=>"100100000",
8911=>"111000100",
8912=>"000000010",
8913=>"000110001",
8914=>"011111001",
8915=>"101100100",
8916=>"000000000",
8917=>"111100110",
8918=>"000010011",
8919=>"000001011",
8920=>"100110100",
8921=>"000000101",
8922=>"011110100",
8923=>"111100100",
8924=>"000010000",
8925=>"000011011",
8926=>"000011001",
8927=>"000000100",
8928=>"111100011",
8929=>"111100100",
8930=>"111100000",
8931=>"000010010",
8932=>"101100110",
8933=>"010011011",
8934=>"000010111",
8935=>"011001110",
8936=>"110110111",
8937=>"100000000",
8938=>"001000100",
8939=>"010100100",
8940=>"001011011",
8941=>"100100111",
8942=>"000000000",
8943=>"010011110",
8944=>"000000100",
8945=>"000001001",
8946=>"011011000",
8947=>"010111000",
8948=>"001011001",
8949=>"101000100",
8950=>"000100000",
8951=>"011001000",
8952=>"011100111",
8953=>"000100110",
8954=>"100100010",
8955=>"000000010",
8956=>"111100100",
8957=>"000000000",
8958=>"100111001",
8959=>"101100101",
8960=>"011010000",
8961=>"000111010",
8962=>"111000110",
8963=>"110111111",
8964=>"101111111",
8965=>"111001000",
8966=>"110101000",
8967=>"000110101",
8968=>"000100110",
8969=>"000000100",
8970=>"110100100",
8971=>"100000000",
8972=>"000111111",
8973=>"010100010",
8974=>"011011110",
8975=>"111111000",
8976=>"111111111",
8977=>"100100100",
8978=>"000101101",
8979=>"111101000",
8980=>"101111110",
8981=>"000111000",
8982=>"011000111",
8983=>"100000100",
8984=>"000101001",
8985=>"111010111",
8986=>"000101110",
8987=>"000000111",
8988=>"100101111",
8989=>"000111110",
8990=>"011000100",
8991=>"100101101",
8992=>"111101000",
8993=>"111111110",
8994=>"010010000",
8995=>"010100000",
8996=>"001001011",
8997=>"111010000",
8998=>"111000101",
8999=>"001000000",
9000=>"100101111",
9001=>"001011000",
9002=>"111101100",
9003=>"111000000",
9004=>"011111111",
9005=>"111010000",
9006=>"101111100",
9007=>"100001001",
9008=>"010100110",
9009=>"111010011",
9010=>"000010000",
9011=>"000011010",
9012=>"010101001",
9013=>"001110100",
9014=>"001000000",
9015=>"111000111",
9016=>"111000000",
9017=>"101001100",
9018=>"010010000",
9019=>"001000000",
9020=>"101000100",
9021=>"111111100",
9022=>"010000101",
9023=>"110111000",
9024=>"000110111",
9025=>"111000000",
9026=>"111111111",
9027=>"101100000",
9028=>"110101010",
9029=>"000110100",
9030=>"001000101",
9031=>"011101000",
9032=>"000101111",
9033=>"000001010",
9034=>"000000101",
9035=>"000000000",
9036=>"111001111",
9037=>"000010110",
9038=>"011011011",
9039=>"111111110",
9040=>"110000101",
9041=>"111000000",
9042=>"111101000",
9043=>"011000000",
9044=>"111001011",
9045=>"011010110",
9046=>"010011011",
9047=>"000000111",
9048=>"010111011",
9049=>"111000011",
9050=>"111101100",
9051=>"100000101",
9052=>"001101001",
9053=>"001001010",
9054=>"000111110",
9055=>"100000000",
9056=>"111101000",
9057=>"101111001",
9058=>"101000111",
9059=>"011001001",
9060=>"111110100",
9061=>"001000000",
9062=>"110111111",
9063=>"001001001",
9064=>"011010000",
9065=>"100101001",
9066=>"000010111",
9067=>"000101000",
9068=>"111111100",
9069=>"000010000",
9070=>"000000000",
9071=>"000010000",
9072=>"000001110",
9073=>"111000101",
9074=>"000000000",
9075=>"000000110",
9076=>"110000000",
9077=>"001000100",
9078=>"000111110",
9079=>"111111000",
9080=>"010110111",
9081=>"101101101",
9082=>"000010110",
9083=>"000001000",
9084=>"100110011",
9085=>"010000100",
9086=>"000000111",
9087=>"000001001",
9088=>"000010000",
9089=>"111100101",
9090=>"100101000",
9091=>"001010010",
9092=>"100100000",
9093=>"000000100",
9094=>"011001100",
9095=>"001011011",
9096=>"011011011",
9097=>"000000000",
9098=>"111111001",
9099=>"100011000",
9100=>"111110010",
9101=>"010100010",
9102=>"110001100",
9103=>"000000010",
9104=>"111000101",
9105=>"110111000",
9106=>"101000111",
9107=>"000000111",
9108=>"000010111",
9109=>"000000101",
9110=>"111101010",
9111=>"000010100",
9112=>"110100000",
9113=>"111110100",
9114=>"111000111",
9115=>"001100110",
9116=>"111101111",
9117=>"000000100",
9118=>"010110110",
9119=>"111000110",
9120=>"000010011",
9121=>"001100000",
9122=>"111011010",
9123=>"011000000",
9124=>"101010000",
9125=>"010110100",
9126=>"000111010",
9127=>"010001111",
9128=>"111000000",
9129=>"001001111",
9130=>"000100000",
9131=>"011000101",
9132=>"000010101",
9133=>"100001101",
9134=>"110000101",
9135=>"111010010",
9136=>"010010010",
9137=>"110101100",
9138=>"110010111",
9139=>"000001000",
9140=>"000011011",
9141=>"111111100",
9142=>"111100000",
9143=>"010011000",
9144=>"000000001",
9145=>"000110110",
9146=>"101000000",
9147=>"010010111",
9148=>"000010000",
9149=>"110111110",
9150=>"001001010",
9151=>"011100101",
9152=>"000000010",
9153=>"111111111",
9154=>"000000100",
9155=>"000001100",
9156=>"000000000",
9157=>"011111101",
9158=>"000000000",
9159=>"001101111",
9160=>"000000000",
9161=>"111101000",
9162=>"111101000",
9163=>"000011010",
9164=>"111000100",
9165=>"011000011",
9166=>"010000111",
9167=>"111000000",
9168=>"100100000",
9169=>"110000111",
9170=>"100111111",
9171=>"111111111",
9172=>"101101111",
9173=>"101000110",
9174=>"111000000",
9175=>"001001111",
9176=>"001000110",
9177=>"000111010",
9178=>"101000010",
9179=>"111000000",
9180=>"010100111",
9181=>"010101100",
9182=>"111111000",
9183=>"000011101",
9184=>"010010011",
9185=>"000100111",
9186=>"101001000",
9187=>"000110110",
9188=>"100100111",
9189=>"101000000",
9190=>"101101111",
9191=>"001001011",
9192=>"111010000",
9193=>"101111111",
9194=>"110010001",
9195=>"001110010",
9196=>"010111110",
9197=>"000000000",
9198=>"000100000",
9199=>"101110000",
9200=>"000100000",
9201=>"111111111",
9202=>"010000011",
9203=>"000100000",
9204=>"011111100",
9205=>"101001101",
9206=>"000000010",
9207=>"001000011",
9208=>"000010010",
9209=>"000000000",
9210=>"001010110",
9211=>"000101111",
9212=>"001000100",
9213=>"001011011",
9214=>"010010011",
9215=>"011100111",
9216=>"000000001",
9217=>"100111111",
9218=>"100000100",
9219=>"000000101",
9220=>"111100000",
9221=>"000000000",
9222=>"111000101",
9223=>"010111110",
9224=>"101100100",
9225=>"010110110",
9226=>"010111010",
9227=>"100000101",
9228=>"000000000",
9229=>"010000011",
9230=>"001001001",
9231=>"111010000",
9232=>"111000010",
9233=>"110010000",
9234=>"010000000",
9235=>"111001000",
9236=>"000000000",
9237=>"000000000",
9238=>"000000011",
9239=>"010011111",
9240=>"001100000",
9241=>"110111101",
9242=>"000111100",
9243=>"011111000",
9244=>"000000011",
9245=>"011110000",
9246=>"111000010",
9247=>"111111010",
9248=>"111111101",
9249=>"100111010",
9250=>"000011011",
9251=>"000011010",
9252=>"110010011",
9253=>"000000000",
9254=>"100000101",
9255=>"000001000",
9256=>"011010111",
9257=>"000000101",
9258=>"001000000",
9259=>"011101000",
9260=>"011011010",
9261=>"000101111",
9262=>"000101111",
9263=>"110100101",
9264=>"000101111",
9265=>"001111111",
9266=>"111011010",
9267=>"111000000",
9268=>"111110110",
9269=>"000000111",
9270=>"000111110",
9271=>"000000111",
9272=>"000110000",
9273=>"101001101",
9274=>"100000100",
9275=>"000101011",
9276=>"000110101",
9277=>"100111010",
9278=>"100000101",
9279=>"101110010",
9280=>"111000000",
9281=>"010000000",
9282=>"000000111",
9283=>"111111100",
9284=>"101101111",
9285=>"000000000",
9286=>"000101111",
9287=>"111110101",
9288=>"001100000",
9289=>"101011111",
9290=>"111101000",
9291=>"100000000",
9292=>"110000010",
9293=>"111100010",
9294=>"111001111",
9295=>"111101111",
9296=>"010110111",
9297=>"010111010",
9298=>"111010101",
9299=>"001000100",
9300=>"010000000",
9301=>"000000100",
9302=>"011011000",
9303=>"111101000",
9304=>"110000010",
9305=>"100100111",
9306=>"001000000",
9307=>"100100000",
9308=>"000111111",
9309=>"001001011",
9310=>"001111000",
9311=>"110111101",
9312=>"111111000",
9313=>"010111011",
9314=>"111111000",
9315=>"100100000",
9316=>"101001100",
9317=>"100001110",
9318=>"111111000",
9319=>"001011111",
9320=>"101001101",
9321=>"111111000",
9322=>"000111111",
9323=>"101000001",
9324=>"000000111",
9325=>"010010000",
9326=>"000000111",
9327=>"101000111",
9328=>"100100100",
9329=>"000101000",
9330=>"010111011",
9331=>"111011101",
9332=>"101011111",
9333=>"000000000",
9334=>"000001001",
9335=>"010000000",
9336=>"001011000",
9337=>"010010000",
9338=>"000011001",
9339=>"000000101",
9340=>"100110010",
9341=>"100000000",
9342=>"000000000",
9343=>"101001100",
9344=>"111000101",
9345=>"011000010",
9346=>"110100110",
9347=>"000000101",
9348=>"111111111",
9349=>"000000100",
9350=>"010000010",
9351=>"000110000",
9352=>"001001001",
9353=>"010010111",
9354=>"101000100",
9355=>"111101100",
9356=>"000000100",
9357=>"010000000",
9358=>"000000100",
9359=>"100000000",
9360=>"011110001",
9361=>"000100000",
9362=>"010111000",
9363=>"111000000",
9364=>"000011111",
9365=>"110011000",
9366=>"111000000",
9367=>"001001111",
9368=>"111111010",
9369=>"000111011",
9370=>"111111111",
9371=>"011001110",
9372=>"101000000",
9373=>"111111000",
9374=>"000000101",
9375=>"010010111",
9376=>"000101101",
9377=>"111000100",
9378=>"110000000",
9379=>"010000111",
9380=>"000000011",
9381=>"111101000",
9382=>"010110000",
9383=>"000010010",
9384=>"110111111",
9385=>"000111111",
9386=>"111000000",
9387=>"111010000",
9388=>"011010000",
9389=>"101101111",
9390=>"010000100",
9391=>"000000111",
9392=>"000000010",
9393=>"111011001",
9394=>"100000000",
9395=>"000000110",
9396=>"110110010",
9397=>"011101000",
9398=>"011011001",
9399=>"000000101",
9400=>"100011000",
9401=>"100111111",
9402=>"000000000",
9403=>"000111100",
9404=>"000110111",
9405=>"010010010",
9406=>"001001000",
9407=>"011110000",
9408=>"000000101",
9409=>"000100111",
9410=>"000111111",
9411=>"100000100",
9412=>"011000001",
9413=>"110110111",
9414=>"000100100",
9415=>"000000111",
9416=>"111000001",
9417=>"000110000",
9418=>"100111111",
9419=>"111101011",
9420=>"101100101",
9421=>"001111110",
9422=>"111111011",
9423=>"111111100",
9424=>"000000000",
9425=>"010110111",
9426=>"011000101",
9427=>"111111010",
9428=>"000000111",
9429=>"110110010",
9430=>"100000110",
9431=>"000111111",
9432=>"000000101",
9433=>"110100111",
9434=>"000100100",
9435=>"000010010",
9436=>"000001000",
9437=>"011010000",
9438=>"111111001",
9439=>"111111000",
9440=>"000000101",
9441=>"000000001",
9442=>"001000000",
9443=>"010000111",
9444=>"111000000",
9445=>"100000000",
9446=>"010000111",
9447=>"011000101",
9448=>"000111111",
9449=>"000111111",
9450=>"000001000",
9451=>"000000001",
9452=>"000100000",
9453=>"111101111",
9454=>"000000000",
9455=>"001010110",
9456=>"111011010",
9457=>"011001001",
9458=>"000000111",
9459=>"001001001",
9460=>"110010011",
9461=>"110000111",
9462=>"000000111",
9463=>"000001001",
9464=>"010111010",
9465=>"001000101",
9466=>"000000000",
9467=>"101011111",
9468=>"111111110",
9469=>"000000011",
9470=>"011011010",
9471=>"000000101",
9472=>"010001000",
9473=>"111011111",
9474=>"100000101",
9475=>"110000001",
9476=>"000100100",
9477=>"000011000",
9478=>"010000010",
9479=>"001010010",
9480=>"110011000",
9481=>"000100100",
9482=>"001001001",
9483=>"000010000",
9484=>"000000000",
9485=>"011111010",
9486=>"000110001",
9487=>"101000111",
9488=>"000000000",
9489=>"000000111",
9490=>"000000000",
9491=>"111111110",
9492=>"001000001",
9493=>"100000101",
9494=>"111000100",
9495=>"010010111",
9496=>"000000000",
9497=>"100001110",
9498=>"101100100",
9499=>"000000111",
9500=>"000000111",
9501=>"000100000",
9502=>"110010000",
9503=>"010010010",
9504=>"101101110",
9505=>"111110100",
9506=>"100111011",
9507=>"101000011",
9508=>"100100100",
9509=>"010010111",
9510=>"000011010",
9511=>"100100111",
9512=>"100100100",
9513=>"001010000",
9514=>"000001000",
9515=>"100000111",
9516=>"000001011",
9517=>"010011101",
9518=>"100000000",
9519=>"000101000",
9520=>"010001000",
9521=>"110100000",
9522=>"001000111",
9523=>"000000111",
9524=>"000000100",
9525=>"010101110",
9526=>"011111000",
9527=>"000000001",
9528=>"111000100",
9529=>"000110000",
9530=>"000110010",
9531=>"101101111",
9532=>"000011111",
9533=>"101111000",
9534=>"111000001",
9535=>"111111101",
9536=>"101100111",
9537=>"111101111",
9538=>"111111000",
9539=>"011011011",
9540=>"111111111",
9541=>"000000100",
9542=>"000000000",
9543=>"000100000",
9544=>"010011001",
9545=>"000000001",
9546=>"010000001",
9547=>"111000000",
9548=>"001000000",
9549=>"001001001",
9550=>"111111110",
9551=>"111001111",
9552=>"111111111",
9553=>"000110111",
9554=>"000000000",
9555=>"110000000",
9556=>"111110101",
9557=>"000001000",
9558=>"100100111",
9559=>"000000000",
9560=>"100000010",
9561=>"001011000",
9562=>"000011000",
9563=>"010111110",
9564=>"000000100",
9565=>"001001010",
9566=>"111111110",
9567=>"110100100",
9568=>"100000000",
9569=>"111101111",
9570=>"100000000",
9571=>"000001111",
9572=>"111111100",
9573=>"011011000",
9574=>"101101111",
9575=>"001111010",
9576=>"010010000",
9577=>"101000111",
9578=>"000010111",
9579=>"101000100",
9580=>"001000000",
9581=>"000101011",
9582=>"101000111",
9583=>"011011011",
9584=>"001011001",
9585=>"000010111",
9586=>"001110100",
9587=>"111111011",
9588=>"100101111",
9589=>"100000111",
9590=>"101011111",
9591=>"111111111",
9592=>"000001111",
9593=>"010000011",
9594=>"111000101",
9595=>"000000100",
9596=>"110011101",
9597=>"110100100",
9598=>"001001010",
9599=>"001000000",
9600=>"111011010",
9601=>"100100000",
9602=>"111111011",
9603=>"111111111",
9604=>"111100100",
9605=>"100001111",
9606=>"100010110",
9607=>"001001101",
9608=>"001110000",
9609=>"111011001",
9610=>"000100100",
9611=>"111000000",
9612=>"010111000",
9613=>"000000000",
9614=>"000000000",
9615=>"000000101",
9616=>"100110110",
9617=>"100101101",
9618=>"110001111",
9619=>"111111000",
9620=>"000110100",
9621=>"100111101",
9622=>"111011000",
9623=>"000011010",
9624=>"111110000",
9625=>"111111111",
9626=>"111111010",
9627=>"101000000",
9628=>"000011011",
9629=>"101101111",
9630=>"100111111",
9631=>"000000000",
9632=>"001101010",
9633=>"000100111",
9634=>"011000010",
9635=>"110010011",
9636=>"100100111",
9637=>"101111111",
9638=>"001001101",
9639=>"011111110",
9640=>"000001011",
9641=>"100100111",
9642=>"101000000",
9643=>"000000000",
9644=>"011011001",
9645=>"111110000",
9646=>"001101001",
9647=>"011010101",
9648=>"000000000",
9649=>"110110100",
9650=>"111011000",
9651=>"101111001",
9652=>"100100111",
9653=>"011110000",
9654=>"101100010",
9655=>"101000011",
9656=>"001110011",
9657=>"000110100",
9658=>"010111011",
9659=>"111010100",
9660=>"111110110",
9661=>"000000000",
9662=>"011111100",
9663=>"000110010",
9664=>"000101111",
9665=>"101101001",
9666=>"110110111",
9667=>"001001111",
9668=>"100001011",
9669=>"100111001",
9670=>"101101100",
9671=>"000011000",
9672=>"000011010",
9673=>"000010010",
9674=>"110000100",
9675=>"101101111",
9676=>"111111111",
9677=>"001011000",
9678=>"000000011",
9679=>"111000000",
9680=>"111111011",
9681=>"010110111",
9682=>"000000101",
9683=>"101100000",
9684=>"000000110",
9685=>"011011011",
9686=>"111010000",
9687=>"111110000",
9688=>"111111010",
9689=>"010000000",
9690=>"110101101",
9691=>"101000100",
9692=>"001001000",
9693=>"100000000",
9694=>"110111111",
9695=>"111011000",
9696=>"111011000",
9697=>"000000101",
9698=>"100000010",
9699=>"011111101",
9700=>"000100111",
9701=>"011100011",
9702=>"000000011",
9703=>"100101011",
9704=>"100000000",
9705=>"101111111",
9706=>"100100101",
9707=>"100101111",
9708=>"110110000",
9709=>"000000000",
9710=>"000000000",
9711=>"000000010",
9712=>"000000110",
9713=>"101010000",
9714=>"100000010",
9715=>"000011100",
9716=>"010100000",
9717=>"111111101",
9718=>"000000000",
9719=>"011100111",
9720=>"101100100",
9721=>"000000100",
9722=>"100100010",
9723=>"000000000",
9724=>"111010000",
9725=>"111100101",
9726=>"100100100",
9727=>"111000000",
9728=>"011100000",
9729=>"000000101",
9730=>"000001000",
9731=>"000111111",
9732=>"011111100",
9733=>"000001111",
9734=>"000111101",
9735=>"010010010",
9736=>"000000000",
9737=>"010010000",
9738=>"110111011",
9739=>"000001000",
9740=>"000000100",
9741=>"000000000",
9742=>"100110100",
9743=>"001111111",
9744=>"001101000",
9745=>"111100101",
9746=>"000000000",
9747=>"111000110",
9748=>"111111111",
9749=>"111000001",
9750=>"000000111",
9751=>"111000101",
9752=>"000000000",
9753=>"000101111",
9754=>"001000000",
9755=>"000000101",
9756=>"111111001",
9757=>"000000000",
9758=>"111101000",
9759=>"100000000",
9760=>"111000011",
9761=>"001000000",
9762=>"010100110",
9763=>"000000000",
9764=>"001111110",
9765=>"011011001",
9766=>"010011011",
9767=>"000111101",
9768=>"010000000",
9769=>"110000000",
9770=>"111111101",
9771=>"111110000",
9772=>"110101100",
9773=>"100000001",
9774=>"011001000",
9775=>"000110110",
9776=>"010000000",
9777=>"000011001",
9778=>"000110011",
9779=>"110000111",
9780=>"111110000",
9781=>"110111111",
9782=>"000000001",
9783=>"101010110",
9784=>"111111010",
9785=>"000000111",
9786=>"010111000",
9787=>"000101111",
9788=>"100111110",
9789=>"111111111",
9790=>"100000100",
9791=>"011111101",
9792=>"100000000",
9793=>"000000101",
9794=>"111100110",
9795=>"000011011",
9796=>"111001101",
9797=>"111110000",
9798=>"010111111",
9799=>"111010000",
9800=>"000001111",
9801=>"101001000",
9802=>"101001111",
9803=>"110110111",
9804=>"111000000",
9805=>"000110110",
9806=>"010011010",
9807=>"111111111",
9808=>"111000000",
9809=>"110110111",
9810=>"100111001",
9811=>"001000000",
9812=>"000000010",
9813=>"001000000",
9814=>"000011111",
9815=>"010111000",
9816=>"001010000",
9817=>"000010011",
9818=>"111011011",
9819=>"110010010",
9820=>"011001000",
9821=>"010010110",
9822=>"000001000",
9823=>"100110000",
9824=>"100101100",
9825=>"010011111",
9826=>"111111111",
9827=>"100100111",
9828=>"000000000",
9829=>"000010100",
9830=>"000101100",
9831=>"111111010",
9832=>"000111111",
9833=>"010000001",
9834=>"111111110",
9835=>"111111000",
9836=>"111111110",
9837=>"101111101",
9838=>"101011011",
9839=>"101000111",
9840=>"010111110",
9841=>"010000000",
9842=>"000000000",
9843=>"110010010",
9844=>"111101000",
9845=>"000000100",
9846=>"000111111",
9847=>"110001000",
9848=>"011011010",
9849=>"000111001",
9850=>"000000111",
9851=>"000000100",
9852=>"000100110",
9853=>"101000000",
9854=>"011111000",
9855=>"000001001",
9856=>"001000000",
9857=>"111100100",
9858=>"111111000",
9859=>"000100111",
9860=>"111010011",
9861=>"100111000",
9862=>"110100100",
9863=>"000110010",
9864=>"000111111",
9865=>"000000001",
9866=>"010010000",
9867=>"011011000",
9868=>"000110000",
9869=>"111110111",
9870=>"010010000",
9871=>"100000000",
9872=>"011111011",
9873=>"111111111",
9874=>"001001101",
9875=>"111000011",
9876=>"000000000",
9877=>"000100000",
9878=>"100010010",
9879=>"100100100",
9880=>"111111000",
9881=>"111000011",
9882=>"000111000",
9883=>"011010110",
9884=>"100000000",
9885=>"101000110",
9886=>"110111110",
9887=>"100101101",
9888=>"000100001",
9889=>"111000000",
9890=>"000111000",
9891=>"000010000",
9892=>"110000111",
9893=>"100011000",
9894=>"000111111",
9895=>"010101000",
9896=>"000000001",
9897=>"000000000",
9898=>"100111000",
9899=>"111110000",
9900=>"011110110",
9901=>"111000000",
9902=>"111000001",
9903=>"110111111",
9904=>"000101111",
9905=>"000000000",
9906=>"100010010",
9907=>"000110111",
9908=>"011111111",
9909=>"010010111",
9910=>"111000000",
9911=>"001001000",
9912=>"000111111",
9913=>"001000010",
9914=>"111111101",
9915=>"111101100",
9916=>"111000000",
9917=>"111111111",
9918=>"100100000",
9919=>"010000000",
9920=>"010000000",
9921=>"000000000",
9922=>"110000100",
9923=>"001011000",
9924=>"000000000",
9925=>"111000000",
9926=>"111011110",
9927=>"000010111",
9928=>"100111100",
9929=>"101000100",
9930=>"111111000",
9931=>"111100111",
9932=>"101001000",
9933=>"000011111",
9934=>"111010000",
9935=>"100111111",
9936=>"001011111",
9937=>"011110111",
9938=>"000110111",
9939=>"000111100",
9940=>"100000011",
9941=>"111110000",
9942=>"000000000",
9943=>"110000100",
9944=>"111001000",
9945=>"010111111",
9946=>"100100110",
9947=>"011000000",
9948=>"000000111",
9949=>"111111111",
9950=>"100111101",
9951=>"111110100",
9952=>"000000000",
9953=>"001000111",
9954=>"000010010",
9955=>"111111111",
9956=>"100000000",
9957=>"011001010",
9958=>"101100000",
9959=>"111000100",
9960=>"100111111",
9961=>"111111111",
9962=>"011111110",
9963=>"001000000",
9964=>"111100100",
9965=>"111001001",
9966=>"001011001",
9967=>"000000000",
9968=>"011111000",
9969=>"111001100",
9970=>"111001001",
9971=>"100100100",
9972=>"110111011",
9973=>"000100111",
9974=>"100101000",
9975=>"010111111",
9976=>"000000111",
9977=>"111000000",
9978=>"001101101",
9979=>"000101101",
9980=>"111110111",
9981=>"011000000",
9982=>"000111100",
9983=>"101101111",
9984=>"001011011",
9985=>"111111000",
9986=>"111001000",
9987=>"110111101",
9988=>"000100100",
9989=>"101001000",
9990=>"000000000",
9991=>"000000101",
9992=>"000110110",
9993=>"000100101",
9994=>"110000100",
9995=>"101001001",
9996=>"111111101",
9997=>"000010111",
9998=>"000100100",
9999=>"101111110",
10000=>"010001000",
10001=>"111000000",
10002=>"110101001",
10003=>"101000010",
10004=>"000100111",
10005=>"001000000",
10006=>"011111001",
10007=>"111111101",
10008=>"101101111",
10009=>"000001011",
10010=>"000000000",
10011=>"000101100",
10012=>"111001011",
10013=>"001001101",
10014=>"110110000",
10015=>"000010110",
10016=>"111000101",
10017=>"001101000",
10018=>"101000010",
10019=>"001110111",
10020=>"111111110",
10021=>"110110100",
10022=>"101000001",
10023=>"100011111",
10024=>"101101111",
10025=>"111001001",
10026=>"001000001",
10027=>"010010111",
10028=>"100100100",
10029=>"000101101",
10030=>"000000000",
10031=>"101100110",
10032=>"011001100",
10033=>"100100100",
10034=>"011010000",
10035=>"101000000",
10036=>"110101001",
10037=>"000111010",
10038=>"000100100",
10039=>"011011000",
10040=>"111111000",
10041=>"010010000",
10042=>"000100000",
10043=>"010000000",
10044=>"000110010",
10045=>"111111111",
10046=>"000000000",
10047=>"000111111",
10048=>"110111101",
10049=>"111111000",
10050=>"011111110",
10051=>"010111011",
10052=>"010000110",
10053=>"010000110",
10054=>"000111001",
10055=>"111000000",
10056=>"100000100",
10057=>"111111111",
10058=>"000000000",
10059=>"000001000",
10060=>"101101101",
10061=>"011111111",
10062=>"010011011",
10063=>"000000000",
10064=>"000000000",
10065=>"111111111",
10066=>"111101010",
10067=>"011011011",
10068=>"100100110",
10069=>"001011010",
10070=>"000011101",
10071=>"111000000",
10072=>"000000101",
10073=>"000110110",
10074=>"010001100",
10075=>"000111100",
10076=>"000010000",
10077=>"000000000",
10078=>"000010111",
10079=>"111100100",
10080=>"000110111",
10081=>"111000001",
10082=>"100101110",
10083=>"000001001",
10084=>"000010011",
10085=>"000010111",
10086=>"000001111",
10087=>"000010010",
10088=>"001101000",
10089=>"111111001",
10090=>"110111111",
10091=>"010110000",
10092=>"111000101",
10093=>"101001101",
10094=>"000010000",
10095=>"010100000",
10096=>"000010111",
10097=>"111111100",
10098=>"010001001",
10099=>"111001000",
10100=>"000011111",
10101=>"010101111",
10102=>"000111110",
10103=>"000000111",
10104=>"101000000",
10105=>"010111111",
10106=>"111111111",
10107=>"111000000",
10108=>"001011010",
10109=>"000110000",
10110=>"100000111",
10111=>"101101111",
10112=>"111010111",
10113=>"111111110",
10114=>"000000111",
10115=>"000000000",
10116=>"000000110",
10117=>"110110100",
10118=>"111111111",
10119=>"000000000",
10120=>"000111111",
10121=>"000000000",
10122=>"000100101",
10123=>"110111000",
10124=>"111000111",
10125=>"000000000",
10126=>"000010111",
10127=>"111001001",
10128=>"000110100",
10129=>"000111110",
10130=>"000101101",
10131=>"011000111",
10132=>"000000000",
10133=>"111011000",
10134=>"111111111",
10135=>"000000011",
10136=>"011011000",
10137=>"010000000",
10138=>"111101000",
10139=>"011000111",
10140=>"000010000",
10141=>"101111111",
10142=>"111011000",
10143=>"111111001",
10144=>"000011011",
10145=>"010000001",
10146=>"011111101",
10147=>"111000000",
10148=>"000001000",
10149=>"000110110",
10150=>"110110100",
10151=>"000010110",
10152=>"111101010",
10153=>"001010111",
10154=>"111111111",
10155=>"111111001",
10156=>"101111110",
10157=>"000111011",
10158=>"100100100",
10159=>"111000000",
10160=>"001011001",
10161=>"001000100",
10162=>"000010010",
10163=>"000011000",
10164=>"101011101",
10165=>"011010000",
10166=>"010111110",
10167=>"010110010",
10168=>"011011010",
10169=>"000000000",
10170=>"010110100",
10171=>"000110100",
10172=>"110000011",
10173=>"101101111",
10174=>"000111111",
10175=>"111000000",
10176=>"010110110",
10177=>"010010000",
10178=>"010100100",
10179=>"111011011",
10180=>"000001101",
10181=>"111101010",
10182=>"111111010",
10183=>"010000010",
10184=>"001000101",
10185=>"001010110",
10186=>"000000110",
10187=>"000111111",
10188=>"000000111",
10189=>"000100111",
10190=>"010111111",
10191=>"111000010",
10192=>"110001001",
10193=>"010011000",
10194=>"000000111",
10195=>"010111101",
10196=>"001001000",
10197=>"000000000",
10198=>"110110100",
10199=>"111110000",
10200=>"001001010",
10201=>"101000011",
10202=>"000111000",
10203=>"111000000",
10204=>"100111110",
10205=>"101000000",
10206=>"000111101",
10207=>"111110111",
10208=>"101001110",
10209=>"000000000",
10210=>"101011111",
10211=>"000000001",
10212=>"111001101",
10213=>"000000110",
10214=>"111001000",
10215=>"010011001",
10216=>"111111111",
10217=>"000000100",
10218=>"001000000",
10219=>"111010100",
10220=>"001000000",
10221=>"000001111",
10222=>"000100001",
10223=>"000110010",
10224=>"111000111",
10225=>"011111111",
10226=>"011111000",
10227=>"000011111",
10228=>"000110110",
10229=>"111000101",
10230=>"111000000",
10231=>"001100111",
10232=>"000010010",
10233=>"101010110",
10234=>"111101000",
10235=>"000000001",
10236=>"000000010",
10237=>"000000000",
10238=>"000011001",
10239=>"111000000",
10240=>"001001011",
10241=>"100101100",
10242=>"101000001",
10243=>"101111100",
10244=>"011011111",
10245=>"000000000",
10246=>"000000001",
10247=>"101110110",
10248=>"110111000",
10249=>"000101101",
10250=>"001000100",
10251=>"111000000",
10252=>"111001101",
10253=>"110100111",
10254=>"110111001",
10255=>"000000110",
10256=>"110010010",
10257=>"100101101",
10258=>"000000101",
10259=>"111010000",
10260=>"101010100",
10261=>"110000000",
10262=>"011100100",
10263=>"111001000",
10264=>"111110000",
10265=>"111110111",
10266=>"000000001",
10267=>"001101111",
10268=>"000111001",
10269=>"001111011",
10270=>"000000000",
10271=>"000000101",
10272=>"111110000",
10273=>"010010110",
10274=>"000000000",
10275=>"010111000",
10276=>"100101100",
10277=>"100100100",
10278=>"111010000",
10279=>"001000000",
10280=>"010011000",
10281=>"100111111",
10282=>"010000000",
10283=>"000000000",
10284=>"111001011",
10285=>"111010101",
10286=>"100101110",
10287=>"000000000",
10288=>"000010000",
10289=>"011000000",
10290=>"000010011",
10291=>"001000010",
10292=>"000000101",
10293=>"111000010",
10294=>"000000000",
10295=>"011111010",
10296=>"111010000",
10297=>"111100100",
10298=>"110110010",
10299=>"100000000",
10300=>"000010110",
10301=>"011011010",
10302=>"100101111",
10303=>"110011010",
10304=>"000011111",
10305=>"111000000",
10306=>"111111100",
10307=>"110110000",
10308=>"101001000",
10309=>"101010010",
10310=>"000101101",
10311=>"111111111",
10312=>"110010001",
10313=>"000010011",
10314=>"101010000",
10315=>"010111100",
10316=>"000101000",
10317=>"001101010",
10318=>"100000101",
10319=>"000000011",
10320=>"000000101",
10321=>"111000111",
10322=>"110111000",
10323=>"011101000",
10324=>"001101111",
10325=>"000100001",
10326=>"011011000",
10327=>"100000111",
10328=>"000001111",
10329=>"001011000",
10330=>"000101101",
10331=>"100011000",
10332=>"101000000",
10333=>"000001111",
10334=>"111101111",
10335=>"110011011",
10336=>"100000000",
10337=>"001000010",
10338=>"000000000",
10339=>"110000101",
10340=>"111110010",
10341=>"000100110",
10342=>"000100110",
10343=>"111111110",
10344=>"101000110",
10345=>"111000000",
10346=>"000111111",
10347=>"110000001",
10348=>"000111010",
10349=>"010110111",
10350=>"000000011",
10351=>"111111000",
10352=>"001101000",
10353=>"100010000",
10354=>"000000000",
10355=>"000000001",
10356=>"111111101",
10357=>"101100100",
10358=>"000110111",
10359=>"010111000",
10360=>"011011010",
10361=>"000100111",
10362=>"011000101",
10363=>"111111010",
10364=>"100110111",
10365=>"100101100",
10366=>"111001010",
10367=>"111000000",
10368=>"111100000",
10369=>"110111111",
10370=>"010111000",
10371=>"000111111",
10372=>"000000111",
10373=>"000001100",
10374=>"001001000",
10375=>"100011001",
10376=>"100100000",
10377=>"000000101",
10378=>"100000000",
10379=>"101111000",
10380=>"010010000",
10381=>"101001111",
10382=>"101111000",
10383=>"001000101",
10384=>"100011001",
10385=>"011001000",
10386=>"111000100",
10387=>"000010111",
10388=>"000101001",
10389=>"010010010",
10390=>"111011000",
10391=>"001001000",
10392=>"100111100",
10393=>"100110111",
10394=>"000000101",
10395=>"000000101",
10396=>"111111101",
10397=>"000101010",
10398=>"111000111",
10399=>"000100010",
10400=>"101011111",
10401=>"000000011",
10402=>"111111111",
10403=>"111110111",
10404=>"010101110",
10405=>"100110000",
10406=>"100110001",
10407=>"001111111",
10408=>"111100000",
10409=>"000010111",
10410=>"111010110",
10411=>"111111000",
10412=>"010111000",
10413=>"110000000",
10414=>"000001101",
10415=>"111101111",
10416=>"010010001",
10417=>"000100010",
10418=>"111111110",
10419=>"001110110",
10420=>"000001000",
10421=>"000001000",
10422=>"111011011",
10423=>"001000100",
10424=>"000010011",
10425=>"000111110",
10426=>"111101111",
10427=>"000000000",
10428=>"010000000",
10429=>"011010010",
10430=>"011011000",
10431=>"101000000",
10432=>"101000000",
10433=>"100000101",
10434=>"010000000",
10435=>"111001001",
10436=>"011000100",
10437=>"001001000",
10438=>"111111000",
10439=>"111111101",
10440=>"011111100",
10441=>"000101111",
10442=>"111111100",
10443=>"000000000",
10444=>"000111111",
10445=>"000011111",
10446=>"000010010",
10447=>"111111000",
10448=>"000000011",
10449=>"000110011",
10450=>"101011111",
10451=>"000011111",
10452=>"000001010",
10453=>"000000000",
10454=>"101000000",
10455=>"000111110",
10456=>"111000000",
10457=>"000000101",
10458=>"000001010",
10459=>"000000000",
10460=>"001111100",
10461=>"111111100",
10462=>"100000100",
10463=>"101111111",
10464=>"001000000",
10465=>"000000111",
10466=>"000101111",
10467=>"101001100",
10468=>"111000011",
10469=>"101000000",
10470=>"011011111",
10471=>"100100111",
10472=>"000001111",
10473=>"001011111",
10474=>"100000000",
10475=>"011010001",
10476=>"000111000",
10477=>"101000000",
10478=>"000000000",
10479=>"110000000",
10480=>"010010000",
10481=>"001011100",
10482=>"010000000",
10483=>"000100100",
10484=>"100101011",
10485=>"111000111",
10486=>"000000100",
10487=>"010001001",
10488=>"000011010",
10489=>"110010111",
10490=>"111111101",
10491=>"000000000",
10492=>"010111000",
10493=>"000000011",
10494=>"100111111",
10495=>"000111101",
10496=>"100100100",
10497=>"011010000",
10498=>"000000000",
10499=>"000000000",
10500=>"100000011",
10501=>"001011101",
10502=>"111111001",
10503=>"101111111",
10504=>"001001001",
10505=>"000000000",
10506=>"111111111",
10507=>"010110001",
10508=>"001001100",
10509=>"000000100",
10510=>"010110111",
10511=>"101111111",
10512=>"111010011",
10513=>"111111110",
10514=>"111010010",
10515=>"111111111",
10516=>"111110111",
10517=>"111111111",
10518=>"001000010",
10519=>"010111110",
10520=>"110000101",
10521=>"111011011",
10522=>"101000111",
10523=>"000000000",
10524=>"011111111",
10525=>"001111111",
10526=>"000000011",
10527=>"000010010",
10528=>"000001001",
10529=>"000000000",
10530=>"000000010",
10531=>"000000000",
10532=>"110111000",
10533=>"011001001",
10534=>"010010011",
10535=>"000000000",
10536=>"000011111",
10537=>"001110000",
10538=>"111111111",
10539=>"110111100",
10540=>"110010000",
10541=>"111000001",
10542=>"001100010",
10543=>"101101000",
10544=>"100000000",
10545=>"001000000",
10546=>"001111000",
10547=>"111111111",
10548=>"111111111",
10549=>"110101011",
10550=>"111111111",
10551=>"001111111",
10552=>"110010101",
10553=>"111010111",
10554=>"011000111",
10555=>"011000000",
10556=>"000001011",
10557=>"111011011",
10558=>"000001001",
10559=>"001000011",
10560=>"111111110",
10561=>"000000011",
10562=>"000000000",
10563=>"000101100",
10564=>"000000000",
10565=>"001011101",
10566=>"101111000",
10567=>"000101111",
10568=>"110000000",
10569=>"000000000",
10570=>"011111101",
10571=>"111111011",
10572=>"111111111",
10573=>"111111001",
10574=>"100100000",
10575=>"000000010",
10576=>"111111111",
10577=>"111011110",
10578=>"111001000",
10579=>"000100100",
10580=>"100001000",
10581=>"001000000",
10582=>"000001011",
10583=>"000000001",
10584=>"011011111",
10585=>"001110110",
10586=>"111111111",
10587=>"100111111",
10588=>"110011001",
10589=>"000000110",
10590=>"001100001",
10591=>"001011101",
10592=>"111111111",
10593=>"000000101",
10594=>"111111111",
10595=>"101100000",
10596=>"000000000",
10597=>"111111111",
10598=>"000001111",
10599=>"000001011",
10600=>"000000000",
10601=>"111101111",
10602=>"111111111",
10603=>"010111111",
10604=>"011000000",
10605=>"111111111",
10606=>"000000000",
10607=>"111110111",
10608=>"110111110",
10609=>"111111111",
10610=>"111111111",
10611=>"000111111",
10612=>"000111111",
10613=>"010111111",
10614=>"000110010",
10615=>"000010110",
10616=>"000001101",
10617=>"110000000",
10618=>"110111111",
10619=>"000000000",
10620=>"011001001",
10621=>"001001001",
10622=>"000011000",
10623=>"000000010",
10624=>"000000101",
10625=>"111111101",
10626=>"000001000",
10627=>"000001000",
10628=>"101101111",
10629=>"000111111",
10630=>"011100010",
10631=>"111010010",
10632=>"111111000",
10633=>"001000111",
10634=>"000100001",
10635=>"000111110",
10636=>"100110000",
10637=>"001101000",
10638=>"101111011",
10639=>"000000101",
10640=>"111111111",
10641=>"111111110",
10642=>"111001000",
10643=>"000101111",
10644=>"000100111",
10645=>"001011111",
10646=>"111111001",
10647=>"000011010",
10648=>"000100100",
10649=>"000111001",
10650=>"000110110",
10651=>"000000001",
10652=>"101000100",
10653=>"110110000",
10654=>"100000101",
10655=>"011000010",
10656=>"000000000",
10657=>"111000000",
10658=>"000000000",
10659=>"111000000",
10660=>"111111111",
10661=>"111011111",
10662=>"000000111",
10663=>"000000000",
10664=>"111000000",
10665=>"000000000",
10666=>"111111111",
10667=>"111111111",
10668=>"001000111",
10669=>"111000111",
10670=>"011011011",
10671=>"001000001",
10672=>"000001101",
10673=>"101111110",
10674=>"001010010",
10675=>"000110110",
10676=>"010110111",
10677=>"011110000",
10678=>"011000000",
10679=>"110111000",
10680=>"000000110",
10681=>"011111100",
10682=>"000001111",
10683=>"110111000",
10684=>"000000001",
10685=>"000110010",
10686=>"000000001",
10687=>"000000000",
10688=>"001001110",
10689=>"110111010",
10690=>"100000101",
10691=>"110110110",
10692=>"110000000",
10693=>"110111001",
10694=>"010000000",
10695=>"000000111",
10696=>"000000101",
10697=>"000001001",
10698=>"110111001",
10699=>"110110000",
10700=>"011111011",
10701=>"111110111",
10702=>"010110111",
10703=>"011110001",
10704=>"010010010",
10705=>"000000011",
10706=>"000010010",
10707=>"111111010",
10708=>"000011011",
10709=>"011011000",
10710=>"000000001",
10711=>"111111111",
10712=>"011001000",
10713=>"000000000",
10714=>"000000000",
10715=>"111110111",
10716=>"000000000",
10717=>"000000000",
10718=>"111111111",
10719=>"010011111",
10720=>"001000000",
10721=>"111111110",
10722=>"001001101",
10723=>"111111100",
10724=>"101001001",
10725=>"111111111",
10726=>"000000111",
10727=>"101010000",
10728=>"000000010",
10729=>"010001001",
10730=>"111111111",
10731=>"111101111",
10732=>"111001001",
10733=>"111111111",
10734=>"111110000",
10735=>"000000001",
10736=>"000100111",
10737=>"111111000",
10738=>"000000000",
10739=>"000000111",
10740=>"000001000",
10741=>"111111111",
10742=>"110111111",
10743=>"000001111",
10744=>"000000110",
10745=>"001000000",
10746=>"000111100",
10747=>"001110110",
10748=>"111111010",
10749=>"000101001",
10750=>"011110110",
10751=>"111111010",
10752=>"011001101",
10753=>"000000011",
10754=>"001000001",
10755=>"010111000",
10756=>"111111101",
10757=>"111111111",
10758=>"111111001",
10759=>"100000000",
10760=>"011111111",
10761=>"010010000",
10762=>"110110100",
10763=>"101111111",
10764=>"000000000",
10765=>"111011111",
10766=>"111011110",
10767=>"000000000",
10768=>"111000110",
10769=>"010000000",
10770=>"000000111",
10771=>"001001000",
10772=>"101111100",
10773=>"111101001",
10774=>"011101101",
10775=>"111111010",
10776=>"000000000",
10777=>"111111111",
10778=>"100100000",
10779=>"010011111",
10780=>"010010111",
10781=>"000000010",
10782=>"111111000",
10783=>"000000000",
10784=>"000010100",
10785=>"001110111",
10786=>"000011111",
10787=>"101111110",
10788=>"000100100",
10789=>"100100100",
10790=>"001111010",
10791=>"110110110",
10792=>"111111010",
10793=>"110111100",
10794=>"000000000",
10795=>"001110010",
10796=>"000011001",
10797=>"111111110",
10798=>"100000000",
10799=>"010000011",
10800=>"000001000",
10801=>"000000001",
10802=>"111111111",
10803=>"010000001",
10804=>"011111110",
10805=>"000010000",
10806=>"011000000",
10807=>"000000000",
10808=>"101000000",
10809=>"000000000",
10810=>"000010011",
10811=>"010000010",
10812=>"001100011",
10813=>"000000101",
10814=>"000000000",
10815=>"100110111",
10816=>"000001101",
10817=>"001000000",
10818=>"010110111",
10819=>"011011100",
10820=>"000010000",
10821=>"000001001",
10822=>"000010000",
10823=>"011000101",
10824=>"100011011",
10825=>"111111111",
10826=>"111001001",
10827=>"001100100",
10828=>"000000000",
10829=>"001001001",
10830=>"001001100",
10831=>"000000101",
10832=>"000000000",
10833=>"100100110",
10834=>"111111100",
10835=>"001000000",
10836=>"000000000",
10837=>"000000111",
10838=>"011101111",
10839=>"110010110",
10840=>"000000101",
10841=>"000000001",
10842=>"000100000",
10843=>"001000111",
10844=>"000010000",
10845=>"000110001",
10846=>"010000000",
10847=>"100101011",
10848=>"111110010",
10849=>"001111111",
10850=>"110010010",
10851=>"010010111",
10852=>"000000001",
10853=>"111111111",
10854=>"111111111",
10855=>"110110111",
10856=>"111111111",
10857=>"111111011",
10858=>"000000100",
10859=>"111111111",
10860=>"001100111",
10861=>"111111111",
10862=>"111000000",
10863=>"000000101",
10864=>"100100100",
10865=>"001001000",
10866=>"110000000",
10867=>"111110110",
10868=>"001000101",
10869=>"000000000",
10870=>"111010101",
10871=>"000000000",
10872=>"000000000",
10873=>"000000000",
10874=>"000111111",
10875=>"111111111",
10876=>"011110111",
10877=>"110100000",
10878=>"111110110",
10879=>"101111001",
10880=>"000010101",
10881=>"111101100",
10882=>"001111011",
10883=>"000000000",
10884=>"101001000",
10885=>"111110110",
10886=>"001011001",
10887=>"000001001",
10888=>"011011010",
10889=>"011000001",
10890=>"101111010",
10891=>"110010000",
10892=>"101000100",
10893=>"110110100",
10894=>"000001000",
10895=>"000000000",
10896=>"110100100",
10897=>"111000000",
10898=>"001000001",
10899=>"001110111",
10900=>"001000011",
10901=>"111000110",
10902=>"010000000",
10903=>"000000000",
10904=>"110000000",
10905=>"111111111",
10906=>"100100100",
10907=>"110000000",
10908=>"111111000",
10909=>"000000011",
10910=>"111000000",
10911=>"001010000",
10912=>"000111101",
10913=>"010010110",
10914=>"000010111",
10915=>"110001000",
10916=>"000000110",
10917=>"000000001",
10918=>"000111001",
10919=>"100100000",
10920=>"111111011",
10921=>"100101000",
10922=>"001010011",
10923=>"111001111",
10924=>"111100111",
10925=>"001001101",
10926=>"100110011",
10927=>"000111100",
10928=>"011110100",
10929=>"000100101",
10930=>"010110010",
10931=>"000000100",
10932=>"101101101",
10933=>"111111110",
10934=>"101000000",
10935=>"110111111",
10936=>"000000110",
10937=>"000000100",
10938=>"010000001",
10939=>"111101011",
10940=>"000000000",
10941=>"111000100",
10942=>"111111110",
10943=>"111001001",
10944=>"111111111",
10945=>"000000000",
10946=>"110000000",
10947=>"001001000",
10948=>"111110010",
10949=>"100010011",
10950=>"101000010",
10951=>"011111111",
10952=>"010111110",
10953=>"000000000",
10954=>"111011100",
10955=>"000100000",
10956=>"000000000",
10957=>"000001110",
10958=>"000000100",
10959=>"000001001",
10960=>"101000000",
10961=>"011111000",
10962=>"000100001",
10963=>"011000000",
10964=>"000000000",
10965=>"001011111",
10966=>"111111000",
10967=>"110000010",
10968=>"000000111",
10969=>"100100000",
10970=>"000111001",
10971=>"000000000",
10972=>"110000100",
10973=>"000101110",
10974=>"101000000",
10975=>"110000000",
10976=>"011001001",
10977=>"000110110",
10978=>"101110111",
10979=>"111111111",
10980=>"111000000",
10981=>"000010000",
10982=>"101011111",
10983=>"010010100",
10984=>"001001110",
10985=>"100010000",
10986=>"011111011",
10987=>"010111110",
10988=>"000000000",
10989=>"111001110",
10990=>"000000000",
10991=>"000000000",
10992=>"101000000",
10993=>"001110100",
10994=>"001000001",
10995=>"000000100",
10996=>"100000001",
10997=>"111111111",
10998=>"010000000",
10999=>"000000001",
11000=>"000001000",
11001=>"111111000",
11002=>"100110110",
11003=>"000010111",
11004=>"010100111",
11005=>"000111000",
11006=>"001001001",
11007=>"011101001",
11008=>"011001001",
11009=>"000000101",
11010=>"101000001",
11011=>"000110011",
11012=>"011011101",
11013=>"000000000",
11014=>"111000000",
11015=>"011001011",
11016=>"000000000",
11017=>"010111000",
11018=>"000000000",
11019=>"000000111",
11020=>"101111111",
11021=>"000100110",
11022=>"011110001",
11023=>"000000000",
11024=>"111000000",
11025=>"110111010",
11026=>"000001000",
11027=>"000001111",
11028=>"111111000",
11029=>"101001000",
11030=>"100100001",
11031=>"000111111",
11032=>"111000101",
11033=>"111001101",
11034=>"010011001",
11035=>"010010110",
11036=>"000000101",
11037=>"000001001",
11038=>"111100001",
11039=>"000111110",
11040=>"000000001",
11041=>"111111011",
11042=>"000110010",
11043=>"111111111",
11044=>"001011011",
11045=>"100111011",
11046=>"110110110",
11047=>"111111000",
11048=>"010010000",
11049=>"110110001",
11050=>"100110000",
11051=>"010000000",
11052=>"001111101",
11053=>"101111111",
11054=>"111000000",
11055=>"000001010",
11056=>"111111111",
11057=>"011011000",
11058=>"001101101",
11059=>"101001001",
11060=>"100000100",
11061=>"000110000",
11062=>"000000011",
11063=>"010000111",
11064=>"111111111",
11065=>"000000100",
11066=>"000001000",
11067=>"010100000",
11068=>"110000001",
11069=>"111111000",
11070=>"000100100",
11071=>"001111100",
11072=>"111001011",
11073=>"110010101",
11074=>"001101101",
11075=>"100011001",
11076=>"000000111",
11077=>"001000000",
11078=>"000101000",
11079=>"001001110",
11080=>"000001111",
11081=>"111111000",
11082=>"000111111",
11083=>"111101110",
11084=>"110111000",
11085=>"100100100",
11086=>"110110100",
11087=>"111011110",
11088=>"000000110",
11089=>"111111010",
11090=>"001000101",
11091=>"001001000",
11092=>"010010000",
11093=>"100100001",
11094=>"100110111",
11095=>"110111001",
11096=>"101101101",
11097=>"100001000",
11098=>"100111110",
11099=>"010000010",
11100=>"010000000",
11101=>"001001000",
11102=>"101011011",
11103=>"010100000",
11104=>"111111111",
11105=>"010011001",
11106=>"011000001",
11107=>"001001101",
11108=>"000101001",
11109=>"001001010",
11110=>"110110000",
11111=>"011111000",
11112=>"011010111",
11113=>"111001000",
11114=>"111100111",
11115=>"001111111",
11116=>"000110111",
11117=>"000011010",
11118=>"000001111",
11119=>"111001111",
11120=>"111111100",
11121=>"000111111",
11122=>"011100100",
11123=>"101101000",
11124=>"010000000",
11125=>"000000001",
11126=>"000111111",
11127=>"110111000",
11128=>"000000111",
11129=>"001111111",
11130=>"000000111",
11131=>"101101100",
11132=>"000110000",
11133=>"100100000",
11134=>"010011001",
11135=>"010000000",
11136=>"111010010",
11137=>"111110000",
11138=>"111001001",
11139=>"100100111",
11140=>"111000000",
11141=>"101111101",
11142=>"011101100",
11143=>"100001001",
11144=>"011001000",
11145=>"001010110",
11146=>"000000000",
11147=>"111001000",
11148=>"000000000",
11149=>"011000000",
11150=>"111001110",
11151=>"000000101",
11152=>"111101111",
11153=>"000110110",
11154=>"010010000",
11155=>"000000110",
11156=>"000000000",
11157=>"000000000",
11158=>"111111111",
11159=>"011011000",
11160=>"010110111",
11161=>"000101111",
11162=>"000001011",
11163=>"010000000",
11164=>"100000000",
11165=>"101000100",
11166=>"111000000",
11167=>"000000010",
11168=>"110100110",
11169=>"000000111",
11170=>"111101100",
11171=>"101111101",
11172=>"010000001",
11173=>"001000101",
11174=>"010110000",
11175=>"000000101",
11176=>"111000001",
11177=>"100111000",
11178=>"000011010",
11179=>"001000000",
11180=>"001001011",
11181=>"110000100",
11182=>"010000110",
11183=>"000000001",
11184=>"000001111",
11185=>"011101101",
11186=>"000000000",
11187=>"111001001",
11188=>"100111011",
11189=>"001111111",
11190=>"000111110",
11191=>"000110000",
11192=>"000100100",
11193=>"001110110",
11194=>"010000010",
11195=>"000010111",
11196=>"011110011",
11197=>"111101000",
11198=>"100000000",
11199=>"000000110",
11200=>"000001111",
11201=>"010010000",
11202=>"111110111",
11203=>"100100000",
11204=>"111111000",
11205=>"010110111",
11206=>"000110111",
11207=>"010010000",
11208=>"101111111",
11209=>"000010000",
11210=>"111101000",
11211=>"000000111",
11212=>"010000000",
11213=>"001011001",
11214=>"001100101",
11215=>"000000000",
11216=>"000000000",
11217=>"001111010",
11218=>"001110011",
11219=>"100000011",
11220=>"110111000",
11221=>"101001101",
11222=>"111110000",
11223=>"000000000",
11224=>"000101111",
11225=>"111000111",
11226=>"011011000",
11227=>"111000000",
11228=>"011001000",
11229=>"011111011",
11230=>"101101101",
11231=>"011001000",
11232=>"010010000",
11233=>"000000001",
11234=>"010111000",
11235=>"110100000",
11236=>"111111000",
11237=>"010010111",
11238=>"101011100",
11239=>"001001001",
11240=>"111111000",
11241=>"101111011",
11242=>"000110001",
11243=>"111111011",
11244=>"111000000",
11245=>"000111111",
11246=>"111000000",
11247=>"100000110",
11248=>"101111011",
11249=>"001001010",
11250=>"010010000",
11251=>"000101111",
11252=>"110100100",
11253=>"101000101",
11254=>"000100000",
11255=>"000000100",
11256=>"000000000",
11257=>"011000100",
11258=>"111100111",
11259=>"000101000",
11260=>"000001111",
11261=>"000000100",
11262=>"100100110",
11263=>"111000110",
11264=>"000111100",
11265=>"101111000",
11266=>"100000100",
11267=>"100110010",
11268=>"000011001",
11269=>"000000111",
11270=>"000000000",
11271=>"000011110",
11272=>"111011000",
11273=>"100000000",
11274=>"000110100",
11275=>"111101101",
11276=>"111000000",
11277=>"111101000",
11278=>"000110001",
11279=>"001000000",
11280=>"000100111",
11281=>"111000111",
11282=>"110110100",
11283=>"000000010",
11284=>"010111111",
11285=>"000010111",
11286=>"011011111",
11287=>"111000101",
11288=>"101000000",
11289=>"110010010",
11290=>"000011001",
11291=>"110111000",
11292=>"100111101",
11293=>"111001000",
11294=>"000011010",
11295=>"001000000",
11296=>"000111000",
11297=>"000111111",
11298=>"100101111",
11299=>"000000111",
11300=>"011001001",
11301=>"011111101",
11302=>"000111111",
11303=>"011110011",
11304=>"100100000",
11305=>"000010010",
11306=>"000000000",
11307=>"101110000",
11308=>"110011011",
11309=>"111111001",
11310=>"000111111",
11311=>"110111001",
11312=>"100000101",
11313=>"011100001",
11314=>"111100000",
11315=>"000111111",
11316=>"000111111",
11317=>"100000111",
11318=>"001000001",
11319=>"111100001",
11320=>"010111111",
11321=>"000000010",
11322=>"111111110",
11323=>"010010000",
11324=>"110110110",
11325=>"111111111",
11326=>"000000101",
11327=>"000000100",
11328=>"001000000",
11329=>"100011000",
11330=>"111111111",
11331=>"000000100",
11332=>"000111111",
11333=>"000000000",
11334=>"001000000",
11335=>"000000111",
11336=>"111111001",
11337=>"101111011",
11338=>"111000000",
11339=>"101111111",
11340=>"000111011",
11341=>"000100110",
11342=>"000011111",
11343=>"000000000",
11344=>"001011001",
11345=>"111111100",
11346=>"000000011",
11347=>"011001011",
11348=>"000100110",
11349=>"110111111",
11350=>"110100100",
11351=>"100000011",
11352=>"000001001",
11353=>"010110110",
11354=>"100110100",
11355=>"000100110",
11356=>"000111010",
11357=>"000001000",
11358=>"110010110",
11359=>"000000001",
11360=>"000000111",
11361=>"000001011",
11362=>"000000000",
11363=>"000001011",
11364=>"001110000",
11365=>"010100000",
11366=>"000111110",
11367=>"111111100",
11368=>"000110010",
11369=>"100100000",
11370=>"111110100",
11371=>"000010100",
11372=>"000010111",
11373=>"000000101",
11374=>"010000101",
11375=>"111011000",
11376=>"100111111",
11377=>"111111101",
11378=>"110100110",
11379=>"100000111",
11380=>"111111100",
11381=>"001000001",
11382=>"001011000",
11383=>"000000000",
11384=>"111100000",
11385=>"001111000",
11386=>"111001111",
11387=>"000110111",
11388=>"001110111",
11389=>"111000000",
11390=>"000100111",
11391=>"000000101",
11392=>"110101110",
11393=>"111001001",
11394=>"000000001",
11395=>"101000010",
11396=>"000010111",
11397=>"111001100",
11398=>"110111011",
11399=>"000011010",
11400=>"100111111",
11401=>"101111100",
11402=>"000010000",
11403=>"000010001",
11404=>"111000101",
11405=>"111000100",
11406=>"000011100",
11407=>"011001011",
11408=>"001011011",
11409=>"011111111",
11410=>"000000000",
11411=>"000111111",
11412=>"010010010",
11413=>"101000000",
11414=>"111100000",
11415=>"000100000",
11416=>"100000100",
11417=>"110100011",
11418=>"111000000",
11419=>"000000000",
11420=>"111111000",
11421=>"010000011",
11422=>"111011011",
11423=>"101111110",
11424=>"011001000",
11425=>"111111101",
11426=>"111101000",
11427=>"010111001",
11428=>"110111111",
11429=>"110100000",
11430=>"011001100",
11431=>"100111111",
11432=>"101010111",
11433=>"001000111",
11434=>"111100100",
11435=>"000000111",
11436=>"111100111",
11437=>"000111111",
11438=>"111111101",
11439=>"101101110",
11440=>"101000100",
11441=>"010101101",
11442=>"000000000",
11443=>"000000000",
11444=>"111000101",
11445=>"111111101",
11446=>"001110000",
11447=>"110111110",
11448=>"011011011",
11449=>"001000110",
11450=>"000011101",
11451=>"110011010",
11452=>"010011001",
11453=>"111000101",
11454=>"100100000",
11455=>"011010101",
11456=>"000010000",
11457=>"110000000",
11458=>"110010000",
11459=>"000110110",
11460=>"000011100",
11461=>"000110111",
11462=>"000000011",
11463=>"101100100",
11464=>"000101001",
11465=>"001111100",
11466=>"000010111",
11467=>"111000111",
11468=>"000010001",
11469=>"001011011",
11470=>"110010100",
11471=>"111011100",
11472=>"111100000",
11473=>"111011011",
11474=>"000011000",
11475=>"000000000",
11476=>"000000111",
11477=>"110000100",
11478=>"000011011",
11479=>"100000011",
11480=>"110011011",
11481=>"000000001",
11482=>"100101000",
11483=>"111100101",
11484=>"011110111",
11485=>"101101110",
11486=>"010111111",
11487=>"000000000",
11488=>"000000000",
11489=>"101100100",
11490=>"111101000",
11491=>"101111101",
11492=>"111000000",
11493=>"000000100",
11494=>"101101101",
11495=>"010111100",
11496=>"101111000",
11497=>"110000000",
11498=>"001111010",
11499=>"100010111",
11500=>"011000000",
11501=>"111001001",
11502=>"000000000",
11503=>"101000000",
11504=>"101100100",
11505=>"011011011",
11506=>"001001110",
11507=>"010011111",
11508=>"011111111",
11509=>"101000001",
11510=>"100000000",
11511=>"010011100",
11512=>"010011000",
11513=>"001101011",
11514=>"111111111",
11515=>"000001011",
11516=>"101000000",
11517=>"000100000",
11518=>"001100001",
11519=>"001100101",
11520=>"111110110",
11521=>"111110011",
11522=>"000000101",
11523=>"011011001",
11524=>"000001100",
11525=>"000111111",
11526=>"010010010",
11527=>"000000000",
11528=>"000010011",
11529=>"100001000",
11530=>"110001000",
11531=>"111001011",
11532=>"111001000",
11533=>"000000010",
11534=>"010110011",
11535=>"000111110",
11536=>"011011101",
11537=>"101111111",
11538=>"101110000",
11539=>"001011000",
11540=>"000100100",
11541=>"100100100",
11542=>"000110011",
11543=>"101001101",
11544=>"000000001",
11545=>"100010110",
11546=>"111111110",
11547=>"000000110",
11548=>"000100110",
11549=>"111000110",
11550=>"000100100",
11551=>"010010000",
11552=>"011000001",
11553=>"011010110",
11554=>"000000101",
11555=>"101000111",
11556=>"101011111",
11557=>"000011011",
11558=>"101000100",
11559=>"111111111",
11560=>"011101101",
11561=>"101111111",
11562=>"100000011",
11563=>"110010010",
11564=>"110011011",
11565=>"000010010",
11566=>"000000100",
11567=>"000111111",
11568=>"000000111",
11569=>"000110010",
11570=>"111111110",
11571=>"000000101",
11572=>"010111110",
11573=>"010100011",
11574=>"000001011",
11575=>"110100111",
11576=>"010000100",
11577=>"000001000",
11578=>"000111000",
11579=>"000000000",
11580=>"000001111",
11581=>"111111111",
11582=>"000100000",
11583=>"100101000",
11584=>"111011011",
11585=>"000000101",
11586=>"010100100",
11587=>"000000110",
11588=>"111111111",
11589=>"000000101",
11590=>"101001011",
11591=>"111011111",
11592=>"000111001",
11593=>"001011001",
11594=>"111111100",
11595=>"111100000",
11596=>"100100111",
11597=>"000111111",
11598=>"000011011",
11599=>"001011111",
11600=>"100000100",
11601=>"111111111",
11602=>"000000011",
11603=>"110111001",
11604=>"000100000",
11605=>"001111111",
11606=>"000100011",
11607=>"000111111",
11608=>"000011010",
11609=>"000110011",
11610=>"010010010",
11611=>"010000110",
11612=>"000011111",
11613=>"010110000",
11614=>"101000000",
11615=>"101101011",
11616=>"100100000",
11617=>"000000000",
11618=>"000111011",
11619=>"011111000",
11620=>"111111100",
11621=>"000101010",
11622=>"000010010",
11623=>"000000000",
11624=>"111010100",
11625=>"000000000",
11626=>"111111000",
11627=>"111111111",
11628=>"100100100",
11629=>"000011010",
11630=>"000010000",
11631=>"100111000",
11632=>"000110110",
11633=>"111000000",
11634=>"000110100",
11635=>"000110110",
11636=>"101000000",
11637=>"010010011",
11638=>"100111101",
11639=>"100000000",
11640=>"011011011",
11641=>"001011010",
11642=>"000011000",
11643=>"111000111",
11644=>"011101001",
11645=>"011011000",
11646=>"001001000",
11647=>"000000110",
11648=>"111110110",
11649=>"000011110",
11650=>"000011011",
11651=>"111100100",
11652=>"111010000",
11653=>"111111111",
11654=>"000110110",
11655=>"000101110",
11656=>"011011001",
11657=>"111000000",
11658=>"001011000",
11659=>"111111111",
11660=>"000000100",
11661=>"101101000",
11662=>"011000100",
11663=>"111000001",
11664=>"100100100",
11665=>"000000000",
11666=>"001011000",
11667=>"110011000",
11668=>"100000000",
11669=>"000000111",
11670=>"101100110",
11671=>"110110101",
11672=>"000100010",
11673=>"010111110",
11674=>"000010000",
11675=>"111010110",
11676=>"000000000",
11677=>"111000000",
11678=>"001001000",
11679=>"110000000",
11680=>"100110010",
11681=>"011010110",
11682=>"011101100",
11683=>"111011110",
11684=>"000111111",
11685=>"101101111",
11686=>"000000000",
11687=>"000010011",
11688=>"000100000",
11689=>"111111101",
11690=>"000000000",
11691=>"000110111",
11692=>"110100000",
11693=>"100101000",
11694=>"101001001",
11695=>"110001000",
11696=>"000100101",
11697=>"001110110",
11698=>"000000000",
11699=>"001011110",
11700=>"011001000",
11701=>"110001100",
11702=>"011011111",
11703=>"001111011",
11704=>"100100001",
11705=>"000000001",
11706=>"000011111",
11707=>"000010000",
11708=>"101101111",
11709=>"000111111",
11710=>"110110100",
11711=>"000000100",
11712=>"000111111",
11713=>"000111011",
11714=>"011000000",
11715=>"001001001",
11716=>"000101110",
11717=>"000100100",
11718=>"111111011",
11719=>"111011000",
11720=>"000100111",
11721=>"100100100",
11722=>"110101111",
11723=>"100000100",
11724=>"110100111",
11725=>"110111011",
11726=>"000111010",
11727=>"111111000",
11728=>"010100101",
11729=>"101111110",
11730=>"110110100",
11731=>"100101111",
11732=>"000000000",
11733=>"010011011",
11734=>"000111011",
11735=>"110000000",
11736=>"001101100",
11737=>"100000000",
11738=>"000001110",
11739=>"111111111",
11740=>"110111110",
11741=>"110110111",
11742=>"010111010",
11743=>"000000010",
11744=>"000100000",
11745=>"010000001",
11746=>"110111111",
11747=>"110111011",
11748=>"111000000",
11749=>"101000101",
11750=>"111011111",
11751=>"000000100",
11752=>"111011111",
11753=>"101100000",
11754=>"111101000",
11755=>"101111111",
11756=>"101111101",
11757=>"000000111",
11758=>"100111001",
11759=>"110001111",
11760=>"111101111",
11761=>"111001000",
11762=>"011100110",
11763=>"011011010",
11764=>"011011011",
11765=>"111100110",
11766=>"000010111",
11767=>"000000000",
11768=>"010111101",
11769=>"001000000",
11770=>"110010011",
11771=>"111111000",
11772=>"100000000",
11773=>"101000100",
11774=>"000111111",
11775=>"111100100",
11776=>"110111111",
11777=>"000000000",
11778=>"100000100",
11779=>"000000001",
11780=>"111101011",
11781=>"001000101",
11782=>"010110111",
11783=>"000101101",
11784=>"010010010",
11785=>"001100111",
11786=>"000000000",
11787=>"000010100",
11788=>"010110011",
11789=>"000000100",
11790=>"100000010",
11791=>"000100000",
11792=>"100001001",
11793=>"000001101",
11794=>"111011011",
11795=>"000000111",
11796=>"111100000",
11797=>"010010010",
11798=>"000000001",
11799=>"000000001",
11800=>"101000000",
11801=>"111111110",
11802=>"000000001",
11803=>"111001000",
11804=>"101111101",
11805=>"001111111",
11806=>"001101001",
11807=>"111110111",
11808=>"010010000",
11809=>"000000000",
11810=>"000010100",
11811=>"000000000",
11812=>"111011011",
11813=>"110010011",
11814=>"001111000",
11815=>"000010111",
11816=>"010010010",
11817=>"001111101",
11818=>"010000010",
11819=>"000010010",
11820=>"110111111",
11821=>"111001111",
11822=>"001001101",
11823=>"010010111",
11824=>"000111111",
11825=>"001001111",
11826=>"000010000",
11827=>"111111011",
11828=>"000001110",
11829=>"000000000",
11830=>"011010101",
11831=>"101101001",
11832=>"001100001",
11833=>"100001101",
11834=>"100111011",
11835=>"000000000",
11836=>"001001100",
11837=>"111111100",
11838=>"000101000",
11839=>"110100101",
11840=>"101101010",
11841=>"110101111",
11842=>"001101111",
11843=>"110010011",
11844=>"010101101",
11845=>"000001001",
11846=>"111111111",
11847=>"000000000",
11848=>"011000111",
11849=>"110101000",
11850=>"000101111",
11851=>"001001101",
11852=>"001000000",
11853=>"111111111",
11854=>"100100111",
11855=>"010000001",
11856=>"111111000",
11857=>"110111111",
11858=>"010011111",
11859=>"111011011",
11860=>"000100000",
11861=>"111011110",
11862=>"110010010",
11863=>"101000101",
11864=>"111111100",
11865=>"011011110",
11866=>"001000000",
11867=>"100001001",
11868=>"010111111",
11869=>"011001110",
11870=>"111110111",
11871=>"011110110",
11872=>"001101100",
11873=>"111111000",
11874=>"101100100",
11875=>"000000000",
11876=>"011000000",
11877=>"110111111",
11878=>"010010010",
11879=>"101000010",
11880=>"101001000",
11881=>"001000101",
11882=>"000000100",
11883=>"000100101",
11884=>"000101111",
11885=>"010101111",
11886=>"001000001",
11887=>"111111010",
11888=>"100100111",
11889=>"000000111",
11890=>"110110111",
11891=>"111110111",
11892=>"011011001",
11893=>"000101001",
11894=>"101111111",
11895=>"100110111",
11896=>"010111000",
11897=>"000000000",
11898=>"110011111",
11899=>"111110100",
11900=>"111010000",
11901=>"110100010",
11902=>"010110000",
11903=>"110010010",
11904=>"000001000",
11905=>"110100000",
11906=>"000000010",
11907=>"000000000",
11908=>"000101001",
11909=>"111111111",
11910=>"010110100",
11911=>"011111010",
11912=>"001110111",
11913=>"000001101",
11914=>"000000101",
11915=>"100001001",
11916=>"100111110",
11917=>"011100000",
11918=>"110010000",
11919=>"101101000",
11920=>"111111011",
11921=>"011000000",
11922=>"000001001",
11923=>"000111011",
11924=>"100000000",
11925=>"000101101",
11926=>"010111011",
11927=>"100111110",
11928=>"011000101",
11929=>"010110101",
11930=>"010010010",
11931=>"010010000",
11932=>"001000101",
11933=>"000001000",
11934=>"000001101",
11935=>"101101110",
11936=>"011011011",
11937=>"000000000",
11938=>"010111110",
11939=>"000100110",
11940=>"001101111",
11941=>"110110111",
11942=>"101001001",
11943=>"010000101",
11944=>"111000001",
11945=>"000000000",
11946=>"101101101",
11947=>"101001001",
11948=>"110100101",
11949=>"110100011",
11950=>"011000001",
11951=>"000011011",
11952=>"000000000",
11953=>"110110101",
11954=>"000101000",
11955=>"100010011",
11956=>"111011111",
11957=>"100101101",
11958=>"000101111",
11959=>"001001000",
11960=>"110100011",
11961=>"100010011",
11962=>"000000000",
11963=>"111101111",
11964=>"111111111",
11965=>"111110101",
11966=>"001000010",
11967=>"000000001",
11968=>"110011011",
11969=>"011111011",
11970=>"101000000",
11971=>"010011111",
11972=>"000010000",
11973=>"001101100",
11974=>"000000100",
11975=>"100111111",
11976=>"010010111",
11977=>"101011010",
11978=>"000000000",
11979=>"011101110",
11980=>"110010010",
11981=>"111011011",
11982=>"101101000",
11983=>"101000000",
11984=>"100101111",
11985=>"110111111",
11986=>"100000000",
11987=>"110100110",
11988=>"011010101",
11989=>"000000001",
11990=>"111110000",
11991=>"000001101",
11992=>"010010111",
11993=>"000000000",
11994=>"100110010",
11995=>"101101101",
11996=>"000111011",
11997=>"001000101",
11998=>"111010111",
11999=>"100100111",
12000=>"000000111",
12001=>"001110101",
12002=>"111110111",
12003=>"001000111",
12004=>"101001000",
12005=>"001011010",
12006=>"000010001",
12007=>"000001000",
12008=>"000000101",
12009=>"010011111",
12010=>"111001000",
12011=>"111110011",
12012=>"010010010",
12013=>"000001101",
12014=>"001101010",
12015=>"000010010",
12016=>"101000001",
12017=>"100000001",
12018=>"000000010",
12019=>"110110110",
12020=>"011011011",
12021=>"010000101",
12022=>"000101001",
12023=>"011111111",
12024=>"000001001",
12025=>"000000101",
12026=>"111011010",
12027=>"000001001",
12028=>"010111000",
12029=>"111011011",
12030=>"011010110",
12031=>"111111111",
12032=>"101100101",
12033=>"000000000",
12034=>"000000100",
12035=>"000001101",
12036=>"000011000",
12037=>"010000101",
12038=>"101111111",
12039=>"010011101",
12040=>"000001001",
12041=>"111110100",
12042=>"000011011",
12043=>"000000010",
12044=>"101000000",
12045=>"001000000",
12046=>"111111100",
12047=>"011001010",
12048=>"010111011",
12049=>"011000000",
12050=>"000011110",
12051=>"010111101",
12052=>"001100110",
12053=>"111111000",
12054=>"011011101",
12055=>"000111111",
12056=>"101000000",
12057=>"111110000",
12058=>"000000000",
12059=>"000010110",
12060=>"000000110",
12061=>"000110111",
12062=>"000000000",
12063=>"000011010",
12064=>"000100111",
12065=>"000010110",
12066=>"000001101",
12067=>"100111111",
12068=>"100100111",
12069=>"110010111",
12070=>"000011011",
12071=>"000111000",
12072=>"001011111",
12073=>"111000111",
12074=>"010100000",
12075=>"101001000",
12076=>"100110110",
12077=>"010001000",
12078=>"011110000",
12079=>"111111111",
12080=>"111100100",
12081=>"010001111",
12082=>"000101100",
12083=>"000001001",
12084=>"000000011",
12085=>"111010000",
12086=>"011011111",
12087=>"000101001",
12088=>"000000111",
12089=>"000000010",
12090=>"000001111",
12091=>"000000110",
12092=>"100100110",
12093=>"110010010",
12094=>"000000100",
12095=>"111011011",
12096=>"110111111",
12097=>"001100111",
12098=>"010111111",
12099=>"011000110",
12100=>"010011010",
12101=>"000101101",
12102=>"000101000",
12103=>"001000111",
12104=>"010011010",
12105=>"101000000",
12106=>"001111001",
12107=>"011000000",
12108=>"000000111",
12109=>"011001001",
12110=>"000110011",
12111=>"000000011",
12112=>"000101111",
12113=>"111111010",
12114=>"111111111",
12115=>"011000001",
12116=>"101000000",
12117=>"010011011",
12118=>"011111110",
12119=>"001111011",
12120=>"111100000",
12121=>"000011111",
12122=>"111101000",
12123=>"000100100",
12124=>"111000000",
12125=>"011000000",
12126=>"111111100",
12127=>"100111111",
12128=>"100100000",
12129=>"111101010",
12130=>"101000100",
12131=>"001011101",
12132=>"001000000",
12133=>"010010000",
12134=>"111111111",
12135=>"111000000",
12136=>"111111010",
12137=>"010111111",
12138=>"111000000",
12139=>"111000000",
12140=>"000010010",
12141=>"111101000",
12142=>"000111100",
12143=>"000111010",
12144=>"011011011",
12145=>"000010110",
12146=>"110011111",
12147=>"000101000",
12148=>"000000010",
12149=>"001000010",
12150=>"010110000",
12151=>"101101001",
12152=>"011111111",
12153=>"111000111",
12154=>"000000000",
12155=>"111011000",
12156=>"000011111",
12157=>"111100000",
12158=>"101111100",
12159=>"000000011",
12160=>"101000000",
12161=>"111111111",
12162=>"110000001",
12163=>"000100101",
12164=>"010000110",
12165=>"001000101",
12166=>"111111011",
12167=>"000100100",
12168=>"100110111",
12169=>"110111000",
12170=>"111111100",
12171=>"100000111",
12172=>"111000000",
12173=>"111100100",
12174=>"010101001",
12175=>"001001010",
12176=>"001011011",
12177=>"011011000",
12178=>"000111111",
12179=>"000100000",
12180=>"111110000",
12181=>"000110111",
12182=>"010000010",
12183=>"011011111",
12184=>"100111100",
12185=>"110001100",
12186=>"111000111",
12187=>"000000000",
12188=>"100010111",
12189=>"111111000",
12190=>"000000000",
12191=>"000001000",
12192=>"011100100",
12193=>"111101111",
12194=>"010000000",
12195=>"011000000",
12196=>"010011000",
12197=>"100001110",
12198=>"001001111",
12199=>"001010011",
12200=>"000000100",
12201=>"011000000",
12202=>"101001000",
12203=>"000010110",
12204=>"101111111",
12205=>"000000000",
12206=>"000000111",
12207=>"111101001",
12208=>"111011000",
12209=>"111001001",
12210=>"000000000",
12211=>"100110011",
12212=>"011111110",
12213=>"111000100",
12214=>"101000000",
12215=>"111111000",
12216=>"101010011",
12217=>"011001000",
12218=>"111010111",
12219=>"111001100",
12220=>"011000000",
12221=>"111111011",
12222=>"110111001",
12223=>"000000000",
12224=>"010100111",
12225=>"000000000",
12226=>"010010011",
12227=>"011011110",
12228=>"000101100",
12229=>"010001101",
12230=>"000111000",
12231=>"111111000",
12232=>"111111100",
12233=>"000011101",
12234=>"111000000",
12235=>"011000001",
12236=>"111110110",
12237=>"000101111",
12238=>"001110111",
12239=>"011001110",
12240=>"000010101",
12241=>"111110110",
12242=>"110000000",
12243=>"110100100",
12244=>"111000000",
12245=>"001100111",
12246=>"000010010",
12247=>"111100000",
12248=>"000000101",
12249=>"000011111",
12250=>"000100011",
12251=>"111101000",
12252=>"110111011",
12253=>"000101111",
12254=>"111101100",
12255=>"000110001",
12256=>"000011010",
12257=>"101000000",
12258=>"000111000",
12259=>"111001001",
12260=>"010000000",
12261=>"111000000",
12262=>"111010000",
12263=>"000101110",
12264=>"000101110",
12265=>"111000010",
12266=>"000000110",
12267=>"011001001",
12268=>"111111010",
12269=>"001111111",
12270=>"110000000",
12271=>"101000000",
12272=>"010010111",
12273=>"011110110",
12274=>"010000000",
12275=>"000011110",
12276=>"101011001",
12277=>"111111000",
12278=>"000000000",
12279=>"010000000",
12280=>"000001111",
12281=>"001111000",
12282=>"000010010",
12283=>"101111010",
12284=>"111000000",
12285=>"111001000",
12286=>"010110010",
12287=>"000110000",
12288=>"011011000",
12289=>"001000111",
12290=>"101000000",
12291=>"100000111",
12292=>"000100100",
12293=>"110000001",
12294=>"010111111",
12295=>"001011010",
12296=>"000000101",
12297=>"000000000",
12298=>"011111010",
12299=>"000111010",
12300=>"010010010",
12301=>"100000000",
12302=>"000011011",
12303=>"101110000",
12304=>"011000101",
12305=>"001100000",
12306=>"111101001",
12307=>"000010010",
12308=>"011101111",
12309=>"101000001",
12310=>"101101001",
12311=>"110101110",
12312=>"100001111",
12313=>"101111001",
12314=>"010100000",
12315=>"000011111",
12316=>"110000001",
12317=>"001100110",
12318=>"111010001",
12319=>"000000000",
12320=>"111101101",
12321=>"111101110",
12322=>"110010010",
12323=>"010010010",
12324=>"100111001",
12325=>"110110001",
12326=>"001000000",
12327=>"101000111",
12328=>"111101111",
12329=>"001011111",
12330=>"011011000",
12331=>"111101111",
12332=>"110111111",
12333=>"111111110",
12334=>"111001001",
12335=>"000100110",
12336=>"100101000",
12337=>"111101101",
12338=>"010000000",
12339=>"001000101",
12340=>"011010000",
12341=>"001110111",
12342=>"110000001",
12343=>"010110101",
12344=>"010000111",
12345=>"000101111",
12346=>"011001000",
12347=>"000111011",
12348=>"001110011",
12349=>"111111111",
12350=>"101001111",
12351=>"000011111",
12352=>"000010111",
12353=>"101111101",
12354=>"000100111",
12355=>"001000010",
12356=>"000101000",
12357=>"111101101",
12358=>"000111010",
12359=>"111010000",
12360=>"111001111",
12361=>"011000111",
12362=>"111000111",
12363=>"101101100",
12364=>"100000000",
12365=>"011101101",
12366=>"100101101",
12367=>"010111111",
12368=>"000100100",
12369=>"111001111",
12370=>"110001010",
12371=>"011001100",
12372=>"000000000",
12373=>"001111111",
12374=>"001101101",
12375=>"111000001",
12376=>"111111000",
12377=>"000100111",
12378=>"101111100",
12379=>"110100100",
12380=>"001000001",
12381=>"010001001",
12382=>"111110001",
12383=>"100000101",
12384=>"011111010",
12385=>"111100101",
12386=>"000111110",
12387=>"001001101",
12388=>"001111001",
12389=>"000101111",
12390=>"000101111",
12391=>"000000101",
12392=>"101000011",
12393=>"011011101",
12394=>"010011110",
12395=>"000000000",
12396=>"111000101",
12397=>"000111000",
12398=>"001010010",
12399=>"111001000",
12400=>"000111001",
12401=>"000111111",
12402=>"011001100",
12403=>"000011000",
12404=>"111100000",
12405=>"000000101",
12406=>"000000111",
12407=>"000111000",
12408=>"011010111",
12409=>"111111000",
12410=>"001001000",
12411=>"100000000",
12412=>"000110110",
12413=>"110100000",
12414=>"110000000",
12415=>"000000000",
12416=>"000101100",
12417=>"001000000",
12418=>"101000111",
12419=>"001000000",
12420=>"111001011",
12421=>"000000001",
12422=>"111111100",
12423=>"000000100",
12424=>"110100000",
12425=>"001000000",
12426=>"000100000",
12427=>"111010000",
12428=>"001000100",
12429=>"111111100",
12430=>"110111111",
12431=>"100001101",
12432=>"111110101",
12433=>"101111010",
12434=>"000001111",
12435=>"111000100",
12436=>"101011001",
12437=>"000000001",
12438=>"100111111",
12439=>"010001011",
12440=>"000111110",
12441=>"010000000",
12442=>"010011000",
12443=>"000010000",
12444=>"111011011",
12445=>"001111001",
12446=>"000000011",
12447=>"000001000",
12448=>"111101011",
12449=>"101000000",
12450=>"010000000",
12451=>"111010010",
12452=>"000001111",
12453=>"110010101",
12454=>"000000001",
12455=>"001111110",
12456=>"000000001",
12457=>"100000000",
12458=>"111101101",
12459=>"011000000",
12460=>"001100000",
12461=>"101001111",
12462=>"111100011",
12463=>"000010111",
12464=>"110000111",
12465=>"010101100",
12466=>"111001101",
12467=>"001100111",
12468=>"001001101",
12469=>"011111010",
12470=>"001001110",
12471=>"000011100",
12472=>"000010010",
12473=>"000110110",
12474=>"000010010",
12475=>"111011000",
12476=>"010010010",
12477=>"111110000",
12478=>"101000000",
12479=>"110000100",
12480=>"100001101",
12481=>"000011111",
12482=>"110000000",
12483=>"000011100",
12484=>"100111000",
12485=>"101100101",
12486=>"111110111",
12487=>"111111111",
12488=>"111111111",
12489=>"000000000",
12490=>"111011111",
12491=>"000111000",
12492=>"100100001",
12493=>"000011011",
12494=>"010001001",
12495=>"100000011",
12496=>"110000000",
12497=>"001111000",
12498=>"010000111",
12499=>"101101101",
12500=>"000101111",
12501=>"010111110",
12502=>"000001001",
12503=>"110110000",
12504=>"000111000",
12505=>"000000101",
12506=>"111001100",
12507=>"000000000",
12508=>"001001111",
12509=>"110000000",
12510=>"000001101",
12511=>"000010101",
12512=>"101101111",
12513=>"111000000",
12514=>"101000100",
12515=>"001100000",
12516=>"101100101",
12517=>"000110110",
12518=>"101011110",
12519=>"111001000",
12520=>"010001111",
12521=>"100100010",
12522=>"110011011",
12523=>"000010000",
12524=>"000000000",
12525=>"001110001",
12526=>"000110000",
12527=>"000000000",
12528=>"010110010",
12529=>"101011111",
12530=>"110010100",
12531=>"001001001",
12532=>"110110100",
12533=>"111000000",
12534=>"000000000",
12535=>"100000000",
12536=>"000001000",
12537=>"110111110",
12538=>"111111110",
12539=>"000100111",
12540=>"000000010",
12541=>"000000010",
12542=>"001111010",
12543=>"000110110",
12544=>"011011001",
12545=>"000000000",
12546=>"101000000",
12547=>"110000000",
12548=>"000100010",
12549=>"110110110",
12550=>"000010010",
12551=>"000010000",
12552=>"111111111",
12553=>"000000101",
12554=>"000000001",
12555=>"111110010",
12556=>"000000000",
12557=>"111111001",
12558=>"000101101",
12559=>"000000010",
12560=>"111111010",
12561=>"000000000",
12562=>"111111000",
12563=>"110101000",
12564=>"000001111",
12565=>"111110100",
12566=>"111011011",
12567=>"000111111",
12568=>"100000000",
12569=>"001010000",
12570=>"111111111",
12571=>"101111111",
12572=>"001111000",
12573=>"111011110",
12574=>"001001110",
12575=>"110011001",
12576=>"011000000",
12577=>"000001110",
12578=>"000000000",
12579=>"110010111",
12580=>"011111011",
12581=>"010001001",
12582=>"110110000",
12583=>"001111111",
12584=>"000000000",
12585=>"110111111",
12586=>"000010010",
12587=>"101010000",
12588=>"111111010",
12589=>"110100011",
12590=>"000001111",
12591=>"001001000",
12592=>"111001011",
12593=>"001011110",
12594=>"011010000",
12595=>"011000000",
12596=>"000000000",
12597=>"000000000",
12598=>"111101111",
12599=>"000101001",
12600=>"011000111",
12601=>"010011011",
12602=>"000000000",
12603=>"000000010",
12604=>"111110011",
12605=>"010111011",
12606=>"000000000",
12607=>"111111111",
12608=>"110011010",
12609=>"101101101",
12610=>"010111111",
12611=>"000001111",
12612=>"000100000",
12613=>"000000000",
12614=>"000010111",
12615=>"010110000",
12616=>"111111111",
12617=>"001111111",
12618=>"111010111",
12619=>"000001000",
12620=>"111111111",
12621=>"010110110",
12622=>"101000110",
12623=>"111101010",
12624=>"111111101",
12625=>"111111011",
12626=>"010001001",
12627=>"111001001",
12628=>"000000010",
12629=>"011111001",
12630=>"111111111",
12631=>"101000111",
12632=>"010110000",
12633=>"001111111",
12634=>"010110100",
12635=>"000011011",
12636=>"001101101",
12637=>"001001001",
12638=>"000000000",
12639=>"111100011",
12640=>"110110110",
12641=>"111111111",
12642=>"000000000",
12643=>"111011011",
12644=>"010110100",
12645=>"101000010",
12646=>"111111101",
12647=>"000000000",
12648=>"111011010",
12649=>"000000110",
12650=>"000111110",
12651=>"110111111",
12652=>"111011110",
12653=>"000000000",
12654=>"011111001",
12655=>"000101101",
12656=>"001101100",
12657=>"001001111",
12658=>"110111111",
12659=>"000000110",
12660=>"011100010",
12661=>"000000001",
12662=>"010000111",
12663=>"000000000",
12664=>"000011001",
12665=>"111011110",
12666=>"011000000",
12667=>"011111110",
12668=>"010111111",
12669=>"110100100",
12670=>"101101000",
12671=>"101100111",
12672=>"100001001",
12673=>"111111010",
12674=>"011111011",
12675=>"000011010",
12676=>"110100101",
12677=>"000011111",
12678=>"000001001",
12679=>"111100010",
12680=>"111111000",
12681=>"001001000",
12682=>"000000100",
12683=>"000000001",
12684=>"111000000",
12685=>"010110010",
12686=>"001001000",
12687=>"001000000",
12688=>"100101100",
12689=>"110100110",
12690=>"010110101",
12691=>"111000000",
12692=>"111000010",
12693=>"100000100",
12694=>"000001001",
12695=>"111111111",
12696=>"000000000",
12697=>"000000000",
12698=>"111111000",
12699=>"000000000",
12700=>"001010111",
12701=>"010000010",
12702=>"111000011",
12703=>"000010011",
12704=>"100111110",
12705=>"001000000",
12706=>"000010001",
12707=>"000000010",
12708=>"011011010",
12709=>"110110110",
12710=>"000000100",
12711=>"000000000",
12712=>"000000000",
12713=>"101001111",
12714=>"111111000",
12715=>"100000000",
12716=>"000000001",
12717=>"110000000",
12718=>"110100001",
12719=>"000000110",
12720=>"110000111",
12721=>"011011011",
12722=>"110101000",
12723=>"001001100",
12724=>"010011011",
12725=>"000000000",
12726=>"011000010",
12727=>"000000100",
12728=>"110000111",
12729=>"111011000",
12730=>"001010000",
12731=>"010011001",
12732=>"000011101",
12733=>"111111111",
12734=>"111111111",
12735=>"001011101",
12736=>"000000000",
12737=>"001000001",
12738=>"110010110",
12739=>"111001110",
12740=>"000010000",
12741=>"111011000",
12742=>"111011110",
12743=>"100100100",
12744=>"000000000",
12745=>"111110010",
12746=>"000100111",
12747=>"100000011",
12748=>"101000000",
12749=>"110110101",
12750=>"000000110",
12751=>"111011000",
12752=>"011111010",
12753=>"110110110",
12754=>"111011000",
12755=>"111111011",
12756=>"000000000",
12757=>"100000000",
12758=>"110111101",
12759=>"110010110",
12760=>"010010010",
12761=>"110100000",
12762=>"011111010",
12763=>"000000000",
12764=>"111001000",
12765=>"010011000",
12766=>"001101001",
12767=>"111111111",
12768=>"000010000",
12769=>"000000001",
12770=>"000000000",
12771=>"111101011",
12772=>"000000000",
12773=>"110111111",
12774=>"011011000",
12775=>"011000000",
12776=>"000000111",
12777=>"000000000",
12778=>"000000000",
12779=>"000000000",
12780=>"101010110",
12781=>"000100010",
12782=>"111010000",
12783=>"111000010",
12784=>"110011000",
12785=>"110100000",
12786=>"111111111",
12787=>"110111111",
12788=>"011100100",
12789=>"101101100",
12790=>"000000000",
12791=>"101111011",
12792=>"101111111",
12793=>"110110010",
12794=>"111111111",
12795=>"010111100",
12796=>"000110111",
12797=>"000000000",
12798=>"110111111",
12799=>"000100111",
12800=>"001001111",
12801=>"111011110",
12802=>"001000001",
12803=>"111111011",
12804=>"000110001",
12805=>"100110110",
12806=>"000110000",
12807=>"110000111",
12808=>"010111101",
12809=>"100100101",
12810=>"011010000",
12811=>"111001101",
12812=>"100000010",
12813=>"111111011",
12814=>"001011111",
12815=>"111110010",
12816=>"111100111",
12817=>"100110100",
12818=>"011010110",
12819=>"100010000",
12820=>"100100011",
12821=>"111111110",
12822=>"011011010",
12823=>"000011000",
12824=>"000010111",
12825=>"001110011",
12826=>"001010000",
12827=>"001011111",
12828=>"000000000",
12829=>"100001001",
12830=>"001001001",
12831=>"011011011",
12832=>"011100001",
12833=>"111101011",
12834=>"100100100",
12835=>"000110110",
12836=>"101011011",
12837=>"000000001",
12838=>"001001011",
12839=>"011100010",
12840=>"000101111",
12841=>"000001111",
12842=>"011000000",
12843=>"100110110",
12844=>"001001101",
12845=>"001011100",
12846=>"100011011",
12847=>"000100000",
12848=>"010110100",
12849=>"011111000",
12850=>"001100100",
12851=>"111100100",
12852=>"011001111",
12853=>"011111101",
12854=>"100111111",
12855=>"001011000",
12856=>"111101111",
12857=>"011001011",
12858=>"111000010",
12859=>"010110110",
12860=>"001101001",
12861=>"011011010",
12862=>"000000000",
12863=>"101001000",
12864=>"011100000",
12865=>"000000011",
12866=>"010010000",
12867=>"011001001",
12868=>"110010110",
12869=>"010000111",
12870=>"001000000",
12871=>"111101011",
12872=>"111001011",
12873=>"110100101",
12874=>"011001011",
12875=>"001011001",
12876=>"111000111",
12877=>"001000000",
12878=>"001001011",
12879=>"011100111",
12880=>"011011011",
12881=>"000001101",
12882=>"010000000",
12883=>"010011111",
12884=>"100000000",
12885=>"011110001",
12886=>"001001101",
12887=>"100100100",
12888=>"010011010",
12889=>"011011010",
12890=>"000001000",
12891=>"111111111",
12892=>"000110100",
12893=>"110000100",
12894=>"100111110",
12895=>"011101111",
12896=>"010010000",
12897=>"011100001",
12898=>"000000001",
12899=>"011111001",
12900=>"101101111",
12901=>"001011000",
12902=>"000100101",
12903=>"011001111",
12904=>"111101011",
12905=>"110110100",
12906=>"111011001",
12907=>"001011000",
12908=>"000001111",
12909=>"110110110",
12910=>"111110000",
12911=>"010000000",
12912=>"000000010",
12913=>"111111100",
12914=>"010010100",
12915=>"111110111",
12916=>"100101001",
12917=>"011001001",
12918=>"011001000",
12919=>"110110000",
12920=>"100000100",
12921=>"100000110",
12922=>"000110100",
12923=>"110110100",
12924=>"000000100",
12925=>"100000111",
12926=>"100111001",
12927=>"001001001",
12928=>"011001000",
12929=>"111001001",
12930=>"110100100",
12931=>"110111101",
12932=>"001111100",
12933=>"011000011",
12934=>"011011001",
12935=>"001110111",
12936=>"111111111",
12937=>"010101001",
12938=>"110000000",
12939=>"110100110",
12940=>"100100100",
12941=>"100100010",
12942=>"001011100",
12943=>"000000000",
12944=>"011001010",
12945=>"001011111",
12946=>"001110010",
12947=>"001011111",
12948=>"001101101",
12949=>"100100110",
12950=>"011011001",
12951=>"001000001",
12952=>"000000000",
12953=>"111000000",
12954=>"000001000",
12955=>"110110110",
12956=>"000010000",
12957=>"001001101",
12958=>"011000001",
12959=>"001001001",
12960=>"111011111",
12961=>"010111010",
12962=>"100010110",
12963=>"011001111",
12964=>"111111010",
12965=>"000000000",
12966=>"110100000",
12967=>"100100100",
12968=>"010100110",
12969=>"011111110",
12970=>"100100111",
12971=>"000000111",
12972=>"000110000",
12973=>"001001001",
12974=>"001011000",
12975=>"110100111",
12976=>"101000000",
12977=>"100100100",
12978=>"010111100",
12979=>"011000000",
12980=>"111111111",
12981=>"111011000",
12982=>"111111111",
12983=>"100110011",
12984=>"010110000",
12985=>"000000011",
12986=>"000011101",
12987=>"001100000",
12988=>"100101111",
12989=>"100110110",
12990=>"111010111",
12991=>"100100100",
12992=>"001011101",
12993=>"000001000",
12994=>"001011011",
12995=>"111011000",
12996=>"110110100",
12997=>"000001001",
12998=>"100100110",
12999=>"111000011",
13000=>"100100111",
13001=>"011011011",
13002=>"100100000",
13003=>"011001000",
13004=>"011001000",
13005=>"001011110",
13006=>"011001000",
13007=>"000100100",
13008=>"000001000",
13009=>"111011110",
13010=>"011100101",
13011=>"001111001",
13012=>"001001011",
13013=>"100110111",
13014=>"001001111",
13015=>"000001011",
13016=>"111011000",
13017=>"100100110",
13018=>"000100000",
13019=>"100100100",
13020=>"011011111",
13021=>"110111110",
13022=>"001000000",
13023=>"000011111",
13024=>"001111001",
13025=>"101100001",
13026=>"100100000",
13027=>"001001101",
13028=>"000000000",
13029=>"110111110",
13030=>"001001001",
13031=>"111011011",
13032=>"100110011",
13033=>"110000100",
13034=>"000110111",
13035=>"110111111",
13036=>"110110100",
13037=>"101110000",
13038=>"000100100",
13039=>"100001000",
13040=>"011011000",
13041=>"011111111",
13042=>"011011001",
13043=>"000000100",
13044=>"000000000",
13045=>"100000110",
13046=>"000000010",
13047=>"100100000",
13048=>"111110110",
13049=>"110100000",
13050=>"111111011",
13051=>"000000110",
13052=>"111001011",
13053=>"100110000",
13054=>"111001011",
13055=>"001001001",
13056=>"110010000",
13057=>"000110000",
13058=>"001001111",
13059=>"000000000",
13060=>"100110110",
13061=>"101001100",
13062=>"110110000",
13063=>"000110110",
13064=>"010011110",
13065=>"000111000",
13066=>"010010011",
13067=>"000001001",
13068=>"110110110",
13069=>"110000000",
13070=>"110110000",
13071=>"100110000",
13072=>"011000100",
13073=>"001000001",
13074=>"001001000",
13075=>"111111111",
13076=>"111111111",
13077=>"001001000",
13078=>"010101011",
13079=>"111111000",
13080=>"000000001",
13081=>"111111111",
13082=>"010000000",
13083=>"000000011",
13084=>"101001001",
13085=>"010111111",
13086=>"110100000",
13087=>"000110110",
13088=>"111001101",
13089=>"011001111",
13090=>"000110110",
13091=>"110111110",
13092=>"100000000",
13093=>"100100000",
13094=>"000000110",
13095=>"100110100",
13096=>"011001000",
13097=>"110111011",
13098=>"110000000",
13099=>"001000011",
13100=>"000000000",
13101=>"001111111",
13102=>"111110000",
13103=>"110111111",
13104=>"000001000",
13105=>"011011000",
13106=>"111011111",
13107=>"111001000",
13108=>"000010000",
13109=>"010011111",
13110=>"110100000",
13111=>"000011100",
13112=>"111110100",
13113=>"011011110",
13114=>"000101111",
13115=>"001111111",
13116=>"100000110",
13117=>"111111000",
13118=>"000000001",
13119=>"010111000",
13120=>"110111111",
13121=>"111110000",
13122=>"111000100",
13123=>"100100011",
13124=>"000001110",
13125=>"000110010",
13126=>"001000000",
13127=>"111001001",
13128=>"000110110",
13129=>"110110000",
13130=>"110000111",
13131=>"111110010",
13132=>"001001000",
13133=>"011001000",
13134=>"100100101",
13135=>"001010111",
13136=>"110000001",
13137=>"110000000",
13138=>"110000000",
13139=>"011011001",
13140=>"110110000",
13141=>"101110010",
13142=>"001111010",
13143=>"111110000",
13144=>"110111110",
13145=>"001011011",
13146=>"000111100",
13147=>"011111111",
13148=>"001000001",
13149=>"001001000",
13150=>"111001011",
13151=>"000111001",
13152=>"110110100",
13153=>"010100101",
13154=>"001000111",
13155=>"011010000",
13156=>"000000000",
13157=>"100001111",
13158=>"000110110",
13159=>"111011000",
13160=>"000110000",
13161=>"111000000",
13162=>"001111111",
13163=>"101000100",
13164=>"011000100",
13165=>"001010111",
13166=>"001001111",
13167=>"000111110",
13168=>"110111001",
13169=>"000010110",
13170=>"011001000",
13171=>"110110010",
13172=>"011000111",
13173=>"000000110",
13174=>"000110110",
13175=>"110110110",
13176=>"001000011",
13177=>"010010010",
13178=>"111001001",
13179=>"011001001",
13180=>"000100100",
13181=>"101000100",
13182=>"000000001",
13183=>"110110000",
13184=>"110111100",
13185=>"000111110",
13186=>"110000110",
13187=>"000101101",
13188=>"111110001",
13189=>"000001000",
13190=>"111011011",
13191=>"000101110",
13192=>"110001101",
13193=>"100100010",
13194=>"011001111",
13195=>"101011100",
13196=>"001001111",
13197=>"000000001",
13198=>"000000111",
13199=>"000000001",
13200=>"101000100",
13201=>"110110000",
13202=>"000100101",
13203=>"110101010",
13204=>"000111111",
13205=>"111001111",
13206=>"110101101",
13207=>"000010011",
13208=>"111111100",
13209=>"001010110",
13210=>"110110000",
13211=>"001110010",
13212=>"000100001",
13213=>"111001111",
13214=>"001001000",
13215=>"101000000",
13216=>"110100000",
13217=>"000000111",
13218=>"100100100",
13219=>"111100000",
13220=>"000001001",
13221=>"101100110",
13222=>"000110100",
13223=>"000000100",
13224=>"101011011",
13225=>"001100100",
13226=>"001000000",
13227=>"110000001",
13228=>"000110111",
13229=>"011000011",
13230=>"000001011",
13231=>"110000000",
13232=>"000100110",
13233=>"000000100",
13234=>"011010000",
13235=>"001100000",
13236=>"001011011",
13237=>"001111110",
13238=>"000111111",
13239=>"000110010",
13240=>"010001111",
13241=>"000100110",
13242=>"010011111",
13243=>"110000001",
13244=>"000010110",
13245=>"011001001",
13246=>"100000011",
13247=>"000001000",
13248=>"000110011",
13249=>"001000111",
13250=>"111101001",
13251=>"100110110",
13252=>"001000000",
13253=>"001001111",
13254=>"110101000",
13255=>"110110000",
13256=>"000010000",
13257=>"000110010",
13258=>"000000101",
13259=>"001001111",
13260=>"100111000",
13261=>"001111000",
13262=>"000000000",
13263=>"011001111",
13264=>"001011011",
13265=>"010110100",
13266=>"011110000",
13267=>"000000010",
13268=>"100100000",
13269=>"111000000",
13270=>"111001111",
13271=>"100000100",
13272=>"000000110",
13273=>"111111111",
13274=>"011110111",
13275=>"001011001",
13276=>"000001100",
13277=>"110111010",
13278=>"110111010",
13279=>"110110100",
13280=>"001000111",
13281=>"000000111",
13282=>"000111110",
13283=>"011111100",
13284=>"001000000",
13285=>"001000000",
13286=>"111001000",
13287=>"010011000",
13288=>"111111111",
13289=>"001000000",
13290=>"000010010",
13291=>"001100110",
13292=>"011110110",
13293=>"000000010",
13294=>"000000001",
13295=>"000000000",
13296=>"110111110",
13297=>"001000111",
13298=>"110110010",
13299=>"100000110",
13300=>"000101000",
13301=>"011111111",
13302=>"110010000",
13303=>"000110000",
13304=>"110111110",
13305=>"111110000",
13306=>"111010111",
13307=>"000110111",
13308=>"001000100",
13309=>"001001000",
13310=>"001001101",
13311=>"000000101",
13312=>"110110010",
13313=>"000001110",
13314=>"101101101",
13315=>"010010100",
13316=>"111110111",
13317=>"011011101",
13318=>"010000111",
13319=>"110011101",
13320=>"101001000",
13321=>"101101000",
13322=>"000001001",
13323=>"000100100",
13324=>"110101100",
13325=>"110000011",
13326=>"110100110",
13327=>"010111011",
13328=>"101001001",
13329=>"001111111",
13330=>"110010000",
13331=>"111010110",
13332=>"011000000",
13333=>"101101101",
13334=>"100110001",
13335=>"101101111",
13336=>"100100000",
13337=>"001001001",
13338=>"100011000",
13339=>"110110010",
13340=>"000000010",
13341=>"001000111",
13342=>"001000000",
13343=>"010010010",
13344=>"101001000",
13345=>"001000111",
13346=>"111100110",
13347=>"111101110",
13348=>"010010010",
13349=>"000000000",
13350=>"101100100",
13351=>"001101111",
13352=>"111011011",
13353=>"111011111",
13354=>"111110101",
13355=>"000001001",
13356=>"110110110",
13357=>"000000000",
13358=>"010100000",
13359=>"111011001",
13360=>"000000000",
13361=>"011010011",
13362=>"111001111",
13363=>"101111101",
13364=>"101111010",
13365=>"100010010",
13366=>"001000010",
13367=>"101100100",
13368=>"000111000",
13369=>"111000100",
13370=>"010010111",
13371=>"101111111",
13372=>"111010111",
13373=>"010010111",
13374=>"100101001",
13375=>"010000000",
13376=>"000001001",
13377=>"000010000",
13378=>"010000111",
13379=>"000100011",
13380=>"010000111",
13381=>"001001000",
13382=>"001001010",
13383=>"110110111",
13384=>"110010000",
13385=>"101001010",
13386=>"101000101",
13387=>"111111110",
13388=>"001101111",
13389=>"111010111",
13390=>"111111101",
13391=>"010001101",
13392=>"000000001",
13393=>"111000110",
13394=>"011000000",
13395=>"011010011",
13396=>"000111000",
13397=>"000001011",
13398=>"110010010",
13399=>"101101101",
13400=>"001011000",
13401=>"011010110",
13402=>"011010010",
13403=>"110110111",
13404=>"101100000",
13405=>"111010011",
13406=>"111101111",
13407=>"101100000",
13408=>"100100000",
13409=>"010010000",
13410=>"001101001",
13411=>"110110010",
13412=>"111111111",
13413=>"010010000",
13414=>"111001111",
13415=>"000000000",
13416=>"000000011",
13417=>"000001101",
13418=>"011100000",
13419=>"000001101",
13420=>"000000000",
13421=>"011111111",
13422=>"001000000",
13423=>"110010111",
13424=>"110110010",
13425=>"010000001",
13426=>"100000011",
13427=>"111111001",
13428=>"000001010",
13429=>"010010110",
13430=>"111000110",
13431=>"101000010",
13432=>"001000001",
13433=>"110010011",
13434=>"111111000",
13435=>"100000000",
13436=>"110010000",
13437=>"011010110",
13438=>"100000111",
13439=>"000000010",
13440=>"101101000",
13441=>"010000101",
13442=>"101000000",
13443=>"010110001",
13444=>"011000100",
13445=>"000100111",
13446=>"000000000",
13447=>"100100000",
13448=>"010010010",
13449=>"101100101",
13450=>"010010111",
13451=>"000001101",
13452=>"111000000",
13453=>"100001111",
13454=>"111111111",
13455=>"100100010",
13456=>"011010011",
13457=>"111110001",
13458=>"111000000",
13459=>"101000000",
13460=>"111001100",
13461=>"101101101",
13462=>"111111011",
13463=>"110110110",
13464=>"111000111",
13465=>"000001101",
13466=>"101000110",
13467=>"101001101",
13468=>"000110010",
13469=>"101100101",
13470=>"000101110",
13471=>"000001000",
13472=>"001100010",
13473=>"000101001",
13474=>"011000001",
13475=>"110111000",
13476=>"010110001",
13477=>"111011111",
13478=>"010110010",
13479=>"110011111",
13480=>"101101101",
13481=>"000001001",
13482=>"110110110",
13483=>"100101111",
13484=>"010000000",
13485=>"110010010",
13486=>"011010110",
13487=>"111101111",
13488=>"100100000",
13489=>"110110010",
13490=>"111011111",
13491=>"000001001",
13492=>"011010110",
13493=>"010010111",
13494=>"111101000",
13495=>"010010101",
13496=>"110000111",
13497=>"100000000",
13498=>"010010011",
13499=>"001000000",
13500=>"111000011",
13501=>"100101100",
13502=>"110000100",
13503=>"001001001",
13504=>"101001000",
13505=>"100101000",
13506=>"000111110",
13507=>"011110010",
13508=>"010000001",
13509=>"000011011",
13510=>"010000111",
13511=>"001001001",
13512=>"000000000",
13513=>"111111111",
13514=>"000010000",
13515=>"101100101",
13516=>"111101111",
13517=>"111000000",
13518=>"000000000",
13519=>"111101001",
13520=>"101001111",
13521=>"110010110",
13522=>"100101000",
13523=>"010110111",
13524=>"101100110",
13525=>"001000010",
13526=>"000010111",
13527=>"000010110",
13528=>"111101101",
13529=>"000101110",
13530=>"101001101",
13531=>"001101101",
13532=>"010000100",
13533=>"000111001",
13534=>"111111000",
13535=>"111000100",
13536=>"100100101",
13537=>"100110101",
13538=>"111111101",
13539=>"011010011",
13540=>"101101101",
13541=>"011010110",
13542=>"111111010",
13543=>"100110110",
13544=>"101111101",
13545=>"100000011",
13546=>"100100100",
13547=>"101111110",
13548=>"100000100",
13549=>"101001100",
13550=>"111000000",
13551=>"000000111",
13552=>"000001010",
13553=>"001001010",
13554=>"010000000",
13555=>"110010010",
13556=>"011011010",
13557=>"000010100",
13558=>"101100001",
13559=>"100110110",
13560=>"101001101",
13561=>"000000101",
13562=>"111101100",
13563=>"111111110",
13564=>"111110111",
13565=>"000111011",
13566=>"110110111",
13567=>"101001000",
13568=>"001000000",
13569=>"011001011",
13570=>"100100100",
13571=>"011010001",
13572=>"110000101",
13573=>"011110110",
13574=>"101111001",
13575=>"011011000",
13576=>"011000111",
13577=>"100100100",
13578=>"000011101",
13579=>"000011000",
13580=>"011011011",
13581=>"001001011",
13582=>"100110101",
13583=>"110010100",
13584=>"101000111",
13585=>"110100110",
13586=>"110110001",
13587=>"111100110",
13588=>"110100111",
13589=>"111100110",
13590=>"100111011",
13591=>"111111110",
13592=>"100100110",
13593=>"111010000",
13594=>"001001011",
13595=>"001001001",
13596=>"100110011",
13597=>"010000000",
13598=>"000100001",
13599=>"011001011",
13600=>"100110110",
13601=>"010001111",
13602=>"100001001",
13603=>"011011011",
13604=>"000000100",
13605=>"001011111",
13606=>"100100110",
13607=>"100000000",
13608=>"110110111",
13609=>"001001111",
13610=>"100110110",
13611=>"001011011",
13612=>"000000000",
13613=>"011100110",
13614=>"001111111",
13615=>"100110010",
13616=>"101100110",
13617=>"100100000",
13618=>"110100110",
13619=>"100110100",
13620=>"001000000",
13621=>"101011010",
13622=>"001011011",
13623=>"011000011",
13624=>"001100100",
13625=>"001000011",
13626=>"000000000",
13627=>"111100010",
13628=>"011011001",
13629=>"001011110",
13630=>"100100000",
13631=>"001000011",
13632=>"100110100",
13633=>"000100110",
13634=>"101111010",
13635=>"001010010",
13636=>"010101111",
13637=>"001001011",
13638=>"000010000",
13639=>"001111010",
13640=>"011111101",
13641=>"001000001",
13642=>"011010001",
13643=>"111011011",
13644=>"000100110",
13645=>"110110101",
13646=>"110110110",
13647=>"100110110",
13648=>"001000001",
13649=>"001100000",
13650=>"100101111",
13651=>"001100000",
13652=>"001111111",
13653=>"011001011",
13654=>"000001101",
13655=>"100000000",
13656=>"001011011",
13657=>"000110111",
13658=>"000000000",
13659=>"101110110",
13660=>"000010111",
13661=>"001001001",
13662=>"110100110",
13663=>"010000010",
13664=>"000001001",
13665=>"010001001",
13666=>"110110001",
13667=>"100011011",
13668=>"010000001",
13669=>"001001000",
13670=>"011001001",
13671=>"100100101",
13672=>"100001000",
13673=>"101110110",
13674=>"100110000",
13675=>"011000001",
13676=>"001001000",
13677=>"110111101",
13678=>"000001000",
13679=>"011011001",
13680=>"101010000",
13681=>"000001000",
13682=>"001001000",
13683=>"000000001",
13684=>"001011000",
13685=>"001110111",
13686=>"100001000",
13687=>"000000011",
13688=>"101101110",
13689=>"001001001",
13690=>"010110100",
13691=>"110110010",
13692=>"011010000",
13693=>"011010001",
13694=>"110110110",
13695=>"000010001",
13696=>"110100100",
13697=>"011001101",
13698=>"001111111",
13699=>"011110011",
13700=>"101000001",
13701=>"001111000",
13702=>"001101001",
13703=>"000011011",
13704=>"010011111",
13705=>"001111001",
13706=>"111011001",
13707=>"001100100",
13708=>"000010000",
13709=>"110110010",
13710=>"110110110",
13711=>"110000000",
13712=>"011011001",
13713=>"100000110",
13714=>"000010100",
13715=>"001010011",
13716=>"000000001",
13717=>"100100000",
13718=>"001001011",
13719=>"001100111",
13720=>"001001011",
13721=>"110000010",
13722=>"100110100",
13723=>"100110001",
13724=>"001010011",
13725=>"000110001",
13726=>"001110110",
13727=>"011010000",
13728=>"100001000",
13729=>"110111111",
13730=>"001001111",
13731=>"100110000",
13732=>"001110011",
13733=>"011000100",
13734=>"010010010",
13735=>"001001111",
13736=>"000100110",
13737=>"010100001",
13738=>"110110111",
13739=>"100000000",
13740=>"010100011",
13741=>"001010110",
13742=>"011010111",
13743=>"000101011",
13744=>"110101001",
13745=>"011001001",
13746=>"110110011",
13747=>"110001001",
13748=>"001000011",
13749=>"001011011",
13750=>"000000001",
13751=>"010111010",
13752=>"001000001",
13753=>"010000000",
13754=>"001001011",
13755=>"001011011",
13756=>"000001101",
13757=>"110111011",
13758=>"100110101",
13759=>"100100100",
13760=>"110110100",
13761=>"000110101",
13762=>"001111011",
13763=>"100110101",
13764=>"000100100",
13765=>"100101110",
13766=>"011001000",
13767=>"001001010",
13768=>"011000111",
13769=>"001001001",
13770=>"001010110",
13771=>"000000111",
13772=>"001110100",
13773=>"000011000",
13774=>"100000101",
13775=>"100000000",
13776=>"100100000",
13777=>"111011111",
13778=>"001000001",
13779=>"001001110",
13780=>"110110100",
13781=>"011011011",
13782=>"001001011",
13783=>"000110000",
13784=>"011001110",
13785=>"001001101",
13786=>"110001100",
13787=>"100110100",
13788=>"011011000",
13789=>"011001001",
13790=>"000000010",
13791=>"110100010",
13792=>"100100101",
13793=>"110110100",
13794=>"110100111",
13795=>"010001001",
13796=>"111000100",
13797=>"011011011",
13798=>"000000011",
13799=>"011010001",
13800=>"000000000",
13801=>"011000100",
13802=>"000000100",
13803=>"010101111",
13804=>"001001011",
13805=>"100001000",
13806=>"000100001",
13807=>"110010011",
13808=>"011001010",
13809=>"111111011",
13810=>"001101110",
13811=>"011001001",
13812=>"011010100",
13813=>"100100101",
13814=>"100100100",
13815=>"100110110",
13816=>"110100000",
13817=>"110110111",
13818=>"011011011",
13819=>"011011011",
13820=>"110100111",
13821=>"000110100",
13822=>"100010111",
13823=>"110110000",
13824=>"011011001",
13825=>"101101100",
13826=>"101000101",
13827=>"000000001",
13828=>"011000000",
13829=>"000100111",
13830=>"000000000",
13831=>"000100111",
13832=>"111100001",
13833=>"001010000",
13834=>"001000111",
13835=>"000000100",
13836=>"011000100",
13837=>"000111111",
13838=>"001011001",
13839=>"111011001",
13840=>"011101101",
13841=>"100001000",
13842=>"001000000",
13843=>"000000110",
13844=>"111111101",
13845=>"000000111",
13846=>"111001101",
13847=>"010110011",
13848=>"000111110",
13849=>"000001110",
13850=>"111111100",
13851=>"111000000",
13852=>"000000110",
13853=>"001111111",
13854=>"110100000",
13855=>"000111111",
13856=>"111100100",
13857=>"111011000",
13858=>"010010000",
13859=>"110111111",
13860=>"001011111",
13861=>"110000000",
13862=>"111010000",
13863=>"111000000",
13864=>"100100110",
13865=>"010100100",
13866=>"000111101",
13867=>"001001001",
13868=>"111011001",
13869=>"000001100",
13870=>"111011111",
13871=>"100000010",
13872=>"110111100",
13873=>"001100111",
13874=>"111111111",
13875=>"011001000",
13876=>"000000000",
13877=>"010001000",
13878=>"111111111",
13879=>"010111111",
13880=>"111111000",
13881=>"000000110",
13882=>"000110111",
13883=>"011001000",
13884=>"110111101",
13885=>"010111010",
13886=>"110111101",
13887=>"000010000",
13888=>"100001111",
13889=>"111101101",
13890=>"100101010",
13891=>"000000000",
13892=>"111011000",
13893=>"111110100",
13894=>"101000110",
13895=>"111000000",
13896=>"101011101",
13897=>"111111100",
13898=>"111001101",
13899=>"000011110",
13900=>"111111000",
13901=>"100001100",
13902=>"100000001",
13903=>"000000111",
13904=>"001000010",
13905=>"000111110",
13906=>"101010101",
13907=>"001001001",
13908=>"000000110",
13909=>"110110100",
13910=>"100110110",
13911=>"110010000",
13912=>"000101111",
13913=>"000111011",
13914=>"110010001",
13915=>"100110110",
13916=>"110010000",
13917=>"001001011",
13918=>"110110011",
13919=>"100000000",
13920=>"111110000",
13921=>"101110110",
13922=>"111110000",
13923=>"110100100",
13924=>"110111110",
13925=>"000011100",
13926=>"010010001",
13927=>"011000000",
13928=>"110000101",
13929=>"011000100",
13930=>"000000011",
13931=>"000110111",
13932=>"111111101",
13933=>"000100101",
13934=>"011101011",
13935=>"000000010",
13936=>"111111001",
13937=>"111111100",
13938=>"011111011",
13939=>"001111100",
13940=>"010000000",
13941=>"111000100",
13942=>"000000010",
13943=>"111010001",
13944=>"111100000",
13945=>"010100010",
13946=>"111011100",
13947=>"000100000",
13948=>"100110111",
13949=>"100100100",
13950=>"111101101",
13951=>"000111100",
13952=>"111100100",
13953=>"100011110",
13954=>"111110000",
13955=>"010000001",
13956=>"010000100",
13957=>"000010101",
13958=>"110101100",
13959=>"001001000",
13960=>"111111010",
13961=>"000000111",
13962=>"110110111",
13963=>"010010111",
13964=>"110000000",
13965=>"000101100",
13966=>"101111101",
13967=>"010000000",
13968=>"101000010",
13969=>"000000101",
13970=>"110111101",
13971=>"001000001",
13972=>"000111111",
13973=>"000000101",
13974=>"000111000",
13975=>"011011001",
13976=>"101111111",
13977=>"000000111",
13978=>"000100111",
13979=>"101101111",
13980=>"111111101",
13981=>"111000111",
13982=>"001101111",
13983=>"000010000",
13984=>"101010111",
13985=>"001000000",
13986=>"011001111",
13987=>"000111000",
13988=>"100000111",
13989=>"110111100",
13990=>"110110000",
13991=>"001101111",
13992=>"100011111",
13993=>"111111000",
13994=>"000000100",
13995=>"000000010",
13996=>"110010100",
13997=>"111000100",
13998=>"011001010",
13999=>"000000000",
14000=>"110001101",
14001=>"101000001",
14002=>"111011011",
14003=>"000100100",
14004=>"111111000",
14005=>"111111000",
14006=>"111111111",
14007=>"111001000",
14008=>"011111011",
14009=>"000110110",
14010=>"000101010",
14011=>"011111000",
14012=>"000100111",
14013=>"111111110",
14014=>"101100010",
14015=>"000000000",
14016=>"011011001",
14017=>"010010000",
14018=>"101111010",
14019=>"100100110",
14020=>"000000000",
14021=>"100110001",
14022=>"111111111",
14023=>"000000000",
14024=>"101101111",
14025=>"111000000",
14026=>"111111111",
14027=>"000001111",
14028=>"000000111",
14029=>"001111110",
14030=>"011011010",
14031=>"000001111",
14032=>"000000000",
14033=>"100111111",
14034=>"000000100",
14035=>"000101101",
14036=>"011010001",
14037=>"110111111",
14038=>"101111000",
14039=>"000001011",
14040=>"000010111",
14041=>"010110000",
14042=>"000110101",
14043=>"010010000",
14044=>"111001001",
14045=>"011000110",
14046=>"011010000",
14047=>"001000000",
14048=>"000101111",
14049=>"101100100",
14050=>"100000111",
14051=>"110100101",
14052=>"000010000",
14053=>"111010000",
14054=>"000010111",
14055=>"101110110",
14056=>"010101111",
14057=>"111010100",
14058=>"100001111",
14059=>"111101000",
14060=>"000000000",
14061=>"111000111",
14062=>"010010000",
14063=>"101101110",
14064=>"000111111",
14065=>"011111111",
14066=>"111000000",
14067=>"100100100",
14068=>"110110000",
14069=>"010000111",
14070=>"001000000",
14071=>"000100001",
14072=>"000111111",
14073=>"000001010",
14074=>"010000011",
14075=>"100101110",
14076=>"000111111",
14077=>"011011000",
14078=>"111111110",
14079=>"000001011",
14080=>"001111111",
14081=>"100111010",
14082=>"000100100",
14083=>"111101000",
14084=>"001101011",
14085=>"000001111",
14086=>"101101011",
14087=>"101111110",
14088=>"111010000",
14089=>"011010000",
14090=>"001000000",
14091=>"000000000",
14092=>"101100100",
14093=>"011110000",
14094=>"011001000",
14095=>"000111111",
14096=>"010000000",
14097=>"010000000",
14098=>"000100011",
14099=>"100000000",
14100=>"100011010",
14101=>"011000110",
14102=>"100100001",
14103=>"001111111",
14104=>"101100000",
14105=>"110001111",
14106=>"000011000",
14107=>"000100010",
14108=>"000000010",
14109=>"000000101",
14110=>"011011111",
14111=>"111111001",
14112=>"110100110",
14113=>"011111011",
14114=>"100000000",
14115=>"110010000",
14116=>"001011001",
14117=>"101011111",
14118=>"011010110",
14119=>"101001010",
14120=>"000111111",
14121=>"010111000",
14122=>"000000000",
14123=>"100100111",
14124=>"001001111",
14125=>"101111001",
14126=>"000101111",
14127=>"100101101",
14128=>"101011010",
14129=>"000001000",
14130=>"010010000",
14131=>"011001101",
14132=>"000000000",
14133=>"010011111",
14134=>"110011010",
14135=>"111101000",
14136=>"110111111",
14137=>"000000000",
14138=>"111100000",
14139=>"001000000",
14140=>"010011110",
14141=>"111111111",
14142=>"010000000",
14143=>"111011000",
14144=>"101000100",
14145=>"000100101",
14146=>"111111000",
14147=>"011000000",
14148=>"100111111",
14149=>"000000011",
14150=>"010010000",
14151=>"111101101",
14152=>"000001001",
14153=>"011010000",
14154=>"000000000",
14155=>"100010111",
14156=>"010000000",
14157=>"101101000",
14158=>"000110110",
14159=>"000011000",
14160=>"001000000",
14161=>"101110001",
14162=>"110111111",
14163=>"000100001",
14164=>"000000000",
14165=>"100100011",
14166=>"101100100",
14167=>"111000000",
14168=>"010000000",
14169=>"111011011",
14170=>"100111011",
14171=>"110100001",
14172=>"111000001",
14173=>"001001011",
14174=>"100010010",
14175=>"101001100",
14176=>"011010000",
14177=>"000000110",
14178=>"111000000",
14179=>"000000110",
14180=>"010010000",
14181=>"001001000",
14182=>"100111011",
14183=>"111101000",
14184=>"101011011",
14185=>"010000110",
14186=>"001111111",
14187=>"111000001",
14188=>"000001100",
14189=>"000010010",
14190=>"111000000",
14191=>"011000111",
14192=>"001011000",
14193=>"010110111",
14194=>"111111011",
14195=>"000000000",
14196=>"001001010",
14197=>"000010000",
14198=>"111010010",
14199=>"111000000",
14200=>"000010111",
14201=>"111100000",
14202=>"100101111",
14203=>"000000101",
14204=>"110010000",
14205=>"100001110",
14206=>"000000010",
14207=>"000000000",
14208=>"110010000",
14209=>"000000111",
14210=>"111000100",
14211=>"110110010",
14212=>"111111110",
14213=>"111000010",
14214=>"111110111",
14215=>"000000100",
14216=>"101111000",
14217=>"000000000",
14218=>"100011011",
14219=>"111001011",
14220=>"111000011",
14221=>"000100111",
14222=>"111111010",
14223=>"000001000",
14224=>"100100101",
14225=>"000001101",
14226=>"001010000",
14227=>"000000101",
14228=>"101011011",
14229=>"011000000",
14230=>"111010010",
14231=>"110011000",
14232=>"000010000",
14233=>"101111011",
14234=>"000000100",
14235=>"000000101",
14236=>"011111000",
14237=>"111011000",
14238=>"011111111",
14239=>"000001111",
14240=>"000101101",
14241=>"100110111",
14242=>"111010011",
14243=>"000011101",
14244=>"111011111",
14245=>"000000000",
14246=>"000010100",
14247=>"100001011",
14248=>"110010010",
14249=>"011011000",
14250=>"000000111",
14251=>"000000111",
14252=>"111010001",
14253=>"011000000",
14254=>"101111100",
14255=>"010000000",
14256=>"001010010",
14257=>"110110000",
14258=>"000100000",
14259=>"110110000",
14260=>"010000011",
14261=>"101001111",
14262=>"000100100",
14263=>"000111111",
14264=>"000100011",
14265=>"101111000",
14266=>"111011011",
14267=>"011010000",
14268=>"010111111",
14269=>"111111100",
14270=>"111000000",
14271=>"000000100",
14272=>"000100100",
14273=>"111100000",
14274=>"011111000",
14275=>"000000000",
14276=>"100110010",
14277=>"001100100",
14278=>"101011010",
14279=>"000000010",
14280=>"000010010",
14281=>"100100101",
14282=>"111101110",
14283=>"111111011",
14284=>"001011001",
14285=>"011011000",
14286=>"100000011",
14287=>"111101100",
14288=>"010011000",
14289=>"110110001",
14290=>"011001000",
14291=>"111110111",
14292=>"000000000",
14293=>"100110011",
14294=>"010010010",
14295=>"001000000",
14296=>"000010011",
14297=>"000000111",
14298=>"100101000",
14299=>"000000101",
14300=>"001101111",
14301=>"101011010",
14302=>"000100101",
14303=>"010100010",
14304=>"001000100",
14305=>"000101000",
14306=>"000000010",
14307=>"111010000",
14308=>"010000000",
14309=>"101111111",
14310=>"111000111",
14311=>"100110010",
14312=>"111111011",
14313=>"010011111",
14314=>"000000000",
14315=>"000100111",
14316=>"111001000",
14317=>"010101111",
14318=>"110000110",
14319=>"000000000",
14320=>"000011011",
14321=>"100100101",
14322=>"010100000",
14323=>"011100110",
14324=>"101001111",
14325=>"001100010",
14326=>"100100000",
14327=>"000000000",
14328=>"101101100",
14329=>"111011010",
14330=>"110100111",
14331=>"110100101",
14332=>"011011000",
14333=>"100011111",
14334=>"101111100",
14335=>"010010000",
14336=>"000000100",
14337=>"101101111",
14338=>"111100000",
14339=>"000111010",
14340=>"000110111",
14341=>"110110101",
14342=>"000000111",
14343=>"011010111",
14344=>"000000010",
14345=>"010000000",
14346=>"111101000",
14347=>"001101000",
14348=>"000000000",
14349=>"001001000",
14350=>"000100101",
14351=>"111111111",
14352=>"111000000",
14353=>"111000011",
14354=>"111111111",
14355=>"000000000",
14356=>"101000001",
14357=>"100100111",
14358=>"000000100",
14359=>"110000110",
14360=>"100101000",
14361=>"001111111",
14362=>"100100110",
14363=>"111000000",
14364=>"101001011",
14365=>"000101010",
14366=>"001000100",
14367=>"000000000",
14368=>"111111000",
14369=>"101010010",
14370=>"010110010",
14371=>"010000100",
14372=>"000001111",
14373=>"100000001",
14374=>"110001100",
14375=>"111111110",
14376=>"111111010",
14377=>"100100000",
14378=>"001000000",
14379=>"111111000",
14380=>"011011011",
14381=>"010010000",
14382=>"011010111",
14383=>"000111010",
14384=>"000110110",
14385=>"010001111",
14386=>"111111101",
14387=>"010000000",
14388=>"001001000",
14389=>"000111000",
14390=>"000000000",
14391=>"000101111",
14392=>"001111111",
14393=>"101000100",
14394=>"111001111",
14395=>"111111111",
14396=>"001000111",
14397=>"111000010",
14398=>"000000100",
14399=>"110111111",
14400=>"000000011",
14401=>"001101001",
14402=>"111111110",
14403=>"111110110",
14404=>"110000000",
14405=>"100000000",
14406=>"000011111",
14407=>"111111010",
14408=>"000000001",
14409=>"111111100",
14410=>"111000000",
14411=>"000010111",
14412=>"111111101",
14413=>"110100101",
14414=>"000000110",
14415=>"000110110",
14416=>"101101101",
14417=>"110010000",
14418=>"000000100",
14419=>"000011001",
14420=>"101101101",
14421=>"000010100",
14422=>"011000100",
14423=>"110111011",
14424=>"010000001",
14425=>"110100111",
14426=>"100110100",
14427=>"011111111",
14428=>"100000111",
14429=>"000100000",
14430=>"100010111",
14431=>"010010011",
14432=>"111111111",
14433=>"101101110",
14434=>"111000000",
14435=>"001011011",
14436=>"000000000",
14437=>"001011111",
14438=>"100111110",
14439=>"101001000",
14440=>"000111111",
14441=>"000000010",
14442=>"111100100",
14443=>"001101000",
14444=>"101001101",
14445=>"110010010",
14446=>"000000011",
14447=>"110101111",
14448=>"011101111",
14449=>"000010100",
14450=>"111000000",
14451=>"110000000",
14452=>"011110100",
14453=>"111101101",
14454=>"111000000",
14455=>"010111111",
14456=>"101101110",
14457=>"011011000",
14458=>"111111111",
14459=>"010010111",
14460=>"000000100",
14461=>"000110000",
14462=>"101010000",
14463=>"101101001",
14464=>"011110101",
14465=>"011011000",
14466=>"101001010",
14467=>"000101001",
14468=>"101000110",
14469=>"000110011",
14470=>"101001111",
14471=>"011001001",
14472=>"100100110",
14473=>"111111110",
14474=>"010010010",
14475=>"111111011",
14476=>"000000111",
14477=>"111111100",
14478=>"011010000",
14479=>"111100000",
14480=>"001100111",
14481=>"000000110",
14482=>"000000000",
14483=>"000000000",
14484=>"010000001",
14485=>"111001000",
14486=>"011011111",
14487=>"000100111",
14488=>"111111010",
14489=>"110001000",
14490=>"000101001",
14491=>"000010000",
14492=>"100101101",
14493=>"010000000",
14494=>"000101111",
14495=>"110000000",
14496=>"001011011",
14497=>"010011111",
14498=>"000000100",
14499=>"111000000",
14500=>"111000111",
14501=>"010111110",
14502=>"101000000",
14503=>"010000110",
14504=>"111000000",
14505=>"000010001",
14506=>"111111001",
14507=>"111000000",
14508=>"000000000",
14509=>"010000000",
14510=>"000101011",
14511=>"010010000",
14512=>"111110110",
14513=>"101000111",
14514=>"000000010",
14515=>"010001000",
14516=>"100011100",
14517=>"000000000",
14518=>"000111111",
14519=>"000111111",
14520=>"101000101",
14521=>"010001110",
14522=>"000101000",
14523=>"001101101",
14524=>"000100010",
14525=>"010110100",
14526=>"001011000",
14527=>"111111111",
14528=>"001100001",
14529=>"111000111",
14530=>"111111001",
14531=>"110010001",
14532=>"010111011",
14533=>"000110100",
14534=>"000000000",
14535=>"111011010",
14536=>"000001010",
14537=>"000000000",
14538=>"000111111",
14539=>"101000100",
14540=>"000100110",
14541=>"100100000",
14542=>"101101101",
14543=>"000000011",
14544=>"101101111",
14545=>"000111111",
14546=>"101101000",
14547=>"010011111",
14548=>"101011111",
14549=>"101001011",
14550=>"111101101",
14551=>"000110111",
14552=>"000000000",
14553=>"100000010",
14554=>"000110110",
14555=>"101101101",
14556=>"111101011",
14557=>"111111111",
14558=>"110111101",
14559=>"111000100",
14560=>"001000010",
14561=>"111011011",
14562=>"101010010",
14563=>"000011111",
14564=>"111000111",
14565=>"000111111",
14566=>"010001001",
14567=>"001001111",
14568=>"111011010",
14569=>"101100111",
14570=>"111100000",
14571=>"000110110",
14572=>"000000000",
14573=>"001111111",
14574=>"110000000",
14575=>"000010000",
14576=>"111000111",
14577=>"010001001",
14578=>"111000100",
14579=>"000111011",
14580=>"000000110",
14581=>"101101101",
14582=>"010010000",
14583=>"101010000",
14584=>"000000111",
14585=>"011111111",
14586=>"000011000",
14587=>"101110001",
14588=>"000110111",
14589=>"000000011",
14590=>"001011110",
14591=>"111111111",
14592=>"000000000",
14593=>"000010010",
14594=>"111000000",
14595=>"101101010",
14596=>"111111101",
14597=>"110000111",
14598=>"000111110",
14599=>"110111111",
14600=>"010010010",
14601=>"101010010",
14602=>"100110111",
14603=>"100000000",
14604=>"000000011",
14605=>"101111001",
14606=>"110011011",
14607=>"000010101",
14608=>"000110110",
14609=>"000010011",
14610=>"010000000",
14611=>"000010111",
14612=>"111011010",
14613=>"101111111",
14614=>"010111100",
14615=>"011011011",
14616=>"111000100",
14617=>"000010000",
14618=>"010001001",
14619=>"000000000",
14620=>"000001001",
14621=>"000010100",
14622=>"111011001",
14623=>"000000101",
14624=>"000100001",
14625=>"011110111",
14626=>"111101111",
14627=>"000111111",
14628=>"011100000",
14629=>"101100001",
14630=>"001101001",
14631=>"000010010",
14632=>"101011010",
14633=>"001111111",
14634=>"100010011",
14635=>"000000100",
14636=>"000101111",
14637=>"111111010",
14638=>"000111111",
14639=>"010001101",
14640=>"111111001",
14641=>"111111100",
14642=>"010001001",
14643=>"111111010",
14644=>"000000000",
14645=>"000000110",
14646=>"001000000",
14647=>"000000000",
14648=>"000011011",
14649=>"000001001",
14650=>"011000101",
14651=>"011011010",
14652=>"010110010",
14653=>"011001000",
14654=>"000100000",
14655=>"110010110",
14656=>"111010111",
14657=>"100100111",
14658=>"111011111",
14659=>"100100011",
14660=>"111000111",
14661=>"000011011",
14662=>"011011111",
14663=>"000000000",
14664=>"110101101",
14665=>"000111111",
14666=>"000000000",
14667=>"101000010",
14668=>"101000011",
14669=>"000001010",
14670=>"011001101",
14671=>"111111111",
14672=>"001000111",
14673=>"101111000",
14674=>"111111100",
14675=>"001001100",
14676=>"101000000",
14677=>"000000000",
14678=>"100111101",
14679=>"100010010",
14680=>"111000001",
14681=>"110101100",
14682=>"111100111",
14683=>"000011110",
14684=>"000010111",
14685=>"000001001",
14686=>"100010010",
14687=>"001011111",
14688=>"111010111",
14689=>"000110111",
14690=>"111000111",
14691=>"110100101",
14692=>"000101111",
14693=>"000011111",
14694=>"000010001",
14695=>"000010011",
14696=>"000100111",
14697=>"111010000",
14698=>"000110000",
14699=>"000101000",
14700=>"110111000",
14701=>"000110111",
14702=>"000110011",
14703=>"101111100",
14704=>"010111111",
14705=>"100011101",
14706=>"000000010",
14707=>"000000000",
14708=>"111101000",
14709=>"011000101",
14710=>"000000010",
14711=>"000110111",
14712=>"111000100",
14713=>"000111100",
14714=>"110000011",
14715=>"000011010",
14716=>"010100010",
14717=>"100100000",
14718=>"001101111",
14719=>"111101111",
14720=>"100100111",
14721=>"010000000",
14722=>"001111010",
14723=>"000101101",
14724=>"000111000",
14725=>"111101101",
14726=>"001011110",
14727=>"100000010",
14728=>"100111011",
14729=>"101011000",
14730=>"000011001",
14731=>"010110011",
14732=>"100000110",
14733=>"000000111",
14734=>"000111111",
14735=>"001100111",
14736=>"011001101",
14737=>"010000111",
14738=>"111000000",
14739=>"000010010",
14740=>"000100111",
14741=>"000010010",
14742=>"111111000",
14743=>"100101101",
14744=>"100100111",
14745=>"010000101",
14746=>"111101101",
14747=>"110101100",
14748=>"000000000",
14749=>"101000000",
14750=>"001110000",
14751=>"000010000",
14752=>"100101000",
14753=>"010010000",
14754=>"000111010",
14755=>"111010101",
14756=>"000110100",
14757=>"000000011",
14758=>"000111011",
14759=>"000101111",
14760=>"100011110",
14761=>"101000010",
14762=>"111101101",
14763=>"000000100",
14764=>"111010011",
14765=>"100011011",
14766=>"111101111",
14767=>"101010110",
14768=>"111000000",
14769=>"011001111",
14770=>"000001111",
14771=>"011001000",
14772=>"000100111",
14773=>"111101001",
14774=>"111100101",
14775=>"000011011",
14776=>"000011000",
14777=>"001011001",
14778=>"000101000",
14779=>"011111010",
14780=>"001000101",
14781=>"111000000",
14782=>"011000011",
14783=>"000110101",
14784=>"000010000",
14785=>"000110111",
14786=>"101101011",
14787=>"000001100",
14788=>"111000111",
14789=>"110110000",
14790=>"011110000",
14791=>"000111111",
14792=>"100010011",
14793=>"000000101",
14794=>"000000001",
14795=>"100101000",
14796=>"000000001",
14797=>"000010010",
14798=>"010000110",
14799=>"111010001",
14800=>"010000000",
14801=>"000001001",
14802=>"100000000",
14803=>"010010010",
14804=>"110111110",
14805=>"000000110",
14806=>"011010000",
14807=>"101111011",
14808=>"001101111",
14809=>"000000101",
14810=>"011001101",
14811=>"111000010",
14812=>"010110000",
14813=>"000010111",
14814=>"011011111",
14815=>"101111001",
14816=>"101000111",
14817=>"111011010",
14818=>"111000111",
14819=>"011111110",
14820=>"000000010",
14821=>"111001000",
14822=>"111111001",
14823=>"100011111",
14824=>"001100110",
14825=>"110110000",
14826=>"001111111",
14827=>"010011111",
14828=>"101000000",
14829=>"111100111",
14830=>"001000000",
14831=>"000100100",
14832=>"011111010",
14833=>"011011001",
14834=>"111111111",
14835=>"000001101",
14836=>"000100100",
14837=>"111101101",
14838=>"101000010",
14839=>"111000000",
14840=>"100000010",
14841=>"010110011",
14842=>"000000100",
14843=>"000000000",
14844=>"111101001",
14845=>"010111000",
14846=>"000100111",
14847=>"110111110",
14848=>"000001000",
14849=>"000000100",
14850=>"111000000",
14851=>"111111111",
14852=>"000000011",
14853=>"000001110",
14854=>"111000101",
14855=>"000101111",
14856=>"101111111",
14857=>"101101111",
14858=>"000000000",
14859=>"011000001",
14860=>"111011000",
14861=>"011011000",
14862=>"011101001",
14863=>"000111111",
14864=>"001011000",
14865=>"000000000",
14866=>"100000000",
14867=>"000000001",
14868=>"101000111",
14869=>"101100000",
14870=>"001111111",
14871=>"100100111",
14872=>"000000000",
14873=>"000010000",
14874=>"000000000",
14875=>"001000000",
14876=>"000000100",
14877=>"000000000",
14878=>"110111001",
14879=>"000111001",
14880=>"111111111",
14881=>"101111011",
14882=>"001111001",
14883=>"111111111",
14884=>"000000000",
14885=>"001101111",
14886=>"111100000",
14887=>"100110010",
14888=>"000111111",
14889=>"101111001",
14890=>"000000000",
14891=>"011111111",
14892=>"001011001",
14893=>"101111000",
14894=>"101111111",
14895=>"000000100",
14896=>"000000000",
14897=>"110110010",
14898=>"001111111",
14899=>"000110000",
14900=>"000000000",
14901=>"000000000",
14902=>"001000000",
14903=>"000110100",
14904=>"111111111",
14905=>"000000000",
14906=>"000000000",
14907=>"000100111",
14908=>"111011111",
14909=>"111111001",
14910=>"000000100",
14911=>"111111110",
14912=>"000000001",
14913=>"000111101",
14914=>"000101011",
14915=>"010110011",
14916=>"111111000",
14917=>"000000000",
14918=>"101101000",
14919=>"111111111",
14920=>"010111101",
14921=>"111111110",
14922=>"000000000",
14923=>"000000000",
14924=>"111100001",
14925=>"000010000",
14926=>"011100101",
14927=>"111111111",
14928=>"000000000",
14929=>"111111110",
14930=>"101111111",
14931=>"111011000",
14932=>"111001110",
14933=>"010100110",
14934=>"001100000",
14935=>"100010000",
14936=>"010000010",
14937=>"011001001",
14938=>"100110000",
14939=>"110010010",
14940=>"111000000",
14941=>"001011111",
14942=>"111111111",
14943=>"011001000",
14944=>"010101100",
14945=>"111110011",
14946=>"110000000",
14947=>"000100000",
14948=>"100000000",
14949=>"000000000",
14950=>"111111111",
14951=>"100100000",
14952=>"100101111",
14953=>"000000000",
14954=>"000100111",
14955=>"111111111",
14956=>"111010111",
14957=>"000000000",
14958=>"000010010",
14959=>"000000110",
14960=>"001011001",
14961=>"000000111",
14962=>"001001000",
14963=>"000000000",
14964=>"111110000",
14965=>"000000100",
14966=>"110000000",
14967=>"101111101",
14968=>"101000111",
14969=>"111011111",
14970=>"000111010",
14971=>"111111111",
14972=>"110110000",
14973=>"110111001",
14974=>"101101110",
14975=>"110000111",
14976=>"000111000",
14977=>"111111010",
14978=>"111111111",
14979=>"011111111",
14980=>"010000000",
14981=>"001000000",
14982=>"000110101",
14983=>"001011001",
14984=>"101101100",
14985=>"000000000",
14986=>"000000000",
14987=>"101101000",
14988=>"001000101",
14989=>"001111111",
14990=>"100000000",
14991=>"000000000",
14992=>"000001001",
14993=>"111111111",
14994=>"000000000",
14995=>"001111111",
14996=>"001001100",
14997=>"000110000",
14998=>"000001001",
14999=>"100101101",
15000=>"101111111",
15001=>"001001111",
15002=>"010011000",
15003=>"110100101",
15004=>"111011000",
15005=>"011000000",
15006=>"111101111",
15007=>"001010111",
15008=>"011011011",
15009=>"000000110",
15010=>"000101111",
15011=>"101100101",
15012=>"100110000",
15013=>"110110000",
15014=>"001100000",
15015=>"000011111",
15016=>"000000111",
15017=>"101100101",
15018=>"000010010",
15019=>"000000000",
15020=>"111111011",
15021=>"111101100",
15022=>"111011111",
15023=>"111111010",
15024=>"111111111",
15025=>"000010000",
15026=>"110101111",
15027=>"110100110",
15028=>"100110000",
15029=>"111111111",
15030=>"100001101",
15031=>"000011111",
15032=>"111100111",
15033=>"100100000",
15034=>"110011000",
15035=>"111111111",
15036=>"000010001",
15037=>"111111111",
15038=>"111111111",
15039=>"011100000",
15040=>"011000100",
15041=>"000001001",
15042=>"101111011",
15043=>"000101001",
15044=>"000000000",
15045=>"100101110",
15046=>"000011111",
15047=>"001000110",
15048=>"100111101",
15049=>"000000100",
15050=>"110001101",
15051=>"000000000",
15052=>"101100101",
15053=>"111001001",
15054=>"000000000",
15055=>"111111000",
15056=>"111001000",
15057=>"011111001",
15058=>"001000010",
15059=>"000000001",
15060=>"111110111",
15061=>"000000101",
15062=>"111111010",
15063=>"000000001",
15064=>"001111101",
15065=>"111111111",
15066=>"110110101",
15067=>"000000000",
15068=>"000001010",
15069=>"111110111",
15070=>"000000000",
15071=>"001101111",
15072=>"111101001",
15073=>"000000000",
15074=>"111111110",
15075=>"000110010",
15076=>"000000000",
15077=>"011001001",
15078=>"011011101",
15079=>"111111111",
15080=>"110101111",
15081=>"100101111",
15082=>"000000000",
15083=>"100000010",
15084=>"110001010",
15085=>"000000000",
15086=>"111111110",
15087=>"111111001",
15088=>"000110110",
15089=>"001011111",
15090=>"111111111",
15091=>"111111001",
15092=>"001011011",
15093=>"000000000",
15094=>"000011111",
15095=>"000011011",
15096=>"010111111",
15097=>"001111111",
15098=>"111111111",
15099=>"000011000",
15100=>"000001001",
15101=>"111111111",
15102=>"000001101",
15103=>"000010000",
15104=>"001100100",
15105=>"111001000",
15106=>"111101111",
15107=>"010111111",
15108=>"011111000",
15109=>"110101111",
15110=>"000000000",
15111=>"110110111",
15112=>"100000101",
15113=>"100111111",
15114=>"111011100",
15115=>"111111000",
15116=>"111000101",
15117=>"001000000",
15118=>"111100000",
15119=>"000001100",
15120=>"010000001",
15121=>"101000000",
15122=>"110111001",
15123=>"000000010",
15124=>"111000100",
15125=>"111001101",
15126=>"111111011",
15127=>"000010111",
15128=>"001110000",
15129=>"000111111",
15130=>"000000010",
15131=>"000111000",
15132=>"111100101",
15133=>"000000010",
15134=>"100000010",
15135=>"111101101",
15136=>"111110000",
15137=>"011010111",
15138=>"010111100",
15139=>"111111111",
15140=>"010011111",
15141=>"000111101",
15142=>"111000000",
15143=>"010101000",
15144=>"010111111",
15145=>"111000100",
15146=>"010001001",
15147=>"010111111",
15148=>"011011011",
15149=>"000001011",
15150=>"010000010",
15151=>"000110101",
15152=>"000011011",
15153=>"111111111",
15154=>"000000100",
15155=>"001010111",
15156=>"000000000",
15157=>"111111111",
15158=>"111011001",
15159=>"101000000",
15160=>"000000010",
15161=>"111001000",
15162=>"100000000",
15163=>"000111111",
15164=>"111101001",
15165=>"111111111",
15166=>"100000000",
15167=>"111110111",
15168=>"000111111",
15169=>"000001110",
15170=>"000000111",
15171=>"000000000",
15172=>"100010010",
15173=>"000101111",
15174=>"000011010",
15175=>"111101111",
15176=>"000100010",
15177=>"000000000",
15178=>"110111111",
15179=>"111001111",
15180=>"000001000",
15181=>"000111011",
15182=>"111111111",
15183=>"010101000",
15184=>"000100101",
15185=>"111110101",
15186=>"000000101",
15187=>"101110010",
15188=>"000000111",
15189=>"111001001",
15190=>"111110110",
15191=>"010000000",
15192=>"000000001",
15193=>"111001000",
15194=>"000000000",
15195=>"101011000",
15196=>"111101101",
15197=>"111010100",
15198=>"000111111",
15199=>"100000000",
15200=>"111000000",
15201=>"000111111",
15202=>"000011011",
15203=>"100000000",
15204=>"011101001",
15205=>"000100100",
15206=>"101000000",
15207=>"111100000",
15208=>"111111111",
15209=>"001011111",
15210=>"010111111",
15211=>"111000100",
15212=>"101110110",
15213=>"001111111",
15214=>"101000000",
15215=>"000000000",
15216=>"000001101",
15217=>"100000000",
15218=>"100110000",
15219=>"111000000",
15220=>"000000000",
15221=>"101100111",
15222=>"111000000",
15223=>"101000000",
15224=>"111101001",
15225=>"111111111",
15226=>"111001000",
15227=>"000111111",
15228=>"000000010",
15229=>"111011010",
15230=>"110100111",
15231=>"000011111",
15232=>"000011111",
15233=>"000000111",
15234=>"000001000",
15235=>"011111111",
15236=>"001001000",
15237=>"110001010",
15238=>"000100110",
15239=>"001010000",
15240=>"100110011",
15241=>"000111111",
15242=>"110111000",
15243=>"011100110",
15244=>"111000000",
15245=>"000101101",
15246=>"000111111",
15247=>"000000000",
15248=>"001011000",
15249=>"010000001",
15250=>"111101000",
15251=>"111101011",
15252=>"000100000",
15253=>"111000000",
15254=>"000010000",
15255=>"100000000",
15256=>"001000000",
15257=>"000010111",
15258=>"010111111",
15259=>"000111000",
15260=>"111100000",
15261=>"000111111",
15262=>"000101111",
15263=>"111000000",
15264=>"011111100",
15265=>"011010000",
15266=>"010000000",
15267=>"000000100",
15268=>"101000000",
15269=>"011011000",
15270=>"110100101",
15271=>"000010000",
15272=>"000110000",
15273=>"010111000",
15274=>"000000000",
15275=>"100000000",
15276=>"011001001",
15277=>"000011111",
15278=>"000000010",
15279=>"000111111",
15280=>"000000111",
15281=>"001100000",
15282=>"001111111",
15283=>"110111001",
15284=>"111011000",
15285=>"010000000",
15286=>"011101000",
15287=>"101100000",
15288=>"111001000",
15289=>"101011001",
15290=>"010000000",
15291=>"010100000",
15292=>"111101000",
15293=>"000111111",
15294=>"110111011",
15295=>"000000000",
15296=>"000010111",
15297=>"000000111",
15298=>"010111000",
15299=>"100000000",
15300=>"111111000",
15301=>"001001001",
15302=>"000000001",
15303=>"100100111",
15304=>"001000101",
15305=>"001101111",
15306=>"111101001",
15307=>"100000000",
15308=>"010000000",
15309=>"000010000",
15310=>"111100000",
15311=>"100011010",
15312=>"111011010",
15313=>"010111110",
15314=>"000001000",
15315=>"010111110",
15316=>"001000110",
15317=>"101000000",
15318=>"011000000",
15319=>"010001111",
15320=>"111100101",
15321=>"111111000",
15322=>"100111001",
15323=>"000111111",
15324=>"111111100",
15325=>"010011001",
15326=>"001000000",
15327=>"111111111",
15328=>"011111111",
15329=>"000000011",
15330=>"000000000",
15331=>"100011111",
15332=>"101000000",
15333=>"000111111",
15334=>"111111101",
15335=>"001000010",
15336=>"111111001",
15337=>"110111110",
15338=>"011100000",
15339=>"000000000",
15340=>"111000000",
15341=>"101101111",
15342=>"110000010",
15343=>"001000000",
15344=>"111010000",
15345=>"110100000",
15346=>"000000100",
15347=>"111111000",
15348=>"101011011",
15349=>"000000000",
15350=>"000101010",
15351=>"110100000",
15352=>"011000000",
15353=>"000010111",
15354=>"110100000",
15355=>"010111000",
15356=>"100000000",
15357=>"010111111",
15358=>"110110110",
15359=>"110101001",
15360=>"000000111",
15361=>"000000001",
15362=>"111111000",
15363=>"111010000",
15364=>"000000110",
15365=>"000001111",
15366=>"000111111",
15367=>"000000000",
15368=>"000000000",
15369=>"111111000",
15370=>"001011011",
15371=>"011001000",
15372=>"011001101",
15373=>"000000000",
15374=>"010010100",
15375=>"000000000",
15376=>"110000111",
15377=>"111000010",
15378=>"111110110",
15379=>"000001011",
15380=>"111101100",
15381=>"001000101",
15382=>"000110010",
15383=>"001000101",
15384=>"000001001",
15385=>"110111101",
15386=>"000000000",
15387=>"111110000",
15388=>"011011101",
15389=>"000000000",
15390=>"111001010",
15391=>"110100111",
15392=>"111110010",
15393=>"010100000",
15394=>"000001001",
15395=>"011111001",
15396=>"010000011",
15397=>"000000000",
15398=>"100100101",
15399=>"111001001",
15400=>"111111111",
15401=>"000000100",
15402=>"000000111",
15403=>"011111001",
15404=>"010111011",
15405=>"000000000",
15406=>"011111111",
15407=>"011000000",
15408=>"000000110",
15409=>"011000110",
15410=>"000000000",
15411=>"000111111",
15412=>"101100111",
15413=>"101101001",
15414=>"000011001",
15415=>"000111111",
15416=>"000000000",
15417=>"000000111",
15418=>"001001000",
15419=>"000000000",
15420=>"000000000",
15421=>"111111111",
15422=>"001001101",
15423=>"100100110",
15424=>"000000010",
15425=>"111001000",
15426=>"010110010",
15427=>"000100110",
15428=>"000000000",
15429=>"000000000",
15430=>"010111111",
15431=>"001001111",
15432=>"000000010",
15433=>"111000111",
15434=>"001101101",
15435=>"111000011",
15436=>"010111111",
15437=>"111011010",
15438=>"000010110",
15439=>"000111110",
15440=>"110110110",
15441=>"111111000",
15442=>"001001111",
15443=>"010110011",
15444=>"110101101",
15445=>"011000000",
15446=>"111010010",
15447=>"111111000",
15448=>"000110111",
15449=>"000010111",
15450=>"011111111",
15451=>"111111110",
15452=>"111110010",
15453=>"001011001",
15454=>"110100111",
15455=>"000111010",
15456=>"010011000",
15457=>"010010000",
15458=>"011001101",
15459=>"110111110",
15460=>"000000110",
15461=>"011010000",
15462=>"101100110",
15463=>"111111000",
15464=>"000001111",
15465=>"000000001",
15466=>"000000000",
15467=>"000001111",
15468=>"000001000",
15469=>"000000010",
15470=>"011000000",
15471=>"010000000",
15472=>"010110110",
15473=>"000001000",
15474=>"000000110",
15475=>"110011111",
15476=>"101000111",
15477=>"101001111",
15478=>"010111111",
15479=>"000010001",
15480=>"111111101",
15481=>"000000000",
15482=>"001000000",
15483=>"000000010",
15484=>"010000000",
15485=>"111111110",
15486=>"000000000",
15487=>"111111111",
15488=>"100111110",
15489=>"000000000",
15490=>"000000000",
15491=>"000000000",
15492=>"011110111",
15493=>"000000111",
15494=>"000000000",
15495=>"001000000",
15496=>"001011001",
15497=>"000001101",
15498=>"000001010",
15499=>"011111111",
15500=>"111111011",
15501=>"010111010",
15502=>"000000000",
15503=>"111000101",
15504=>"111111111",
15505=>"010010010",
15506=>"001000101",
15507=>"011101110",
15508=>"000101101",
15509=>"010000000",
15510=>"100100100",
15511=>"000000001",
15512=>"110000000",
15513=>"111111101",
15514=>"001000101",
15515=>"111110000",
15516=>"110000010",
15517=>"011110010",
15518=>"000000111",
15519=>"110111110",
15520=>"000000010",
15521=>"000000000",
15522=>"001001000",
15523=>"000010000",
15524=>"000000100",
15525=>"000000000",
15526=>"000001001",
15527=>"100000111",
15528=>"000011011",
15529=>"000001001",
15530=>"111101100",
15531=>"100110110",
15532=>"111111011",
15533=>"111111111",
15534=>"001011011",
15535=>"111111110",
15536=>"111111111",
15537=>"000000110",
15538=>"000010010",
15539=>"011000000",
15540=>"010000010",
15541=>"000000111",
15542=>"111110100",
15543=>"110010000",
15544=>"000000000",
15545=>"001010101",
15546=>"000000000",
15547=>"100000110",
15548=>"001101111",
15549=>"000111111",
15550=>"000001001",
15551=>"000100000",
15552=>"111111111",
15553=>"000010111",
15554=>"000000000",
15555=>"000010000",
15556=>"001001101",
15557=>"010000001",
15558=>"000000001",
15559=>"111111111",
15560=>"001001101",
15561=>"000000001",
15562=>"111111111",
15563=>"000000000",
15564=>"011110111",
15565=>"001011000",
15566=>"111001100",
15567=>"011001111",
15568=>"111111111",
15569=>"110110110",
15570=>"111110101",
15571=>"011101111",
15572=>"111111111",
15573=>"001011011",
15574=>"111111111",
15575=>"110111111",
15576=>"001000001",
15577=>"000110010",
15578=>"000000100",
15579=>"111100000",
15580=>"001111110",
15581=>"111111001",
15582=>"010111111",
15583=>"000000000",
15584=>"110000001",
15585=>"111111111",
15586=>"111000000",
15587=>"011111011",
15588=>"001000000",
15589=>"010111010",
15590=>"001000000",
15591=>"100110110",
15592=>"000000000",
15593=>"000101000",
15594=>"100100110",
15595=>"111111110",
15596=>"000000000",
15597=>"011111011",
15598=>"010010000",
15599=>"001000001",
15600=>"001001101",
15601=>"000000100",
15602=>"011111111",
15603=>"100001101",
15604=>"001001011",
15605=>"110111111",
15606=>"110111110",
15607=>"011000000",
15608=>"001000001",
15609=>"000101000",
15610=>"111000001",
15611=>"101111111",
15612=>"111100111",
15613=>"010000000",
15614=>"000000000",
15615=>"000111111",
15616=>"011011011",
15617=>"001111110",
15618=>"101000000",
15619=>"100111000",
15620=>"001001110",
15621=>"000000110",
15622=>"000000010",
15623=>"000100100",
15624=>"000000000",
15625=>"011001111",
15626=>"001001011",
15627=>"111101010",
15628=>"101100110",
15629=>"111111001",
15630=>"001000001",
15631=>"001111111",
15632=>"000001110",
15633=>"010000101",
15634=>"000111100",
15635=>"111000000",
15636=>"110000000",
15637=>"111110010",
15638=>"111111011",
15639=>"001000111",
15640=>"001100111",
15641=>"011000001",
15642=>"010001111",
15643=>"011001001",
15644=>"001000100",
15645=>"100000100",
15646=>"111000000",
15647=>"000110111",
15648=>"000000000",
15649=>"000001111",
15650=>"111111111",
15651=>"111110110",
15652=>"001011111",
15653=>"110010111",
15654=>"110110010",
15655=>"101010101",
15656=>"110011000",
15657=>"110110000",
15658=>"001000111",
15659=>"010000000",
15660=>"111100000",
15661=>"111011101",
15662=>"101001000",
15663=>"011111100",
15664=>"000000001",
15665=>"011100011",
15666=>"101111001",
15667=>"100000000",
15668=>"000000000",
15669=>"111101000",
15670=>"100010111",
15671=>"000111100",
15672=>"111111010",
15673=>"001000101",
15674=>"000101000",
15675=>"110111111",
15676=>"110001000",
15677=>"010111010",
15678=>"000000101",
15679=>"000000000",
15680=>"100101101",
15681=>"111110010",
15682=>"110001000",
15683=>"011000000",
15684=>"011110000",
15685=>"101000000",
15686=>"000000001",
15687=>"110000010",
15688=>"111111111",
15689=>"001001000",
15690=>"000001001",
15691=>"001000101",
15692=>"111110110",
15693=>"110111100",
15694=>"010110001",
15695=>"110111111",
15696=>"000000000",
15697=>"010011111",
15698=>"111000001",
15699=>"011001011",
15700=>"001000011",
15701=>"110111110",
15702=>"111111011",
15703=>"000000000",
15704=>"000000111",
15705=>"100001000",
15706=>"001111101",
15707=>"010100000",
15708=>"100110110",
15709=>"000011111",
15710=>"111111111",
15711=>"110000000",
15712=>"000000000",
15713=>"000000001",
15714=>"001001011",
15715=>"111110000",
15716=>"100111111",
15717=>"110011100",
15718=>"001001111",
15719=>"110110000",
15720=>"000000000",
15721=>"110000101",
15722=>"000111101",
15723=>"111110000",
15724=>"110110101",
15725=>"000000001",
15726=>"111111000",
15727=>"000100110",
15728=>"011101101",
15729=>"000000000",
15730=>"001100111",
15731=>"111000000",
15732=>"001100110",
15733=>"000001000",
15734=>"000001001",
15735=>"111110001",
15736=>"011011111",
15737=>"110010010",
15738=>"111111001",
15739=>"101000000",
15740=>"010111101",
15741=>"100100100",
15742=>"110000000",
15743=>"001001000",
15744=>"110101110",
15745=>"100100001",
15746=>"111001011",
15747=>"111101111",
15748=>"011111101",
15749=>"000000000",
15750=>"110100111",
15751=>"000001010",
15752=>"100111011",
15753=>"001000000",
15754=>"000000111",
15755=>"010000000",
15756=>"000000100",
15757=>"101000000",
15758=>"000101011",
15759=>"011000000",
15760=>"111111111",
15761=>"010110110",
15762=>"000000010",
15763=>"001000000",
15764=>"000000000",
15765=>"010000000",
15766=>"001111111",
15767=>"010011101",
15768=>"111111111",
15769=>"001110110",
15770=>"110000000",
15771=>"001001000",
15772=>"000000000",
15773=>"001001011",
15774=>"110111111",
15775=>"111010000",
15776=>"100101110",
15777=>"000110110",
15778=>"100000001",
15779=>"001001011",
15780=>"110000011",
15781=>"110111100",
15782=>"110110000",
15783=>"111001101",
15784=>"110000000",
15785=>"000110111",
15786=>"101001111",
15787=>"011000001",
15788=>"001001011",
15789=>"000000011",
15790=>"100100100",
15791=>"110100100",
15792=>"000001001",
15793=>"000111011",
15794=>"000000000",
15795=>"000000011",
15796=>"111111111",
15797=>"000000011",
15798=>"111111111",
15799=>"111110010",
15800=>"011101001",
15801=>"110011100",
15802=>"111010110",
15803=>"011001001",
15804=>"100010000",
15805=>"000110111",
15806=>"000000001",
15807=>"010111111",
15808=>"000000111",
15809=>"000000100",
15810=>"101000010",
15811=>"010111010",
15812=>"011000000",
15813=>"001001111",
15814=>"100000000",
15815=>"101010111",
15816=>"101101001",
15817=>"110111000",
15818=>"001101111",
15819=>"001101001",
15820=>"001001000",
15821=>"110101011",
15822=>"001101010",
15823=>"001111001",
15824=>"111111000",
15825=>"100111010",
15826=>"001010000",
15827=>"111111011",
15828=>"111000001",
15829=>"001100110",
15830=>"111110110",
15831=>"111111111",
15832=>"111110010",
15833=>"111111111",
15834=>"110100000",
15835=>"001000001",
15836=>"110111001",
15837=>"111010000",
15838=>"111110000",
15839=>"111111000",
15840=>"001000101",
15841=>"001001001",
15842=>"111111101",
15843=>"000000101",
15844=>"001000110",
15845=>"110010000",
15846=>"101011000",
15847=>"001001011",
15848=>"111100100",
15849=>"010010110",
15850=>"001000001",
15851=>"001001011",
15852=>"010100000",
15853=>"110110100",
15854=>"110000000",
15855=>"100110011",
15856=>"000000000",
15857=>"010100111",
15858=>"111011110",
15859=>"010011110",
15860=>"100100100",
15861=>"001001111",
15862=>"000000010",
15863=>"001001101",
15864=>"001000000",
15865=>"000001111",
15866=>"001111111",
15867=>"011111111",
15868=>"001011001",
15869=>"000000000",
15870=>"000110111",
15871=>"000000001",
15872=>"011011111",
15873=>"100101011",
15874=>"001001011",
15875=>"000011101",
15876=>"100010100",
15877=>"000000111",
15878=>"011111010",
15879=>"100010111",
15880=>"000110111",
15881=>"000100000",
15882=>"000100100",
15883=>"110000111",
15884=>"110110100",
15885=>"011001100",
15886=>"011000110",
15887=>"000000000",
15888=>"000110110",
15889=>"011000111",
15890=>"001011100",
15891=>"111001010",
15892=>"011111111",
15893=>"101001101",
15894=>"110111111",
15895=>"111110111",
15896=>"001011111",
15897=>"001110110",
15898=>"000111010",
15899=>"100110000",
15900=>"001001101",
15901=>"110100000",
15902=>"000011001",
15903=>"110110000",
15904=>"001010111",
15905=>"110111011",
15906=>"111001010",
15907=>"110100111",
15908=>"111011000",
15909=>"000000000",
15910=>"001011111",
15911=>"101000000",
15912=>"011111111",
15913=>"011111110",
15914=>"000000001",
15915=>"010110100",
15916=>"100110001",
15917=>"100110100",
15918=>"001001101",
15919=>"111111110",
15920=>"111000100",
15921=>"111011011",
15922=>"100001000",
15923=>"110000100",
15924=>"110100000",
15925=>"000100000",
15926=>"100100100",
15927=>"000100100",
15928=>"000011011",
15929=>"000000000",
15930=>"100000000",
15931=>"100001000",
15932=>"110110110",
15933=>"110011011",
15934=>"000000001",
15935=>"100000010",
15936=>"011011111",
15937=>"000010011",
15938=>"110100100",
15939=>"011000000",
15940=>"001011000",
15941=>"000000010",
15942=>"100100000",
15943=>"001111001",
15944=>"000000000",
15945=>"110010100",
15946=>"010011111",
15947=>"010001001",
15948=>"001001110",
15949=>"000000100",
15950=>"001000000",
15951=>"111111110",
15952=>"011011010",
15953=>"101111110",
15954=>"100100000",
15955=>"101101001",
15956=>"111001000",
15957=>"001101111",
15958=>"100000101",
15959=>"010110000",
15960=>"010111110",
15961=>"111100000",
15962=>"101110100",
15963=>"100010001",
15964=>"000010100",
15965=>"011100010",
15966=>"101111010",
15967=>"101111111",
15968=>"000011111",
15969=>"111011000",
15970=>"011010101",
15971=>"110111011",
15972=>"100100100",
15973=>"100100110",
15974=>"110000000",
15975=>"011111011",
15976=>"011010110",
15977=>"000000000",
15978=>"110000110",
15979=>"101110101",
15980=>"011011110",
15981=>"011000000",
15982=>"100000000",
15983=>"100000001",
15984=>"001101100",
15985=>"100100000",
15986=>"100000110",
15987=>"000000110",
15988=>"000000000",
15989=>"000011001",
15990=>"111101001",
15991=>"100011010",
15992=>"110111111",
15993=>"110100001",
15994=>"011000111",
15995=>"111001010",
15996=>"110010100",
15997=>"000000101",
15998=>"100100111",
15999=>"111000000",
16000=>"001001000",
16001=>"111001000",
16002=>"101111000",
16003=>"100111111",
16004=>"110010100",
16005=>"011100000",
16006=>"001010110",
16007=>"110011111",
16008=>"010111111",
16009=>"001100100",
16010=>"100100010",
16011=>"001010001",
16012=>"000111110",
16013=>"000000100",
16014=>"001100000",
16015=>"010000000",
16016=>"100100110",
16017=>"100100000",
16018=>"000000001",
16019=>"011011111",
16020=>"110111010",
16021=>"001000000",
16022=>"000100000",
16023=>"100000110",
16024=>"110100110",
16025=>"011111011",
16026=>"001011111",
16027=>"001100100",
16028=>"110100000",
16029=>"011011100",
16030=>"000101100",
16031=>"111001111",
16032=>"100100001",
16033=>"010010100",
16034=>"011110111",
16035=>"001011111",
16036=>"011010110",
16037=>"000100100",
16038=>"111011010",
16039=>"000110110",
16040=>"111110000",
16041=>"100111110",
16042=>"001001001",
16043=>"011011011",
16044=>"001111111",
16045=>"010100000",
16046=>"010000000",
16047=>"100100101",
16048=>"010100100",
16049=>"011110111",
16050=>"001010000",
16051=>"000000110",
16052=>"111111111",
16053=>"111100000",
16054=>"100000100",
16055=>"011100001",
16056=>"111000010",
16057=>"100110000",
16058=>"100000000",
16059=>"010111111",
16060=>"100100010",
16061=>"001001110",
16062=>"111111111",
16063=>"110010000",
16064=>"001000000",
16065=>"001001100",
16066=>"001001000",
16067=>"010011001",
16068=>"000000000",
16069=>"011101111",
16070=>"100110010",
16071=>"011011011",
16072=>"100000001",
16073=>"110010010",
16074=>"000110100",
16075=>"100100000",
16076=>"011011100",
16077=>"111000100",
16078=>"110011111",
16079=>"100100111",
16080=>"101001000",
16081=>"110100001",
16082=>"100110100",
16083=>"100000000",
16084=>"001000000",
16085=>"000100100",
16086=>"111110010",
16087=>"100000000",
16088=>"000000000",
16089=>"110100000",
16090=>"100111011",
16091=>"001011111",
16092=>"100111111",
16093=>"011011101",
16094=>"000110100",
16095=>"000111001",
16096=>"100100100",
16097=>"011001001",
16098=>"100000000",
16099=>"000100010",
16100=>"000010100",
16101=>"000110000",
16102=>"100100000",
16103=>"110010101",
16104=>"010000000",
16105=>"010010000",
16106=>"111100000",
16107=>"011000000",
16108=>"110100000",
16109=>"000010000",
16110=>"010011010",
16111=>"000000110",
16112=>"010110111",
16113=>"011011110",
16114=>"000111111",
16115=>"100100000",
16116=>"100100111",
16117=>"000111011",
16118=>"000110011",
16119=>"000000010",
16120=>"011001111",
16121=>"100110000",
16122=>"011111100",
16123=>"110011111",
16124=>"001001100",
16125=>"000000100",
16126=>"100110110",
16127=>"010011111",
16128=>"111111001",
16129=>"000111111",
16130=>"100000100",
16131=>"110111111",
16132=>"001011001",
16133=>"000001000",
16134=>"000000110",
16135=>"111111111",
16136=>"010000000",
16137=>"000000000",
16138=>"000000011",
16139=>"010111111",
16140=>"110111111",
16141=>"111111000",
16142=>"000111111",
16143=>"000000000",
16144=>"110000000",
16145=>"000000000",
16146=>"111000000",
16147=>"000100111",
16148=>"111001000",
16149=>"111111111",
16150=>"101001100",
16151=>"111010010",
16152=>"000111111",
16153=>"000000000",
16154=>"000010000",
16155=>"000000111",
16156=>"111101111",
16157=>"000001100",
16158=>"011000010",
16159=>"000111111",
16160=>"000000000",
16161=>"011111010",
16162=>"101000101",
16163=>"101111111",
16164=>"101101001",
16165=>"110110100",
16166=>"000000001",
16167=>"111111111",
16168=>"111110111",
16169=>"001101111",
16170=>"111111111",
16171=>"111100111",
16172=>"000111111",
16173=>"001011001",
16174=>"111100111",
16175=>"110111111",
16176=>"000000010",
16177=>"011011010",
16178=>"111111111",
16179=>"111101111",
16180=>"001000000",
16181=>"011101111",
16182=>"111111111",
16183=>"000000001",
16184=>"111000000",
16185=>"011001000",
16186=>"000000010",
16187=>"111000110",
16188=>"100100110",
16189=>"000111111",
16190=>"000000111",
16191=>"000000000",
16192=>"100000001",
16193=>"101111010",
16194=>"000000111",
16195=>"010000000",
16196=>"110111111",
16197=>"000001000",
16198=>"000000000",
16199=>"010000011",
16200=>"111110111",
16201=>"000000000",
16202=>"111010000",
16203=>"000000000",
16204=>"000000000",
16205=>"110000001",
16206=>"000000111",
16207=>"101111010",
16208=>"111111110",
16209=>"111111001",
16210=>"000000000",
16211=>"001011010",
16212=>"000110111",
16213=>"010110110",
16214=>"000000000",
16215=>"000000000",
16216=>"000000000",
16217=>"001001000",
16218=>"000001100",
16219=>"000001000",
16220=>"111111000",
16221=>"001011000",
16222=>"101101000",
16223=>"101000010",
16224=>"000000000",
16225=>"000100000",
16226=>"111010010",
16227=>"000000000",
16228=>"000100000",
16229=>"100000000",
16230=>"001000010",
16231=>"001000100",
16232=>"000000000",
16233=>"001001111",
16234=>"111100010",
16235=>"110111110",
16236=>"111111101",
16237=>"000000100",
16238=>"110000000",
16239=>"000011101",
16240=>"100100100",
16241=>"111000000",
16242=>"111111110",
16243=>"100000101",
16244=>"111111000",
16245=>"000000000",
16246=>"001111111",
16247=>"101111111",
16248=>"000000000",
16249=>"001111111",
16250=>"000000000",
16251=>"111111000",
16252=>"100100110",
16253=>"110110000",
16254=>"001000001",
16255=>"000000000",
16256=>"110101000",
16257=>"111111000",
16258=>"000000001",
16259=>"010001001",
16260=>"111111111",
16261=>"001000011",
16262=>"110001011",
16263=>"001001001",
16264=>"011011111",
16265=>"001000000",
16266=>"100000000",
16267=>"111010000",
16268=>"000000000",
16269=>"000000001",
16270=>"000111101",
16271=>"000100110",
16272=>"011011011",
16273=>"010111111",
16274=>"111111000",
16275=>"110111111",
16276=>"000001111",
16277=>"111110010",
16278=>"111011000",
16279=>"000000000",
16280=>"000001001",
16281=>"000110111",
16282=>"110000000",
16283=>"111000000",
16284=>"111100010",
16285=>"000110111",
16286=>"111110000",
16287=>"101000000",
16288=>"011011100",
16289=>"001111010",
16290=>"111111111",
16291=>"010000010",
16292=>"111111111",
16293=>"000000000",
16294=>"111100101",
16295=>"111111101",
16296=>"000000111",
16297=>"000111111",
16298=>"111000100",
16299=>"000111111",
16300=>"001000011",
16301=>"000010111",
16302=>"110111100",
16303=>"001101111",
16304=>"000000000",
16305=>"001000100",
16306=>"000000000",
16307=>"010100100",
16308=>"000011011",
16309=>"111111111",
16310=>"001000100",
16311=>"111101111",
16312=>"011001001",
16313=>"000100111",
16314=>"000110101",
16315=>"000110010",
16316=>"000100000",
16317=>"111000000",
16318=>"000000000",
16319=>"011011111",
16320=>"000110000",
16321=>"000000001",
16322=>"111101011",
16323=>"111011111",
16324=>"000000000",
16325=>"010101111",
16326=>"000000011",
16327=>"111110100",
16328=>"111000111",
16329=>"000000001",
16330=>"010110111",
16331=>"000000000",
16332=>"000000000",
16333=>"001001011",
16334=>"000000011",
16335=>"111101011",
16336=>"000000000",
16337=>"001000000",
16338=>"001000001",
16339=>"000000001",
16340=>"100110100",
16341=>"101011111",
16342=>"110101000",
16343=>"000000011",
16344=>"111111100",
16345=>"001100111",
16346=>"110000001",
16347=>"111000100",
16348=>"000000011",
16349=>"100110111",
16350=>"000000000",
16351=>"111010111",
16352=>"000011001",
16353=>"111001010",
16354=>"101111111",
16355=>"000100100",
16356=>"111000000",
16357=>"001111111",
16358=>"011000000",
16359=>"110110010",
16360=>"111000001",
16361=>"011111101",
16362=>"000000000",
16363=>"001001111",
16364=>"111111111",
16365=>"111111101",
16366=>"000000000",
16367=>"111001000",
16368=>"000000000",
16369=>"111111111",
16370=>"111001001",
16371=>"000111011",
16372=>"110110110",
16373=>"111000001",
16374=>"101001001",
16375=>"000001000",
16376=>"110110010",
16377=>"111111111",
16378=>"011111110",
16379=>"001000111",
16380=>"000000000",
16381=>"111111011",
16382=>"110110101",
16383=>"111101111",
16384=>"000000000",
16385=>"000000001",
16386=>"010000001",
16387=>"110000010",
16388=>"011011010",
16389=>"100000011",
16390=>"111010110",
16391=>"000111010",
16392=>"110011000",
16393=>"001000000",
16394=>"000011110",
16395=>"101000000",
16396=>"111000000",
16397=>"111101101",
16398=>"100010110",
16399=>"001000001",
16400=>"000000110",
16401=>"000110001",
16402=>"101000000",
16403=>"111000001",
16404=>"111001111",
16405=>"100000000",
16406=>"101111000",
16407=>"111010001",
16408=>"000000001",
16409=>"111111111",
16410=>"111100101",
16411=>"000110010",
16412=>"000001101",
16413=>"101000000",
16414=>"110100100",
16415=>"111000000",
16416=>"110111100",
16417=>"111111110",
16418=>"000000001",
16419=>"100110000",
16420=>"111111111",
16421=>"100001111",
16422=>"000000111",
16423=>"111110001",
16424=>"000111110",
16425=>"000110110",
16426=>"111000001",
16427=>"000000111",
16428=>"011111011",
16429=>"111000000",
16430=>"100101011",
16431=>"100111111",
16432=>"110110101",
16433=>"001111111",
16434=>"110111101",
16435=>"010110110",
16436=>"110000111",
16437=>"010110011",
16438=>"001010000",
16439=>"100000000",
16440=>"010111011",
16441=>"001000101",
16442=>"011001001",
16443=>"000010101",
16444=>"010011100",
16445=>"111011000",
16446=>"111000000",
16447=>"100001000",
16448=>"010110000",
16449=>"110000101",
16450=>"101010010",
16451=>"011010011",
16452=>"100000101",
16453=>"001000000",
16454=>"001111010",
16455=>"110000000",
16456=>"101001101",
16457=>"110010000",
16458=>"001001000",
16459=>"000000110",
16460=>"111110110",
16461=>"010011111",
16462=>"000100110",
16463=>"000001110",
16464=>"000000110",
16465=>"111001000",
16466=>"011000010",
16467=>"011011100",
16468=>"101100110",
16469=>"111100000",
16470=>"000111111",
16471=>"111101111",
16472=>"000000100",
16473=>"011000010",
16474=>"111001001",
16475=>"111011110",
16476=>"100001001",
16477=>"110001011",
16478=>"001111111",
16479=>"111100001",
16480=>"001001111",
16481=>"000100000",
16482=>"101111111",
16483=>"101000100",
16484=>"000110100",
16485=>"011100100",
16486=>"101000010",
16487=>"010101111",
16488=>"000011111",
16489=>"110000111",
16490=>"011111000",
16491=>"000000111",
16492=>"110100111",
16493=>"000110110",
16494=>"111000000",
16495=>"101111111",
16496=>"100111101",
16497=>"110110011",
16498=>"001100000",
16499=>"000001001",
16500=>"000110000",
16501=>"100000111",
16502=>"000000010",
16503=>"100001110",
16504=>"111000110",
16505=>"010110001",
16506=>"111111001",
16507=>"000001000",
16508=>"100110100",
16509=>"100100101",
16510=>"110111011",
16511=>"001001110",
16512=>"011010010",
16513=>"111000001",
16514=>"101011100",
16515=>"111101000",
16516=>"110000100",
16517=>"001111111",
16518=>"110000100",
16519=>"001100001",
16520=>"001101011",
16521=>"000110010",
16522=>"000001001",
16523=>"000000000",
16524=>"000000100",
16525=>"001001111",
16526=>"110111000",
16527=>"100000100",
16528=>"101111111",
16529=>"110000111",
16530=>"010010101",
16531=>"000001111",
16532=>"000111110",
16533=>"110110000",
16534=>"000111111",
16535=>"110000000",
16536=>"001000110",
16537=>"110001000",
16538=>"010000000",
16539=>"000010010",
16540=>"101000010",
16541=>"001010010",
16542=>"110100000",
16543=>"101001000",
16544=>"101001100",
16545=>"111110111",
16546=>"001001111",
16547=>"110000001",
16548=>"110111111",
16549=>"000011111",
16550=>"101001001",
16551=>"101000000",
16552=>"001110111",
16553=>"000000111",
16554=>"111111001",
16555=>"001110001",
16556=>"111101101",
16557=>"001000000",
16558=>"110011011",
16559=>"000000010",
16560=>"111000000",
16561=>"000001010",
16562=>"111110000",
16563=>"100001101",
16564=>"111101101",
16565=>"000001001",
16566=>"000011100",
16567=>"110010000",
16568=>"011000101",
16569=>"100010110",
16570=>"011001110",
16571=>"111011001",
16572=>"011101010",
16573=>"111111011",
16574=>"001000001",
16575=>"110110111",
16576=>"101001000",
16577=>"000010000",
16578=>"010110000",
16579=>"001011111",
16580=>"000010111",
16581=>"111110101",
16582=>"111110011",
16583=>"010111111",
16584=>"101101010",
16585=>"000010100",
16586=>"001011000",
16587=>"001110111",
16588=>"000001110",
16589=>"011110110",
16590=>"111110000",
16591=>"010010111",
16592=>"000011000",
16593=>"000111111",
16594=>"000011010",
16595=>"101001100",
16596=>"100110010",
16597=>"111000100",
16598=>"101001101",
16599=>"000000001",
16600=>"101001001",
16601=>"000000000",
16602=>"011000000",
16603=>"001000010",
16604=>"011110000",
16605=>"000000111",
16606=>"000111101",
16607=>"000000110",
16608=>"001000110",
16609=>"111111010",
16610=>"110001001",
16611=>"000111111",
16612=>"001000000",
16613=>"110110110",
16614=>"000111110",
16615=>"101101101",
16616=>"111110000",
16617=>"111000000",
16618=>"000100100",
16619=>"111100000",
16620=>"110000000",
16621=>"010001001",
16622=>"110000100",
16623=>"010111101",
16624=>"000001000",
16625=>"111011101",
16626=>"100001000",
16627=>"000011000",
16628=>"100001011",
16629=>"000000010",
16630=>"000100111",
16631=>"010101001",
16632=>"101000100",
16633=>"111101111",
16634=>"011111101",
16635=>"000111110",
16636=>"111111111",
16637=>"000010000",
16638=>"110100100",
16639=>"000111111",
16640=>"100100100",
16641=>"000000000",
16642=>"010010010",
16643=>"000000011",
16644=>"111111111",
16645=>"000001011",
16646=>"001111011",
16647=>"000101000",
16648=>"001111111",
16649=>"000100001",
16650=>"110110100",
16651=>"101001000",
16652=>"101101101",
16653=>"101111010",
16654=>"110000100",
16655=>"000010001",
16656=>"100000101",
16657=>"001011010",
16658=>"010010000",
16659=>"000110111",
16660=>"111111111",
16661=>"001111111",
16662=>"100100100",
16663=>"000101001",
16664=>"110010000",
16665=>"111111010",
16666=>"000000100",
16667=>"110110011",
16668=>"110001110",
16669=>"000000010",
16670=>"001101111",
16671=>"000010011",
16672=>"111111111",
16673=>"111111010",
16674=>"000000101",
16675=>"101001101",
16676=>"010111000",
16677=>"001001111",
16678=>"010011111",
16679=>"111111011",
16680=>"111101000",
16681=>"001111111",
16682=>"100000100",
16683=>"000000001",
16684=>"000100100",
16685=>"111101100",
16686=>"000101111",
16687=>"000100101",
16688=>"101001000",
16689=>"111110010",
16690=>"110000000",
16691=>"101000000",
16692=>"001001111",
16693=>"000101100",
16694=>"000100100",
16695=>"101101000",
16696=>"000000000",
16697=>"000000000",
16698=>"000000000",
16699=>"111111111",
16700=>"001001011",
16701=>"011011001",
16702=>"100000000",
16703=>"100101001",
16704=>"111001001",
16705=>"001101101",
16706=>"101100000",
16707=>"100001000",
16708=>"111110011",
16709=>"000001111",
16710=>"001001000",
16711=>"001101110",
16712=>"011011001",
16713=>"101101001",
16714=>"000101101",
16715=>"011001101",
16716=>"000000100",
16717=>"011011000",
16718=>"111001000",
16719=>"000000001",
16720=>"101101111",
16721=>"110000001",
16722=>"000011000",
16723=>"110000000",
16724=>"010111101",
16725=>"011101011",
16726=>"011011010",
16727=>"101000100",
16728=>"010000100",
16729=>"111110010",
16730=>"011011011",
16731=>"101110111",
16732=>"101101100",
16733=>"110110100",
16734=>"101111111",
16735=>"001000100",
16736=>"010010010",
16737=>"001101111",
16738=>"110010101",
16739=>"110110110",
16740=>"011011011",
16741=>"101100110",
16742=>"001111001",
16743=>"010010000",
16744=>"101000001",
16745=>"000000000",
16746=>"001000001",
16747=>"000011010",
16748=>"111101100",
16749=>"010000000",
16750=>"101101100",
16751=>"010010000",
16752=>"101001100",
16753=>"000111100",
16754=>"100000000",
16755=>"000000111",
16756=>"000000101",
16757=>"000100100",
16758=>"101000000",
16759=>"000010111",
16760=>"100111100",
16761=>"010100001",
16762=>"111000000",
16763=>"011001001",
16764=>"011001001",
16765=>"011001000",
16766=>"101001111",
16767=>"010010011",
16768=>"101111000",
16769=>"010010000",
16770=>"000000110",
16771=>"001001111",
16772=>"101101001",
16773=>"000111010",
16774=>"100100110",
16775=>"110100100",
16776=>"110111011",
16777=>"111010010",
16778=>"000100100",
16779=>"101111011",
16780=>"000000000",
16781=>"010010111",
16782=>"101100111",
16783=>"111000011",
16784=>"111001111",
16785=>"000010000",
16786=>"001000001",
16787=>"101001000",
16788=>"111000000",
16789=>"000000100",
16790=>"111100101",
16791=>"010100110",
16792=>"001111111",
16793=>"110111000",
16794=>"000000110",
16795=>"000000110",
16796=>"100100100",
16797=>"010110010",
16798=>"101101000",
16799=>"010011000",
16800=>"100110000",
16801=>"000010000",
16802=>"100101011",
16803=>"000000000",
16804=>"000101101",
16805=>"011111001",
16806=>"111101110",
16807=>"000100111",
16808=>"101101001",
16809=>"000000111",
16810=>"000000000",
16811=>"111101010",
16812=>"101111111",
16813=>"110010000",
16814=>"011110100",
16815=>"101011001",
16816=>"000111111",
16817=>"011100001",
16818=>"000010010",
16819=>"011011011",
16820=>"000000000",
16821=>"101101111",
16822=>"111011011",
16823=>"101111011",
16824=>"110100110",
16825=>"011001000",
16826=>"100000000",
16827=>"101111111",
16828=>"110010011",
16829=>"111010011",
16830=>"100100100",
16831=>"000101101",
16832=>"001111000",
16833=>"000100100",
16834=>"111110010",
16835=>"110100111",
16836=>"111101000",
16837=>"011011000",
16838=>"110101000",
16839=>"010100100",
16840=>"111000010",
16841=>"000010110",
16842=>"000000111",
16843=>"000000100",
16844=>"100111111",
16845=>"110100100",
16846=>"011111111",
16847=>"110101000",
16848=>"111110000",
16849=>"010011010",
16850=>"101000001",
16851=>"100001000",
16852=>"111111111",
16853=>"001111111",
16854=>"110111001",
16855=>"101000110",
16856=>"001111101",
16857=>"010000000",
16858=>"010001000",
16859=>"011000000",
16860=>"000111110",
16861=>"000100110",
16862=>"100101111",
16863=>"111111100",
16864=>"101101101",
16865=>"110000000",
16866=>"101111111",
16867=>"111000011",
16868=>"000000000",
16869=>"111111111",
16870=>"101000000",
16871=>"101111010",
16872=>"000000000",
16873=>"111111101",
16874=>"101101001",
16875=>"001100111",
16876=>"100101101",
16877=>"110111011",
16878=>"111011011",
16879=>"001111101",
16880=>"000000001",
16881=>"110110110",
16882=>"101101111",
16883=>"000000100",
16884=>"001101101",
16885=>"010010110",
16886=>"011010111",
16887=>"000000000",
16888=>"111001001",
16889=>"001000000",
16890=>"010010011",
16891=>"111000001",
16892=>"000111111",
16893=>"100100111",
16894=>"111110111",
16895=>"100110000",
16896=>"011100000",
16897=>"111111000",
16898=>"111000101",
16899=>"101111110",
16900=>"001111011",
16901=>"110111110",
16902=>"011000000",
16903=>"000000000",
16904=>"000010010",
16905=>"010010000",
16906=>"110000000",
16907=>"100000001",
16908=>"101111011",
16909=>"111111000",
16910=>"101011100",
16911=>"000000000",
16912=>"001111011",
16913=>"111000000",
16914=>"001001111",
16915=>"000010001",
16916=>"000000010",
16917=>"110110000",
16918=>"001001101",
16919=>"001000110",
16920=>"101101000",
16921=>"000000000",
16922=>"001011010",
16923=>"111110101",
16924=>"101111111",
16925=>"010111111",
16926=>"111111011",
16927=>"111000011",
16928=>"001000000",
16929=>"101111111",
16930=>"001000101",
16931=>"000100111",
16932=>"001000010",
16933=>"111010000",
16934=>"000000111",
16935=>"000000110",
16936=>"101111000",
16937=>"000101100",
16938=>"011000010",
16939=>"001101111",
16940=>"000100111",
16941=>"100111111",
16942=>"100111111",
16943=>"000110110",
16944=>"001111100",
16945=>"000011011",
16946=>"010010010",
16947=>"010110000",
16948=>"000000101",
16949=>"000000100",
16950=>"111111100",
16951=>"000001111",
16952=>"111100000",
16953=>"001000111",
16954=>"111000100",
16955=>"000000100",
16956=>"100111001",
16957=>"111111111",
16958=>"101000101",
16959=>"001000010",
16960=>"111001000",
16961=>"110010000",
16962=>"111111000",
16963=>"010001000",
16964=>"000010000",
16965=>"000000010",
16966=>"000010010",
16967=>"001111101",
16968=>"000011011",
16969=>"111111100",
16970=>"101101101",
16971=>"001001111",
16972=>"111010101",
16973=>"001100000",
16974=>"110111110",
16975=>"100111111",
16976=>"110010000",
16977=>"111111111",
16978=>"000100111",
16979=>"001000001",
16980=>"101001101",
16981=>"000010110",
16982=>"111001000",
16983=>"111111000",
16984=>"100000000",
16985=>"110000001",
16986=>"000001111",
16987=>"100000011",
16988=>"011010000",
16989=>"000001011",
16990=>"011111000",
16991=>"110001000",
16992=>"000000000",
16993=>"111110000",
16994=>"000000000",
16995=>"000101111",
16996=>"101101000",
16997=>"111101001",
16998=>"011110000",
16999=>"000110010",
17000=>"100101001",
17001=>"010000100",
17002=>"011111111",
17003=>"000010000",
17004=>"111101101",
17005=>"011011001",
17006=>"000110011",
17007=>"111100111",
17008=>"110110010",
17009=>"111000000",
17010=>"111111001",
17011=>"000000010",
17012=>"001111011",
17013=>"000100100",
17014=>"100110101",
17015=>"101100001",
17016=>"110000101",
17017=>"000000000",
17018=>"111111111",
17019=>"111111000",
17020=>"110111011",
17021=>"100000000",
17022=>"100110111",
17023=>"010010000",
17024=>"010101111",
17025=>"111010000",
17026=>"001010101",
17027=>"001111111",
17028=>"000000011",
17029=>"000000101",
17030=>"011010011",
17031=>"000000001",
17032=>"001011010",
17033=>"101101101",
17034=>"000000000",
17035=>"000111101",
17036=>"111011000",
17037=>"101000111",
17038=>"111010000",
17039=>"000000101",
17040=>"000100110",
17041=>"111000000",
17042=>"011110000",
17043=>"000000001",
17044=>"000010110",
17045=>"111111001",
17046=>"001000101",
17047=>"001001011",
17048=>"000101000",
17049=>"000000111",
17050=>"111010000",
17051=>"000100100",
17052=>"000011000",
17053=>"000001111",
17054=>"000111111",
17055=>"000000111",
17056=>"110110011",
17057=>"000000111",
17058=>"011111000",
17059=>"100101111",
17060=>"111111111",
17061=>"000001110",
17062=>"000001111",
17063=>"011111000",
17064=>"111011111",
17065=>"111111000",
17066=>"111111000",
17067=>"100100100",
17068=>"111001111",
17069=>"010010000",
17070=>"011011100",
17071=>"000101111",
17072=>"000000001",
17073=>"001100110",
17074=>"000101000",
17075=>"001100010",
17076=>"110011111",
17077=>"011110100",
17078=>"101110110",
17079=>"001000000",
17080=>"100111100",
17081=>"000110010",
17082=>"011010100",
17083=>"111111110",
17084=>"000000001",
17085=>"111111000",
17086=>"111011100",
17087=>"110000000",
17088=>"010011111",
17089=>"000000111",
17090=>"110110011",
17091=>"011011011",
17092=>"000000001",
17093=>"001010101",
17094=>"010000000",
17095=>"110101000",
17096=>"010000000",
17097=>"000000100",
17098=>"000001000",
17099=>"111111010",
17100=>"100000001",
17101=>"101111110",
17102=>"000001111",
17103=>"001111111",
17104=>"000001111",
17105=>"100110011",
17106=>"110010011",
17107=>"001001011",
17108=>"001101111",
17109=>"100001011",
17110=>"111110000",
17111=>"001000111",
17112=>"000000011",
17113=>"111111010",
17114=>"111100100",
17115=>"100000100",
17116=>"001100011",
17117=>"001111111",
17118=>"110001110",
17119=>"101001011",
17120=>"111111000",
17121=>"111111001",
17122=>"000000111",
17123=>"101110100",
17124=>"101000000",
17125=>"110111111",
17126=>"000000010",
17127=>"001110011",
17128=>"100111111",
17129=>"100100101",
17130=>"011010000",
17131=>"000000000",
17132=>"111110000",
17133=>"011100111",
17134=>"010000000",
17135=>"000101111",
17136=>"100000101",
17137=>"100110111",
17138=>"011101011",
17139=>"001010010",
17140=>"010001001",
17141=>"010000111",
17142=>"000000000",
17143=>"000000110",
17144=>"000011010",
17145=>"001110000",
17146=>"000010010",
17147=>"101110111",
17148=>"000010000",
17149=>"000000111",
17150=>"000000000",
17151=>"000101111",
17152=>"000011001",
17153=>"111000000",
17154=>"001001000",
17155=>"001111010",
17156=>"010110111",
17157=>"111000101",
17158=>"000111111",
17159=>"000110110",
17160=>"111001000",
17161=>"000001000",
17162=>"100000110",
17163=>"111111110",
17164=>"111001000",
17165=>"101000000",
17166=>"100100000",
17167=>"000101001",
17168=>"000101101",
17169=>"000001100",
17170=>"000001110",
17171=>"111110111",
17172=>"110111111",
17173=>"111001110",
17174=>"001110000",
17175=>"101101111",
17176=>"101101100",
17177=>"000111110",
17178=>"111000000",
17179=>"000001111",
17180=>"100111111",
17181=>"101010111",
17182=>"111111000",
17183=>"000000001",
17184=>"000111110",
17185=>"110000000",
17186=>"111110001",
17187=>"000000001",
17188=>"001111111",
17189=>"011110100",
17190=>"001000111",
17191=>"000100000",
17192=>"110110100",
17193=>"000100110",
17194=>"000011110",
17195=>"111001001",
17196=>"000110101",
17197=>"111111001",
17198=>"100010011",
17199=>"000010111",
17200=>"111111000",
17201=>"100110100",
17202=>"000111000",
17203=>"111110111",
17204=>"000000111",
17205=>"011011010",
17206=>"000100000",
17207=>"000000010",
17208=>"111111000",
17209=>"000000010",
17210=>"010000101",
17211=>"001001000",
17212=>"100110011",
17213=>"111010110",
17214=>"000000101",
17215=>"010000001",
17216=>"111111000",
17217=>"111100000",
17218=>"111111111",
17219=>"100011110",
17220=>"111000000",
17221=>"000001101",
17222=>"001111110",
17223=>"111000001",
17224=>"000000000",
17225=>"000110111",
17226=>"000111111",
17227=>"001001010",
17228=>"000111111",
17229=>"000110101",
17230=>"001011111",
17231=>"100010111",
17232=>"111001001",
17233=>"111111000",
17234=>"000000101",
17235=>"011011001",
17236=>"111101001",
17237=>"010000110",
17238=>"000111100",
17239=>"000111101",
17240=>"111001000",
17241=>"000100111",
17242=>"000001101",
17243=>"111110001",
17244=>"000110000",
17245=>"000011001",
17246=>"111111000",
17247=>"111110111",
17248=>"000000000",
17249=>"001000010",
17250=>"111001000",
17251=>"001101100",
17252=>"000000111",
17253=>"000010011",
17254=>"000110110",
17255=>"000010110",
17256=>"001011011",
17257=>"001101111",
17258=>"000000111",
17259=>"000100110",
17260=>"000000001",
17261=>"001000101",
17262=>"000000111",
17263=>"000001101",
17264=>"011110111",
17265=>"000010111",
17266=>"000011001",
17267=>"001111001",
17268=>"111110011",
17269=>"011001100",
17270=>"111111110",
17271=>"110000000",
17272=>"101101110",
17273=>"000000000",
17274=>"001000000",
17275=>"101001000",
17276=>"001100100",
17277=>"000100100",
17278=>"000001011",
17279=>"101000011",
17280=>"101000000",
17281=>"000111000",
17282=>"000111011",
17283=>"000001011",
17284=>"000111101",
17285=>"111011000",
17286=>"100011001",
17287=>"000000001",
17288=>"000110101",
17289=>"001000011",
17290=>"000110111",
17291=>"000000000",
17292=>"011000000",
17293=>"111011111",
17294=>"000101001",
17295=>"000001001",
17296=>"000011101",
17297=>"000000000",
17298=>"100000111",
17299=>"000000000",
17300=>"000000111",
17301=>"000001001",
17302=>"101111000",
17303=>"010100100",
17304=>"000111111",
17305=>"111111110",
17306=>"111111111",
17307=>"111000001",
17308=>"000111011",
17309=>"000010000",
17310=>"111111100",
17311=>"000000111",
17312=>"001010001",
17313=>"011010111",
17314=>"000000000",
17315=>"100010000",
17316=>"010000000",
17317=>"001111000",
17318=>"001001011",
17319=>"000110100",
17320=>"000000000",
17321=>"111111101",
17322=>"111101001",
17323=>"000010100",
17324=>"100100110",
17325=>"000100111",
17326=>"010110110",
17327=>"111001000",
17328=>"000110010",
17329=>"000001000",
17330=>"111111000",
17331=>"011011100",
17332=>"000110111",
17333=>"110101101",
17334=>"010000001",
17335=>"010111101",
17336=>"000011111",
17337=>"000000000",
17338=>"000010100",
17339=>"110111000",
17340=>"000000000",
17341=>"111001001",
17342=>"100000000",
17343=>"000000010",
17344=>"001011110",
17345=>"000001010",
17346=>"111110001",
17347=>"000111111",
17348=>"000000000",
17349=>"111111110",
17350=>"000000000",
17351=>"111111000",
17352=>"001101111",
17353=>"000100100",
17354=>"000100110",
17355=>"001110110",
17356=>"000010010",
17357=>"000001010",
17358=>"000000001",
17359=>"101101101",
17360=>"101000001",
17361=>"010011001",
17362=>"000000000",
17363=>"001101001",
17364=>"001111111",
17365=>"000000000",
17366=>"000111110",
17367=>"110110100",
17368=>"000011000",
17369=>"000110101",
17370=>"000000100",
17371=>"111001101",
17372=>"110111011",
17373=>"001101101",
17374=>"000000000",
17375=>"000010110",
17376=>"001000111",
17377=>"111001000",
17378=>"111000000",
17379=>"011010100",
17380=>"000001111",
17381=>"111000001",
17382=>"110000000",
17383=>"000111110",
17384=>"000001001",
17385=>"011111111",
17386=>"001000011",
17387=>"000001000",
17388=>"111101001",
17389=>"111101101",
17390=>"010001000",
17391=>"010001101",
17392=>"001001001",
17393=>"000111101",
17394=>"000000000",
17395=>"000011111",
17396=>"000110111",
17397=>"111001101",
17398=>"000010110",
17399=>"010000010",
17400=>"111011000",
17401=>"001001011",
17402=>"010111111",
17403=>"000110111",
17404=>"000111110",
17405=>"111000111",
17406=>"000111111",
17407=>"000110110",
17408=>"110101111",
17409=>"011011111",
17410=>"100100111",
17411=>"100011011",
17412=>"000000000",
17413=>"001000010",
17414=>"001001100",
17415=>"001001001",
17416=>"111100111",
17417=>"100001001",
17418=>"000100110",
17419=>"011011011",
17420=>"111111111",
17421=>"011010011",
17422=>"110011001",
17423=>"011011000",
17424=>"011010000",
17425=>"011001011",
17426=>"100110111",
17427=>"011000000",
17428=>"100001100",
17429=>"100100111",
17430=>"110101100",
17431=>"011111110",
17432=>"000000101",
17433=>"110000101",
17434=>"000000111",
17435=>"101101111",
17436=>"000100111",
17437=>"110010001",
17438=>"111100100",
17439=>"100010000",
17440=>"111100111",
17441=>"011111110",
17442=>"000011100",
17443=>"011011011",
17444=>"000001000",
17445=>"111000001",
17446=>"001011000",
17447=>"011111100",
17448=>"110110100",
17449=>"011001000",
17450=>"010000111",
17451=>"011011100",
17452=>"011001001",
17453=>"100001111",
17454=>"111001000",
17455=>"000100111",
17456=>"110111011",
17457=>"100001000",
17458=>"000000000",
17459=>"100110100",
17460=>"101111001",
17461=>"011011100",
17462=>"110010000",
17463=>"110110111",
17464=>"111110110",
17465=>"100100111",
17466=>"011110000",
17467=>"011111000",
17468=>"011111010",
17469=>"101011100",
17470=>"101000001",
17471=>"001101001",
17472=>"100100010",
17473=>"000000000",
17474=>"100100001",
17475=>"110000110",
17476=>"001011000",
17477=>"100110000",
17478=>"000100010",
17479=>"010011000",
17480=>"000000001",
17481=>"110111110",
17482=>"100100111",
17483=>"100100000",
17484=>"100100100",
17485=>"111110100",
17486=>"110011110",
17487=>"001111111",
17488=>"111101100",
17489=>"000111111",
17490=>"001000000",
17491=>"000000001",
17492=>"111000000",
17493=>"110111101",
17494=>"111110011",
17495=>"001001011",
17496=>"000110000",
17497=>"000110010",
17498=>"010011001",
17499=>"011011100",
17500=>"100001100",
17501=>"001001001",
17502=>"111101100",
17503=>"101101001",
17504=>"011011000",
17505=>"111100111",
17506=>"100000011",
17507=>"110110110",
17508=>"111101111",
17509=>"110100000",
17510=>"000110100",
17511=>"110111110",
17512=>"011110001",
17513=>"000001001",
17514=>"001000000",
17515=>"010000000",
17516=>"000011011",
17517=>"111101001",
17518=>"110110011",
17519=>"001011000",
17520=>"111111101",
17521=>"010111111",
17522=>"000100110",
17523=>"000001000",
17524=>"011011000",
17525=>"100000000",
17526=>"100001000",
17527=>"011010000",
17528=>"000100001",
17529=>"001101000",
17530=>"111101000",
17531=>"011010011",
17532=>"100001000",
17533=>"100000000",
17534=>"100100111",
17535=>"000000101",
17536=>"001000100",
17537=>"100100100",
17538=>"000001000",
17539=>"011001011",
17540=>"011010000",
17541=>"101100111",
17542=>"010001010",
17543=>"000100100",
17544=>"111111001",
17545=>"010111011",
17546=>"110111111",
17547=>"111101100",
17548=>"111111100",
17549=>"000000010",
17550=>"110100110",
17551=>"000000001",
17552=>"000001000",
17553=>"100111110",
17554=>"011011001",
17555=>"011110010",
17556=>"000011111",
17557=>"111100110",
17558=>"000110001",
17559=>"001001011",
17560=>"000001000",
17561=>"011011000",
17562=>"100100110",
17563=>"000000111",
17564=>"110110111",
17565=>"011000001",
17566=>"100000111",
17567=>"000001111",
17568=>"000100000",
17569=>"101101111",
17570=>"100011110",
17571=>"000000111",
17572=>"100100101",
17573=>"110011011",
17574=>"011011000",
17575=>"111011110",
17576=>"111100111",
17577=>"011011110",
17578=>"100110111",
17579=>"111100001",
17580=>"011111101",
17581=>"100110001",
17582=>"101101101",
17583=>"001001000",
17584=>"101011111",
17585=>"000001001",
17586=>"000011000",
17587=>"000000100",
17588=>"000001000",
17589=>"000100100",
17590=>"001010010",
17591=>"111111011",
17592=>"100000000",
17593=>"011011100",
17594=>"111010011",
17595=>"110110111",
17596=>"100111111",
17597=>"101111101",
17598=>"101111110",
17599=>"001011011",
17600=>"110100101",
17601=>"010110111",
17602=>"100000000",
17603=>"110100110",
17604=>"000011011",
17605=>"110111100",
17606=>"000001001",
17607=>"000000101",
17608=>"000100100",
17609=>"001000000",
17610=>"100110100",
17611=>"100100111",
17612=>"110100000",
17613=>"001001000",
17614=>"100000000",
17615=>"001000110",
17616=>"110100000",
17617=>"111011011",
17618=>"000010011",
17619=>"110110111",
17620=>"000000000",
17621=>"001011000",
17622=>"000011000",
17623=>"111100101",
17624=>"111011001",
17625=>"000100010",
17626=>"101111110",
17627=>"000100111",
17628=>"101001010",
17629=>"010011011",
17630=>"011000000",
17631=>"011110000",
17632=>"111110111",
17633=>"100100110",
17634=>"001000000",
17635=>"001100100",
17636=>"110100111",
17637=>"011011000",
17638=>"011100000",
17639=>"000000000",
17640=>"000010001",
17641=>"111111110",
17642=>"100000000",
17643=>"101111111",
17644=>"011001100",
17645=>"000010011",
17646=>"000100000",
17647=>"111011001",
17648=>"011011000",
17649=>"000110100",
17650=>"111001100",
17651=>"111111011",
17652=>"110111101",
17653=>"000010111",
17654=>"000001001",
17655=>"000001000",
17656=>"000110000",
17657=>"010000000",
17658=>"000110000",
17659=>"110111000",
17660=>"100100111",
17661=>"001001000",
17662=>"000000000",
17663=>"100000111",
17664=>"111111011",
17665=>"000110100",
17666=>"001100100",
17667=>"000100011",
17668=>"101110001",
17669=>"001101000",
17670=>"000111111",
17671=>"010010111",
17672=>"000000111",
17673=>"000100111",
17674=>"010011100",
17675=>"111011011",
17676=>"101111001",
17677=>"000010000",
17678=>"000000000",
17679=>"101111100",
17680=>"100000100",
17681=>"001001011",
17682=>"011000000",
17683=>"010100011",
17684=>"101101111",
17685=>"010000100",
17686=>"110111001",
17687=>"111111111",
17688=>"101101100",
17689=>"110111111",
17690=>"001000010",
17691=>"110110111",
17692=>"000111110",
17693=>"111110000",
17694=>"000000000",
17695=>"001011000",
17696=>"011000101",
17697=>"011011110",
17698=>"011000000",
17699=>"000000110",
17700=>"101111101",
17701=>"100000000",
17702=>"000100101",
17703=>"000011111",
17704=>"001001111",
17705=>"010110111",
17706=>"000001111",
17707=>"010000000",
17708=>"000000000",
17709=>"100110100",
17710=>"111001001",
17711=>"110000000",
17712=>"011001001",
17713=>"110111001",
17714=>"111001000",
17715=>"001000000",
17716=>"000100011",
17717=>"101000010",
17718=>"000000000",
17719=>"110110011",
17720=>"011011010",
17721=>"111110010",
17722=>"101100110",
17723=>"000100000",
17724=>"000011011",
17725=>"110011111",
17726=>"001000000",
17727=>"110111011",
17728=>"110100100",
17729=>"011001111",
17730=>"001010001",
17731=>"111011011",
17732=>"111100100",
17733=>"001000000",
17734=>"000100011",
17735=>"001001000",
17736=>"000000010",
17737=>"000111111",
17738=>"011000001",
17739=>"001100110",
17740=>"000000000",
17741=>"111111101",
17742=>"110111111",
17743=>"000011100",
17744=>"011111000",
17745=>"110100110",
17746=>"100001010",
17747=>"111101101",
17748=>"011000000",
17749=>"100011111",
17750=>"111111111",
17751=>"011111110",
17752=>"100010111",
17753=>"000000000",
17754=>"000100110",
17755=>"101011110",
17756=>"001001010",
17757=>"011000000",
17758=>"101100111",
17759=>"000000000",
17760=>"100011001",
17761=>"111110110",
17762=>"001100100",
17763=>"110010110",
17764=>"010000001",
17765=>"000001001",
17766=>"111111111",
17767=>"110111110",
17768=>"100000000",
17769=>"111001000",
17770=>"100010011",
17771=>"101111111",
17772=>"110001100",
17773=>"001100110",
17774=>"110000100",
17775=>"000110101",
17776=>"111101101",
17777=>"110110011",
17778=>"110110001",
17779=>"001001011",
17780=>"001011010",
17781=>"000000000",
17782=>"000100111",
17783=>"000111011",
17784=>"111001010",
17785=>"110111011",
17786=>"010011001",
17787=>"001000000",
17788=>"111100111",
17789=>"000000000",
17790=>"111001100",
17791=>"101100110",
17792=>"011001011",
17793=>"000000000",
17794=>"101011011",
17795=>"100110011",
17796=>"011001001",
17797=>"100001101",
17798=>"001001001",
17799=>"110100000",
17800=>"000011111",
17801=>"000001000",
17802=>"110000001",
17803=>"100000000",
17804=>"110110010",
17805=>"111001100",
17806=>"111100110",
17807=>"000001010",
17808=>"111100111",
17809=>"100100110",
17810=>"000000001",
17811=>"110110111",
17812=>"000000001",
17813=>"011110110",
17814=>"110111010",
17815=>"100000000",
17816=>"100011011",
17817=>"000000111",
17818=>"000010100",
17819=>"011000101",
17820=>"100110011",
17821=>"100100000",
17822=>"111111110",
17823=>"000100100",
17824=>"111111000",
17825=>"011000100",
17826=>"000000000",
17827=>"100100000",
17828=>"110011001",
17829=>"000001111",
17830=>"001001100",
17831=>"110001001",
17832=>"001001010",
17833=>"101100100",
17834=>"011101110",
17835=>"000000100",
17836=>"100101100",
17837=>"111001000",
17838=>"000000000",
17839=>"100100110",
17840=>"000000000",
17841=>"111111111",
17842=>"010010000",
17843=>"111111111",
17844=>"110000000",
17845=>"010010000",
17846=>"100110000",
17847=>"011111101",
17848=>"100101000",
17849=>"100110010",
17850=>"110101110",
17851=>"010011011",
17852=>"101001001",
17853=>"110110001",
17854=>"101100011",
17855=>"000000011",
17856=>"010000000",
17857=>"100111000",
17858=>"110111111",
17859=>"011111111",
17860=>"000000000",
17861=>"010111110",
17862=>"100000000",
17863=>"000010010",
17864=>"000000000",
17865=>"000000000",
17866=>"010001110",
17867=>"100110111",
17868=>"110110111",
17869=>"000000000",
17870=>"001101111",
17871=>"000000100",
17872=>"100110010",
17873=>"011110111",
17874=>"100000000",
17875=>"110011011",
17876=>"011001100",
17877=>"011010000",
17878=>"011011110",
17879=>"000000000",
17880=>"110011001",
17881=>"000000101",
17882=>"001111111",
17883=>"011100110",
17884=>"000000000",
17885=>"000000000",
17886=>"100111000",
17887=>"100010011",
17888=>"000000100",
17889=>"001000100",
17890=>"110011001",
17891=>"111011101",
17892=>"000000001",
17893=>"011110011",
17894=>"100011111",
17895=>"111011111",
17896=>"000001011",
17897=>"000000000",
17898=>"000100011",
17899=>"100101110",
17900=>"100100111",
17901=>"011000100",
17902=>"110000000",
17903=>"001000011",
17904=>"000001011",
17905=>"000000000",
17906=>"111001011",
17907=>"000011001",
17908=>"000000000",
17909=>"001000100",
17910=>"001100011",
17911=>"111000000",
17912=>"010010001",
17913=>"010000111",
17914=>"101110101",
17915=>"001111011",
17916=>"111011011",
17917=>"001001001",
17918=>"000100000",
17919=>"111011001",
17920=>"111011000",
17921=>"100110010",
17922=>"110110110",
17923=>"000111001",
17924=>"110011011",
17925=>"100000111",
17926=>"100100000",
17927=>"100111110",
17928=>"011001001",
17929=>"111110001",
17930=>"101100000",
17931=>"111000000",
17932=>"000000000",
17933=>"000000000",
17934=>"110111110",
17935=>"000001011",
17936=>"111111001",
17937=>"011000000",
17938=>"111111101",
17939=>"100101000",
17940=>"111111100",
17941=>"111111111",
17942=>"111111001",
17943=>"111111000",
17944=>"111111111",
17945=>"001000011",
17946=>"000100000",
17947=>"111000000",
17948=>"001000000",
17949=>"000000010",
17950=>"101001110",
17951=>"010000001",
17952=>"100000000",
17953=>"010000000",
17954=>"010000100",
17955=>"000001111",
17956=>"100100000",
17957=>"101010001",
17958=>"111111011",
17959=>"111011101",
17960=>"111111000",
17961=>"000000000",
17962=>"110111111",
17963=>"110000010",
17964=>"110100000",
17965=>"111111001",
17966=>"000000101",
17967=>"111011111",
17968=>"111111111",
17969=>"011000111",
17970=>"000000010",
17971=>"000000111",
17972=>"111010000",
17973=>"111011101",
17974=>"011011000",
17975=>"000000000",
17976=>"111010000",
17977=>"111111000",
17978=>"000000001",
17979=>"111000011",
17980=>"000110000",
17981=>"001001001",
17982=>"100111000",
17983=>"111111101",
17984=>"110000000",
17985=>"011000001",
17986=>"000111100",
17987=>"111111011",
17988=>"000011001",
17989=>"000000111",
17990=>"000100100",
17991=>"001000011",
17992=>"000000000",
17993=>"011111000",
17994=>"111100101",
17995=>"000010111",
17996=>"001000011",
17997=>"110000001",
17998=>"010111001",
17999=>"000000111",
18000=>"000101101",
18001=>"000111001",
18002=>"010111111",
18003=>"101000000",
18004=>"111111011",
18005=>"110111001",
18006=>"010110011",
18007=>"111001001",
18008=>"110110000",
18009=>"001001011",
18010=>"001111110",
18011=>"011100100",
18012=>"111111000",
18013=>"001010000",
18014=>"110100111",
18015=>"111111000",
18016=>"100100000",
18017=>"111111111",
18018=>"001100111",
18019=>"110111001",
18020=>"010011000",
18021=>"000100111",
18022=>"111001111",
18023=>"000000111",
18024=>"111111000",
18025=>"000000000",
18026=>"110101101",
18027=>"000000011",
18028=>"000100000",
18029=>"000011111",
18030=>"111010110",
18031=>"000011000",
18032=>"100100011",
18033=>"000110111",
18034=>"111100000",
18035=>"000000111",
18036=>"100001101",
18037=>"101010011",
18038=>"110011000",
18039=>"000110110",
18040=>"011111010",
18041=>"000000000",
18042=>"010001100",
18043=>"111000000",
18044=>"111000000",
18045=>"000000101",
18046=>"001100000",
18047=>"111101000",
18048=>"111011010",
18049=>"001000000",
18050=>"111111100",
18051=>"000000010",
18052=>"000000000",
18053=>"111111001",
18054=>"101100000",
18055=>"000100000",
18056=>"000110010",
18057=>"111111000",
18058=>"001101111",
18059=>"000000111",
18060=>"001111111",
18061=>"111101001",
18062=>"111111100",
18063=>"000010000",
18064=>"001001110",
18065=>"111111000",
18066=>"000010000",
18067=>"110111000",
18068=>"111111100",
18069=>"000101000",
18070=>"000110110",
18071=>"010100101",
18072=>"111100101",
18073=>"011111010",
18074=>"111110100",
18075=>"111101100",
18076=>"111111111",
18077=>"111100000",
18078=>"111110101",
18079=>"000000110",
18080=>"111100100",
18081=>"111111111",
18082=>"000101110",
18083=>"110000111",
18084=>"111000000",
18085=>"100110000",
18086=>"001001111",
18087=>"111111101",
18088=>"101111100",
18089=>"111110111",
18090=>"111000111",
18091=>"000111111",
18092=>"000001100",
18093=>"000000011",
18094=>"111110000",
18095=>"000000111",
18096=>"100000000",
18097=>"000000000",
18098=>"000110000",
18099=>"010100000",
18100=>"001110000",
18101=>"111101001",
18102=>"010010010",
18103=>"000000111",
18104=>"010001000",
18105=>"111111101",
18106=>"111101111",
18107=>"100000111",
18108=>"000000101",
18109=>"011111111",
18110=>"110110000",
18111=>"000000100",
18112=>"111110000",
18113=>"000000110",
18114=>"000011110",
18115=>"111110111",
18116=>"000000100",
18117=>"101011011",
18118=>"011011110",
18119=>"101000000",
18120=>"100000000",
18121=>"111001011",
18122=>"000001011",
18123=>"111000000",
18124=>"111011111",
18125=>"110011000",
18126=>"000010110",
18127=>"101000000",
18128=>"111100100",
18129=>"000000010",
18130=>"000001010",
18131=>"010010111",
18132=>"111000000",
18133=>"100010011",
18134=>"111000000",
18135=>"111011000",
18136=>"111111000",
18137=>"011111001",
18138=>"111001010",
18139=>"000000111",
18140=>"001111100",
18141=>"000101111",
18142=>"001011111",
18143=>"101110000",
18144=>"111111111",
18145=>"100000111",
18146=>"110000100",
18147=>"010110000",
18148=>"000000010",
18149=>"111000000",
18150=>"110011000",
18151=>"110100110",
18152=>"000000011",
18153=>"000000001",
18154=>"111001000",
18155=>"000000101",
18156=>"111111111",
18157=>"000000011",
18158=>"000000011",
18159=>"111000000",
18160=>"100011000",
18161=>"011111100",
18162=>"111101101",
18163=>"100110000",
18164=>"001000000",
18165=>"000111111",
18166=>"000000111",
18167=>"111101111",
18168=>"111101000",
18169=>"111101111",
18170=>"000011011",
18171=>"010001000",
18172=>"111111000",
18173=>"101101111",
18174=>"001000110",
18175=>"000000000",
18176=>"000000111",
18177=>"000011000",
18178=>"000001001",
18179=>"110000000",
18180=>"010011001",
18181=>"100000000",
18182=>"111111111",
18183=>"000011001",
18184=>"100000000",
18185=>"111111001",
18186=>"000111001",
18187=>"100000000",
18188=>"111000000",
18189=>"000111111",
18190=>"001110100",
18191=>"000000000",
18192=>"111101001",
18193=>"101111000",
18194=>"111111110",
18195=>"110010000",
18196=>"000000000",
18197=>"111111111",
18198=>"000011110",
18199=>"111011111",
18200=>"111111111",
18201=>"000000000",
18202=>"000011000",
18203=>"111111000",
18204=>"000000010",
18205=>"000000000",
18206=>"111101111",
18207=>"011000000",
18208=>"000000000",
18209=>"000111000",
18210=>"000100000",
18211=>"111000100",
18212=>"111111111",
18213=>"111001110",
18214=>"111111111",
18215=>"111111111",
18216=>"111111000",
18217=>"111111001",
18218=>"000110000",
18219=>"000011010",
18220=>"110100110",
18221=>"111010111",
18222=>"000011100",
18223=>"000010000",
18224=>"111111110",
18225=>"111011011",
18226=>"111111100",
18227=>"000111000",
18228=>"110010101",
18229=>"111111110",
18230=>"001011101",
18231=>"000001000",
18232=>"010000011",
18233=>"000110000",
18234=>"110100111",
18235=>"100110000",
18236=>"100111011",
18237=>"001111111",
18238=>"000100000",
18239=>"011011011",
18240=>"000010001",
18241=>"001111111",
18242=>"000000000",
18243=>"100000100",
18244=>"110110000",
18245=>"111101110",
18246=>"111111111",
18247=>"111111101",
18248=>"000000010",
18249=>"001000000",
18250=>"100101110",
18251=>"000111111",
18252=>"111011000",
18253=>"110000000",
18254=>"001000010",
18255=>"111000101",
18256=>"111001000",
18257=>"010111010",
18258=>"000010000",
18259=>"011111001",
18260=>"000000000",
18261=>"110110111",
18262=>"110010010",
18263=>"001001000",
18264=>"001000101",
18265=>"000010011",
18266=>"110110001",
18267=>"111111111",
18268=>"000000000",
18269=>"000111110",
18270=>"010110000",
18271=>"011100000",
18272=>"101101000",
18273=>"000110010",
18274=>"000001000",
18275=>"101111111",
18276=>"111111111",
18277=>"000000000",
18278=>"000000000",
18279=>"000000010",
18280=>"010110100",
18281=>"000100111",
18282=>"000000001",
18283=>"010111111",
18284=>"000000000",
18285=>"111010000",
18286=>"111111011",
18287=>"111111111",
18288=>"011011110",
18289=>"000000100",
18290=>"000110110",
18291=>"000000000",
18292=>"000010000",
18293=>"110000111",
18294=>"100110100",
18295=>"000000011",
18296=>"100101000",
18297=>"110111110",
18298=>"111111111",
18299=>"111000001",
18300=>"001011001",
18301=>"001011011",
18302=>"010111111",
18303=>"000000010",
18304=>"000000000",
18305=>"000111111",
18306=>"010011011",
18307=>"011101111",
18308=>"111011001",
18309=>"111101111",
18310=>"110100110",
18311=>"110101000",
18312=>"111111111",
18313=>"000101000",
18314=>"111110111",
18315=>"111101001",
18316=>"000010000",
18317=>"000011110",
18318=>"000000000",
18319=>"000000000",
18320=>"110111011",
18321=>"010111111",
18322=>"000001001",
18323=>"111101101",
18324=>"000001001",
18325=>"100101100",
18326=>"000000000",
18327=>"100111110",
18328=>"111000000",
18329=>"000001001",
18330=>"111111111",
18331=>"101011000",
18332=>"000000000",
18333=>"111000010",
18334=>"001111110",
18335=>"011010000",
18336=>"111111111",
18337=>"001011010",
18338=>"011111110",
18339=>"000001111",
18340=>"000111111",
18341=>"110100100",
18342=>"111101010",
18343=>"111000000",
18344=>"101000111",
18345=>"000101010",
18346=>"010110000",
18347=>"011011000",
18348=>"111001111",
18349=>"000001111",
18350=>"100011000",
18351=>"000111011",
18352=>"010000001",
18353=>"001100000",
18354=>"000000000",
18355=>"000011001",
18356=>"011000111",
18357=>"111111110",
18358=>"000001001",
18359=>"010000000",
18360=>"001110000",
18361=>"100111101",
18362=>"111010001",
18363=>"010001110",
18364=>"110110111",
18365=>"011111010",
18366=>"000000000",
18367=>"000111011",
18368=>"000111111",
18369=>"000000000",
18370=>"111111101",
18371=>"011011011",
18372=>"000100100",
18373=>"000110110",
18374=>"000010000",
18375=>"000101000",
18376=>"111110010",
18377=>"101101111",
18378=>"101100101",
18379=>"111111111",
18380=>"010010010",
18381=>"000101100",
18382=>"110111010",
18383=>"111111111",
18384=>"010010010",
18385=>"111111111",
18386=>"100010000",
18387=>"000000000",
18388=>"000000000",
18389=>"000000000",
18390=>"111111000",
18391=>"010111000",
18392=>"000000010",
18393=>"010010000",
18394=>"111111111",
18395=>"010111000",
18396=>"110111110",
18397=>"000001101",
18398=>"000000100",
18399=>"000000011",
18400=>"000000000",
18401=>"010010001",
18402=>"010000111",
18403=>"000000011",
18404=>"000000000",
18405=>"000010010",
18406=>"011111111",
18407=>"000111101",
18408=>"111000001",
18409=>"110110001",
18410=>"011111000",
18411=>"001001000",
18412=>"001000000",
18413=>"101101100",
18414=>"000011000",
18415=>"000000000",
18416=>"000000000",
18417=>"011011111",
18418=>"111101111",
18419=>"110110000",
18420=>"010000111",
18421=>"110010010",
18422=>"111000111",
18423=>"000010000",
18424=>"000010011",
18425=>"111101010",
18426=>"111001000",
18427=>"000010000",
18428=>"111111111",
18429=>"000011000",
18430=>"111111011",
18431=>"101111000",
18432=>"101111001",
18433=>"111011011",
18434=>"111000001",
18435=>"000000110",
18436=>"010011111",
18437=>"010100001",
18438=>"011001001",
18439=>"110111010",
18440=>"111011011",
18441=>"001111001",
18442=>"000000001",
18443=>"011001001",
18444=>"000100100",
18445=>"100100000",
18446=>"001101110",
18447=>"000010000",
18448=>"001111001",
18449=>"000000110",
18450=>"010000000",
18451=>"001000100",
18452=>"111100100",
18453=>"011000000",
18454=>"001001011",
18455=>"100001111",
18456=>"011001011",
18457=>"111011001",
18458=>"100110001",
18459=>"000000110",
18460=>"001011111",
18461=>"000000110",
18462=>"110100010",
18463=>"110100000",
18464=>"001001001",
18465=>"101110001",
18466=>"000111111",
18467=>"010000011",
18468=>"111111101",
18469=>"011010111",
18470=>"001011001",
18471=>"000110110",
18472=>"100110000",
18473=>"100100000",
18474=>"001001001",
18475=>"110011011",
18476=>"001111111",
18477=>"110010001",
18478=>"001101101",
18479=>"110111110",
18480=>"000101110",
18481=>"011111111",
18482=>"111101101",
18483=>"110110101",
18484=>"000100111",
18485=>"001000101",
18486=>"001010000",
18487=>"011001011",
18488=>"100000000",
18489=>"011001011",
18490=>"000101110",
18491=>"001011100",
18492=>"110111111",
18493=>"100011011",
18494=>"011001001",
18495=>"111101111",
18496=>"001000000",
18497=>"001111011",
18498=>"001000001",
18499=>"001011011",
18500=>"100000110",
18501=>"011000001",
18502=>"100001011",
18503=>"110010000",
18504=>"010111111",
18505=>"111110110",
18506=>"011001011",
18507=>"011001011",
18508=>"011001001",
18509=>"001111100",
18510=>"010000000",
18511=>"110010111",
18512=>"001110100",
18513=>"110101000",
18514=>"011001000",
18515=>"110011001",
18516=>"010000110",
18517=>"111010111",
18518=>"111111011",
18519=>"011111111",
18520=>"110001101",
18521=>"001101010",
18522=>"100001011",
18523=>"000000110",
18524=>"001000010",
18525=>"100100000",
18526=>"000110110",
18527=>"011001011",
18528=>"011001111",
18529=>"100010011",
18530=>"100000001",
18531=>"110101000",
18532=>"111100100",
18533=>"011001001",
18534=>"000110110",
18535=>"011011010",
18536=>"011000110",
18537=>"110100001",
18538=>"110110100",
18539=>"110111001",
18540=>"001011001",
18541=>"111100100",
18542=>"001001001",
18543=>"001110110",
18544=>"100000000",
18545=>"010001100",
18546=>"100111011",
18547=>"001001010",
18548=>"000101110",
18549=>"011001011",
18550=>"100100100",
18551=>"100110100",
18552=>"110010000",
18553=>"110110010",
18554=>"100000001",
18555=>"110111000",
18556=>"000100011",
18557=>"110000000",
18558=>"101001011",
18559=>"100000000",
18560=>"001011111",
18561=>"010000000",
18562=>"111001111",
18563=>"100111111",
18564=>"100110000",
18565=>"011000110",
18566=>"001011110",
18567=>"011001001",
18568=>"110111111",
18569=>"010000110",
18570=>"111011011",
18571=>"011011001",
18572=>"011000000",
18573=>"001000001",
18574=>"011001000",
18575=>"010001001",
18576=>"001001001",
18577=>"001111010",
18578=>"001001000",
18579=>"111011001",
18580=>"001001001",
18581=>"111100001",
18582=>"011011011",
18583=>"111111101",
18584=>"011100001",
18585=>"010100111",
18586=>"101001000",
18587=>"000000000",
18588=>"111010000",
18589=>"111011101",
18590=>"000000111",
18591=>"011001011",
18592=>"001111111",
18593=>"011111000",
18594=>"000001001",
18595=>"000001001",
18596=>"100100110",
18597=>"000001011",
18598=>"110100110",
18599=>"100110100",
18600=>"111000001",
18601=>"010100100",
18602=>"100100000",
18603=>"101100000",
18604=>"101100100",
18605=>"001100100",
18606=>"110001110",
18607=>"111110110",
18608=>"011001011",
18609=>"110110011",
18610=>"110001111",
18611=>"110101000",
18612=>"111111101",
18613=>"111011010",
18614=>"111111001",
18615=>"101111110",
18616=>"000100111",
18617=>"000100011",
18618=>"010011100",
18619=>"001100100",
18620=>"011011010",
18621=>"110110110",
18622=>"100111111",
18623=>"000001111",
18624=>"011001001",
18625=>"000001001",
18626=>"000100110",
18627=>"100111111",
18628=>"011001001",
18629=>"101100001",
18630=>"110100100",
18631=>"110110001",
18632=>"100001101",
18633=>"011001011",
18634=>"000011001",
18635=>"011011111",
18636=>"111001001",
18637=>"111111001",
18638=>"011001011",
18639=>"010001001",
18640=>"111001000",
18641=>"000000000",
18642=>"000000000",
18643=>"100000000",
18644=>"011001011",
18645=>"110011001",
18646=>"001011000",
18647=>"001011111",
18648=>"011011111",
18649=>"100100110",
18650=>"000010100",
18651=>"111001001",
18652=>"001111000",
18653=>"000110110",
18654=>"011010010",
18655=>"100000000",
18656=>"011010101",
18657=>"101110110",
18658=>"111110100",
18659=>"011011101",
18660=>"111001001",
18661=>"000001111",
18662=>"111001101",
18663=>"000011111",
18664=>"100100101",
18665=>"000100000",
18666=>"000000101",
18667=>"000010101",
18668=>"110110100",
18669=>"011001000",
18670=>"100100100",
18671=>"000000001",
18672=>"011001011",
18673=>"011010011",
18674=>"011111111",
18675=>"000000110",
18676=>"011100101",
18677=>"100001000",
18678=>"001001001",
18679=>"100011110",
18680=>"000101010",
18681=>"100001100",
18682=>"101001001",
18683=>"000010010",
18684=>"011001001",
18685=>"010000000",
18686=>"111001001",
18687=>"010001001",
18688=>"000000100",
18689=>"101000000",
18690=>"010110110",
18691=>"101000000",
18692=>"110100110",
18693=>"111100111",
18694=>"111001000",
18695=>"100111111",
18696=>"000000000",
18697=>"001111001",
18698=>"000000000",
18699=>"101000000",
18700=>"100110111",
18701=>"000000000",
18702=>"000000000",
18703=>"011111000",
18704=>"100000000",
18705=>"000000000",
18706=>"000001000",
18707=>"000101101",
18708=>"111111000",
18709=>"000011010",
18710=>"111111111",
18711=>"111111111",
18712=>"000000000",
18713=>"000000000",
18714=>"111100101",
18715=>"000011000",
18716=>"101000000",
18717=>"000000000",
18718=>"000100111",
18719=>"111111111",
18720=>"010111111",
18721=>"101000100",
18722=>"101000000",
18723=>"101111101",
18724=>"110111100",
18725=>"000000101",
18726=>"000000000",
18727=>"100000000",
18728=>"011111011",
18729=>"111111111",
18730=>"000000110",
18731=>"111100001",
18732=>"110010010",
18733=>"000000000",
18734=>"000100000",
18735=>"001111111",
18736=>"111101101",
18737=>"110100110",
18738=>"101000101",
18739=>"000000111",
18740=>"000000000",
18741=>"100000000",
18742=>"001000000",
18743=>"011011111",
18744=>"011111001",
18745=>"000000000",
18746=>"000000111",
18747=>"111111111",
18748=>"100101000",
18749=>"101111111",
18750=>"000000000",
18751=>"011011111",
18752=>"111101111",
18753=>"010010111",
18754=>"101101100",
18755=>"111110111",
18756=>"000100100",
18757=>"000010111",
18758=>"101000000",
18759=>"100101101",
18760=>"000000010",
18761=>"000000000",
18762=>"000000000",
18763=>"000111111",
18764=>"010111011",
18765=>"011001100",
18766=>"100000111",
18767=>"000000111",
18768=>"100000000",
18769=>"011011111",
18770=>"000000000",
18771=>"100100100",
18772=>"111001101",
18773=>"111111111",
18774=>"010000000",
18775=>"101000000",
18776=>"000000000",
18777=>"000000000",
18778=>"111111111",
18779=>"101011110",
18780=>"000000000",
18781=>"010000100",
18782=>"010111111",
18783=>"100001001",
18784=>"101001000",
18785=>"111000000",
18786=>"000110000",
18787=>"110111101",
18788=>"001000000",
18789=>"000000000",
18790=>"000000000",
18791=>"011111111",
18792=>"010111011",
18793=>"000000000",
18794=>"100000111",
18795=>"000000000",
18796=>"011101111",
18797=>"000000000",
18798=>"111111010",
18799=>"010000000",
18800=>"011000000",
18801=>"100111110",
18802=>"001100000",
18803=>"000000000",
18804=>"000101100",
18805=>"000000000",
18806=>"000011010",
18807=>"010010111",
18808=>"111111111",
18809=>"101001000",
18810=>"001001001",
18811=>"111100100",
18812=>"011000100",
18813=>"010001101",
18814=>"000111111",
18815=>"100100000",
18816=>"000101100",
18817=>"111111111",
18818=>"110111000",
18819=>"000101000",
18820=>"000000111",
18821=>"000000001",
18822=>"000000001",
18823=>"000000000",
18824=>"001000001",
18825=>"000100100",
18826=>"000000000",
18827=>"000000110",
18828=>"011111011",
18829=>"101110000",
18830=>"010000000",
18831=>"111100100",
18832=>"000000000",
18833=>"111111111",
18834=>"111111111",
18835=>"100100101",
18836=>"000000000",
18837=>"000111010",
18838=>"111000000",
18839=>"110110110",
18840=>"001000001",
18841=>"000111101",
18842=>"000000011",
18843=>"111111001",
18844=>"000000000",
18845=>"111111100",
18846=>"000000101",
18847=>"010000010",
18848=>"111111111",
18849=>"111101100",
18850=>"000000000",
18851=>"100000000",
18852=>"000000010",
18853=>"000000000",
18854=>"001000001",
18855=>"101011100",
18856=>"100000000",
18857=>"101001000",
18858=>"001000111",
18859=>"110000000",
18860=>"111011111",
18861=>"000100000",
18862=>"011011110",
18863=>"001111001",
18864=>"111111111",
18865=>"100000000",
18866=>"010111111",
18867=>"001000001",
18868=>"110100000",
18869=>"000000111",
18870=>"111100000",
18871=>"100000100",
18872=>"001110100",
18873=>"000000000",
18874=>"000101000",
18875=>"111101000",
18876=>"000000000",
18877=>"010111111",
18878=>"110110110",
18879=>"110111111",
18880=>"000111001",
18881=>"001001000",
18882=>"000000000",
18883=>"111111011",
18884=>"000000000",
18885=>"001101111",
18886=>"111101100",
18887=>"000011111",
18888=>"100100001",
18889=>"111111111",
18890=>"000000000",
18891=>"000010010",
18892=>"000010010",
18893=>"010000000",
18894=>"111000110",
18895=>"001100000",
18896=>"000010011",
18897=>"111010001",
18898=>"000000000",
18899=>"000000000",
18900=>"000000111",
18901=>"111000000",
18902=>"011111000",
18903=>"000000000",
18904=>"011111111",
18905=>"011100111",
18906=>"111101101",
18907=>"000010000",
18908=>"011111111",
18909=>"101001100",
18910=>"000000000",
18911=>"001111011",
18912=>"000000111",
18913=>"100000101",
18914=>"100000000",
18915=>"111000000",
18916=>"110111000",
18917=>"111111011",
18918=>"111000000",
18919=>"100100110",
18920=>"100111111",
18921=>"111111111",
18922=>"100000000",
18923=>"100000100",
18924=>"101001000",
18925=>"111111110",
18926=>"110111000",
18927=>"010110000",
18928=>"000111011",
18929=>"010000110",
18930=>"111111111",
18931=>"000000000",
18932=>"000000000",
18933=>"001111000",
18934=>"000000000",
18935=>"000000001",
18936=>"000000000",
18937=>"111001000",
18938=>"100000000",
18939=>"000000000",
18940=>"111111110",
18941=>"100110100",
18942=>"100000110",
18943=>"000000100",
18944=>"011001000",
18945=>"000000100",
18946=>"101000101",
18947=>"000000001",
18948=>"000011011",
18949=>"010010111",
18950=>"010111010",
18951=>"000010000",
18952=>"000110000",
18953=>"101011000",
18954=>"000110010",
18955=>"000000100",
18956=>"000000000",
18957=>"010011000",
18958=>"000000110",
18959=>"010010000",
18960=>"110111000",
18961=>"110111001",
18962=>"000000100",
18963=>"000000010",
18964=>"000000100",
18965=>"111101111",
18966=>"000100101",
18967=>"101111010",
18968=>"101000000",
18969=>"111101101",
18970=>"000001101",
18971=>"000000001",
18972=>"100100100",
18973=>"111110000",
18974=>"111101111",
18975=>"000010010",
18976=>"010000101",
18977=>"101100101",
18978=>"000001111",
18979=>"000000000",
18980=>"001001001",
18981=>"011010110",
18982=>"001111111",
18983=>"000111111",
18984=>"111000000",
18985=>"011000000",
18986=>"000011000",
18987=>"001000000",
18988=>"010011011",
18989=>"111011110",
18990=>"011101100",
18991=>"100010110",
18992=>"000000110",
18993=>"011101000",
18994=>"101000000",
18995=>"111111000",
18996=>"000000000",
18997=>"000000100",
18998=>"000111110",
18999=>"000000000",
19000=>"111010000",
19001=>"000111110",
19002=>"010000000",
19003=>"111111111",
19004=>"001111110",
19005=>"111111110",
19006=>"000000000",
19007=>"110111100",
19008=>"001000100",
19009=>"100000111",
19010=>"000010010",
19011=>"110100001",
19012=>"111111111",
19013=>"000101111",
19014=>"000000000",
19015=>"100101000",
19016=>"000010011",
19017=>"001011111",
19018=>"111001100",
19019=>"000111111",
19020=>"100100100",
19021=>"110110100",
19022=>"100111111",
19023=>"110111010",
19024=>"111111101",
19025=>"111000010",
19026=>"000010111",
19027=>"111111001",
19028=>"000000000",
19029=>"000011011",
19030=>"000110110",
19031=>"001000000",
19032=>"100111111",
19033=>"000010011",
19034=>"000001100",
19035=>"101101111",
19036=>"001010000",
19037=>"000000010",
19038=>"010111111",
19039=>"010100110",
19040=>"101111111",
19041=>"001001000",
19042=>"111101101",
19043=>"000101000",
19044=>"000111010",
19045=>"000011001",
19046=>"000100101",
19047=>"100000000",
19048=>"000000111",
19049=>"111000011",
19050=>"011111000",
19051=>"000011011",
19052=>"000000111",
19053=>"010110000",
19054=>"101000000",
19055=>"010111111",
19056=>"100111101",
19057=>"010000010",
19058=>"111111011",
19059=>"011101000",
19060=>"111010000",
19061=>"000001000",
19062=>"000111111",
19063=>"010101011",
19064=>"001100011",
19065=>"010000000",
19066=>"110110111",
19067=>"111100111",
19068=>"110110010",
19069=>"111100000",
19070=>"101000001",
19071=>"001001101",
19072=>"111001101",
19073=>"110100000",
19074=>"011011111",
19075=>"010010011",
19076=>"111111101",
19077=>"111101000",
19078=>"110110001",
19079=>"010110010",
19080=>"110101100",
19081=>"000110101",
19082=>"010111000",
19083=>"110001100",
19084=>"101001101",
19085=>"001010010",
19086=>"000011110",
19087=>"000000000",
19088=>"001011001",
19089=>"100101100",
19090=>"000010000",
19091=>"001101000",
19092=>"000111111",
19093=>"000111001",
19094=>"000001111",
19095=>"000010000",
19096=>"000000000",
19097=>"001101101",
19098=>"000011011",
19099=>"111100000",
19100=>"000000000",
19101=>"111101111",
19102=>"011010000",
19103=>"000000100",
19104=>"001011111",
19105=>"111011111",
19106=>"111001000",
19107=>"000000001",
19108=>"000000011",
19109=>"000000000",
19110=>"100110110",
19111=>"000011010",
19112=>"011000111",
19113=>"111111111",
19114=>"000001101",
19115=>"010111111",
19116=>"111000000",
19117=>"011011011",
19118=>"100111111",
19119=>"010010000",
19120=>"000010000",
19121=>"010111000",
19122=>"000000010",
19123=>"110000010",
19124=>"000111000",
19125=>"100011010",
19126=>"000011111",
19127=>"110110010",
19128=>"000011011",
19129=>"000111111",
19130=>"000111110",
19131=>"000000000",
19132=>"110100111",
19133=>"111101111",
19134=>"011001111",
19135=>"011010010",
19136=>"001010000",
19137=>"101000000",
19138=>"011111000",
19139=>"000011000",
19140=>"000010000",
19141=>"111110000",
19142=>"000000111",
19143=>"011111000",
19144=>"111111111",
19145=>"000101001",
19146=>"110101101",
19147=>"101100111",
19148=>"000110000",
19149=>"100011111",
19150=>"010000101",
19151=>"111111111",
19152=>"111100101",
19153=>"110111001",
19154=>"000000111",
19155=>"100100100",
19156=>"000000001",
19157=>"110100000",
19158=>"000110000",
19159=>"010010000",
19160=>"100000000",
19161=>"000010010",
19162=>"001111011",
19163=>"111101000",
19164=>"000101110",
19165=>"001001000",
19166=>"000000000",
19167=>"000000111",
19168=>"000001001",
19169=>"011011101",
19170=>"000000000",
19171=>"000011000",
19172=>"010000000",
19173=>"101000011",
19174=>"000111111",
19175=>"000111011",
19176=>"100001111",
19177=>"010010110",
19178=>"000000100",
19179=>"111000101",
19180=>"111000000",
19181=>"000100000",
19182=>"100000000",
19183=>"111000000",
19184=>"010111111",
19185=>"100011001",
19186=>"111111011",
19187=>"000111010",
19188=>"000110001",
19189=>"101000000",
19190=>"000000000",
19191=>"000011111",
19192=>"000000100",
19193=>"110111111",
19194=>"110000000",
19195=>"101001111",
19196=>"111101111",
19197=>"000000000",
19198=>"000110000",
19199=>"111100000",
19200=>"001001100",
19201=>"001000010",
19202=>"111100101",
19203=>"000010100",
19204=>"000101111",
19205=>"000000111",
19206=>"001000111",
19207=>"000100111",
19208=>"011101000",
19209=>"111001000",
19210=>"001110110",
19211=>"111101110",
19212=>"111000000",
19213=>"001000000",
19214=>"001101101",
19215=>"001000000",
19216=>"000110101",
19217=>"000000000",
19218=>"110100000",
19219=>"100000000",
19220=>"111011100",
19221=>"010100111",
19222=>"001000000",
19223=>"111000000",
19224=>"000000001",
19225=>"111100000",
19226=>"000000010",
19227=>"100000111",
19228=>"000000000",
19229=>"111111111",
19230=>"010000101",
19231=>"000000001",
19232=>"011111011",
19233=>"111011010",
19234=>"000100010",
19235=>"011011101",
19236=>"110110000",
19237=>"110100100",
19238=>"010110110",
19239=>"000010101",
19240=>"010000000",
19241=>"000001111",
19242=>"111111101",
19243=>"010010010",
19244=>"111001101",
19245=>"111111000",
19246=>"010000111",
19247=>"111111001",
19248=>"000000101",
19249=>"000100110",
19250=>"000000010",
19251=>"000000111",
19252=>"010010010",
19253=>"011010010",
19254=>"101000000",
19255=>"011111111",
19256=>"110100001",
19257=>"101100101",
19258=>"010110100",
19259=>"001011010",
19260=>"000011101",
19261=>"111111010",
19262=>"000000000",
19263=>"110000001",
19264=>"111100001",
19265=>"110000100",
19266=>"100000010",
19267=>"001100111",
19268=>"001001000",
19269=>"010000000",
19270=>"000101111",
19271=>"010011111",
19272=>"100111111",
19273=>"010111000",
19274=>"101001111",
19275=>"111010011",
19276=>"111000000",
19277=>"001100100",
19278=>"001101001",
19279=>"000000011",
19280=>"000010011",
19281=>"111110101",
19282=>"101111111",
19283=>"011101100",
19284=>"000000000",
19285=>"110110100",
19286=>"010011000",
19287=>"000000111",
19288=>"000010010",
19289=>"100101100",
19290=>"000100011",
19291=>"111111011",
19292=>"111111010",
19293=>"000011011",
19294=>"111100100",
19295=>"000000111",
19296=>"000011010",
19297=>"000001011",
19298=>"101101101",
19299=>"000010110",
19300=>"001111101",
19301=>"101011100",
19302=>"000010011",
19303=>"000100000",
19304=>"010011111",
19305=>"000000000",
19306=>"111011101",
19307=>"000000111",
19308=>"000010010",
19309=>"000111111",
19310=>"011000000",
19311=>"001000000",
19312=>"111110001",
19313=>"011000101",
19314=>"101000001",
19315=>"010100000",
19316=>"000010011",
19317=>"101000000",
19318=>"000100001",
19319=>"010000001",
19320=>"111000010",
19321=>"000010011",
19322=>"110011101",
19323=>"111111010",
19324=>"011000000",
19325=>"100001110",
19326=>"010010010",
19327=>"000000011",
19328=>"111111101",
19329=>"010100111",
19330=>"000010010",
19331=>"010111111",
19332=>"100010011",
19333=>"111111010",
19334=>"011001001",
19335=>"101111111",
19336=>"001001100",
19337=>"001010010",
19338=>"111000001",
19339=>"000010000",
19340=>"000101010",
19341=>"000101100",
19342=>"101111100",
19343=>"000001000",
19344=>"100000001",
19345=>"000000100",
19346=>"101011010",
19347=>"000101111",
19348=>"000111011",
19349=>"101100100",
19350=>"100100110",
19351=>"010110100",
19352=>"000010111",
19353=>"000000100",
19354=>"010111000",
19355=>"011001010",
19356=>"100100100",
19357=>"000011011",
19358=>"011110111",
19359=>"101100110",
19360=>"101001000",
19361=>"010000111",
19362=>"100001111",
19363=>"000000000",
19364=>"010000100",
19365=>"110110010",
19366=>"110110001",
19367=>"000000010",
19368=>"010010010",
19369=>"101010000",
19370=>"000101100",
19371=>"000000101",
19372=>"011111001",
19373=>"100100100",
19374=>"000011111",
19375=>"011101110",
19376=>"000000000",
19377=>"000111011",
19378=>"100100000",
19379=>"000000001",
19380=>"001001010",
19381=>"100001010",
19382=>"111011000",
19383=>"011011101",
19384=>"100100001",
19385=>"010110110",
19386=>"110010010",
19387=>"011100110",
19388=>"010110110",
19389=>"010111011",
19390=>"011001000",
19391=>"011000101",
19392=>"110101000",
19393=>"011101011",
19394=>"011010001",
19395=>"000100000",
19396=>"011010000",
19397=>"011110000",
19398=>"011101000",
19399=>"011111010",
19400=>"110011000",
19401=>"111000000",
19402=>"011101000",
19403=>"110000100",
19404=>"100000001",
19405=>"111100000",
19406=>"000000000",
19407=>"111010100",
19408=>"111101101",
19409=>"000001111",
19410=>"100010111",
19411=>"011000011",
19412=>"100100000",
19413=>"000000110",
19414=>"101100111",
19415=>"001000111",
19416=>"000001001",
19417=>"100000000",
19418=>"111111010",
19419=>"000000000",
19420=>"001001000",
19421=>"111100011",
19422=>"000000011",
19423=>"011000000",
19424=>"101100010",
19425=>"101100100",
19426=>"001010111",
19427=>"000101111",
19428=>"000000001",
19429=>"101111111",
19430=>"000010111",
19431=>"000001111",
19432=>"111000011",
19433=>"000000011",
19434=>"110011111",
19435=>"111110000",
19436=>"111100000",
19437=>"011010000",
19438=>"110000000",
19439=>"001111111",
19440=>"001000010",
19441=>"111001001",
19442=>"111000000",
19443=>"100101110",
19444=>"011001001",
19445=>"000000111",
19446=>"000000011",
19447=>"001001100",
19448=>"111000000",
19449=>"110110010",
19450=>"101111101",
19451=>"000111111",
19452=>"000000000",
19453=>"011011111",
19454=>"001011000",
19455=>"111000111",
19456=>"000011100",
19457=>"000100111",
19458=>"101000100",
19459=>"101101100",
19460=>"101000011",
19461=>"110000100",
19462=>"000000000",
19463=>"000010111",
19464=>"001100000",
19465=>"101000100",
19466=>"101001001",
19467=>"000100100",
19468=>"111100100",
19469=>"111100000",
19470=>"100100000",
19471=>"010011111",
19472=>"100100100",
19473=>"001001000",
19474=>"010001011",
19475=>"000000000",
19476=>"111101000",
19477=>"111000000",
19478=>"010000101",
19479=>"000100000",
19480=>"100100010",
19481=>"001111111",
19482=>"101100000",
19483=>"000010000",
19484=>"000100000",
19485=>"011111011",
19486=>"111101100",
19487=>"001101101",
19488=>"101000000",
19489=>"101010001",
19490=>"100011000",
19491=>"000000100",
19492=>"101001000",
19493=>"001011110",
19494=>"111000000",
19495=>"100100000",
19496=>"101011011",
19497=>"001100000",
19498=>"110100100",
19499=>"010010011",
19500=>"111111011",
19501=>"101000100",
19502=>"111011111",
19503=>"000110100",
19504=>"000100111",
19505=>"000101011",
19506=>"101000000",
19507=>"000000111",
19508=>"000011100",
19509=>"000010111",
19510=>"000110110",
19511=>"111100100",
19512=>"011011110",
19513=>"101100100",
19514=>"101100100",
19515=>"000011010",
19516=>"011000011",
19517=>"111101110",
19518=>"000100000",
19519=>"110011011",
19520=>"000000000",
19521=>"010111011",
19522=>"011100000",
19523=>"111100100",
19524=>"111100101",
19525=>"111101100",
19526=>"001100100",
19527=>"010000111",
19528=>"010011100",
19529=>"111011000",
19530=>"000101101",
19531=>"101100100",
19532=>"010010100",
19533=>"000000110",
19534=>"101111111",
19535=>"110011010",
19536=>"111011011",
19537=>"111010111",
19538=>"110100100",
19539=>"011001000",
19540=>"100101111",
19541=>"010010010",
19542=>"111100111",
19543=>"101101101",
19544=>"000000000",
19545=>"110100000",
19546=>"001001000",
19547=>"100010011",
19548=>"100000100",
19549=>"001001001",
19550=>"100111111",
19551=>"100100100",
19552=>"111000000",
19553=>"111111101",
19554=>"101100100",
19555=>"110101100",
19556=>"000000010",
19557=>"000100100",
19558=>"000110001",
19559=>"010010100",
19560=>"111000000",
19561=>"111011101",
19562=>"111111101",
19563=>"011111010",
19564=>"100000111",
19565=>"000000010",
19566=>"101100100",
19567=>"000000011",
19568=>"100111111",
19569=>"100111101",
19570=>"000011001",
19571=>"000000000",
19572=>"111111111",
19573=>"000100100",
19574=>"100000111",
19575=>"000001000",
19576=>"111000000",
19577=>"010000000",
19578=>"100111011",
19579=>"111000000",
19580=>"000011011",
19581=>"111000000",
19582=>"011010000",
19583=>"101000000",
19584=>"000010110",
19585=>"000011000",
19586=>"000011001",
19587=>"000000000",
19588=>"111111111",
19589=>"111100000",
19590=>"010010011",
19591=>"100001110",
19592=>"100111111",
19593=>"011100010",
19594=>"100100111",
19595=>"111111101",
19596=>"100011011",
19597=>"000011011",
19598=>"010000000",
19599=>"010000000",
19600=>"001001001",
19601=>"000111011",
19602=>"000111011",
19603=>"100100010",
19604=>"000100111",
19605=>"111100100",
19606=>"111100111",
19607=>"100100100",
19608=>"001011111",
19609=>"000011011",
19610=>"101011011",
19611=>"010000000",
19612=>"011100100",
19613=>"000000001",
19614=>"000100100",
19615=>"111100111",
19616=>"000010011",
19617=>"001000010",
19618=>"000011011",
19619=>"011010000",
19620=>"000000001",
19621=>"001111110",
19622=>"001000101",
19623=>"000010011",
19624=>"000000100",
19625=>"111000101",
19626=>"001000000",
19627=>"111100100",
19628=>"100000000",
19629=>"101100101",
19630=>"011110101",
19631=>"000000011",
19632=>"101000001",
19633=>"001011000",
19634=>"010001011",
19635=>"001010011",
19636=>"110111011",
19637=>"000000000",
19638=>"000010011",
19639=>"110011110",
19640=>"010011010",
19641=>"000000011",
19642=>"000011011",
19643=>"111111011",
19644=>"111111111",
19645=>"111111111",
19646=>"101000000",
19647=>"010011111",
19648=>"000000000",
19649=>"110000000",
19650=>"010111011",
19651=>"001001001",
19652=>"111101000",
19653=>"001000010",
19654=>"000110111",
19655=>"111000100",
19656=>"111111110",
19657=>"000000000",
19658=>"001111111",
19659=>"111100100",
19660=>"100011001",
19661=>"000011111",
19662=>"010111111",
19663=>"000000001",
19664=>"011100000",
19665=>"101001101",
19666=>"000010011",
19667=>"111110110",
19668=>"101011000",
19669=>"100100111",
19670=>"111100100",
19671=>"000100100",
19672=>"000010010",
19673=>"000100111",
19674=>"101000011",
19675=>"100000000",
19676=>"111110011",
19677=>"111111000",
19678=>"100111000",
19679=>"100100111",
19680=>"111100001",
19681=>"101100100",
19682=>"100000000",
19683=>"111100101",
19684=>"100000000",
19685=>"110111111",
19686=>"000000011",
19687=>"010000110",
19688=>"010000000",
19689=>"011111111",
19690=>"110000000",
19691=>"111100100",
19692=>"000011011",
19693=>"111100100",
19694=>"001001001",
19695=>"000000111",
19696=>"000000000",
19697=>"100110111",
19698=>"010000000",
19699=>"011101010",
19700=>"101000001",
19701=>"011000011",
19702=>"000000000",
19703=>"010011011",
19704=>"000010000",
19705=>"010010100",
19706=>"111000001",
19707=>"000101101",
19708=>"111100100",
19709=>"000011011",
19710=>"011111111",
19711=>"000000001",
19712=>"011001100",
19713=>"000000100",
19714=>"000010000",
19715=>"101101100",
19716=>"111100001",
19717=>"001001000",
19718=>"010101101",
19719=>"111000101",
19720=>"111100101",
19721=>"000001000",
19722=>"000010110",
19723=>"111000110",
19724=>"000100100",
19725=>"111111111",
19726=>"100000001",
19727=>"001101001",
19728=>"000000010",
19729=>"000000111",
19730=>"000000000",
19731=>"000100111",
19732=>"001110010",
19733=>"000110111",
19734=>"011000010",
19735=>"001111110",
19736=>"000000000",
19737=>"000001111",
19738=>"001000100",
19739=>"000011000",
19740=>"111111111",
19741=>"111000000",
19742=>"111111010",
19743=>"000101101",
19744=>"000000110",
19745=>"001101100",
19746=>"000111100",
19747=>"011101111",
19748=>"100100010",
19749=>"110111111",
19750=>"000000111",
19751=>"000010111",
19752=>"111010111",
19753=>"111111111",
19754=>"000111011",
19755=>"100111000",
19756=>"110011011",
19757=>"011111011",
19758=>"111101000",
19759=>"000000000",
19760=>"011111000",
19761=>"011110100",
19762=>"111000000",
19763=>"111011010",
19764=>"000001011",
19765=>"101111111",
19766=>"000100111",
19767=>"000111000",
19768=>"111111000",
19769=>"011111001",
19770=>"111000000",
19771=>"111111000",
19772=>"001101011",
19773=>"010010111",
19774=>"000010010",
19775=>"000001011",
19776=>"111101101",
19777=>"101101001",
19778=>"001111000",
19779=>"000100110",
19780=>"110000000",
19781=>"111000000",
19782=>"000011110",
19783=>"010100000",
19784=>"111100001",
19785=>"111001001",
19786=>"010000101",
19787=>"000010110",
19788=>"000100101",
19789=>"011000111",
19790=>"110001000",
19791=>"100110100",
19792=>"000000111",
19793=>"111100000",
19794=>"100110111",
19795=>"001000110",
19796=>"101100010",
19797=>"101111100",
19798=>"100101111",
19799=>"000010000",
19800=>"111000111",
19801=>"110011111",
19802=>"001100110",
19803=>"000110111",
19804=>"000101111",
19805=>"011000000",
19806=>"010111111",
19807=>"000001011",
19808=>"100000000",
19809=>"000010010",
19810=>"100111011",
19811=>"000000111",
19812=>"010000000",
19813=>"111011101",
19814=>"010101101",
19815=>"000000100",
19816=>"010000000",
19817=>"011111000",
19818=>"011100010",
19819=>"001000101",
19820=>"011011001",
19821=>"010010111",
19822=>"000000000",
19823=>"011001001",
19824=>"110101101",
19825=>"111111000",
19826=>"000001111",
19827=>"111000110",
19828=>"000000101",
19829=>"100000101",
19830=>"001000110",
19831=>"000111111",
19832=>"000010010",
19833=>"000111111",
19834=>"010010101",
19835=>"011010000",
19836=>"110000000",
19837=>"100100001",
19838=>"111111011",
19839=>"000000011",
19840=>"101001011",
19841=>"110000001",
19842=>"111111001",
19843=>"110111000",
19844=>"011001101",
19845=>"000000001",
19846=>"111101100",
19847=>"000000110",
19848=>"001100000",
19849=>"010000000",
19850=>"111000011",
19851=>"100100110",
19852=>"110111000",
19853=>"010111111",
19854=>"000111101",
19855=>"000001001",
19856=>"111100110",
19857=>"100000100",
19858=>"000101111",
19859=>"111000010",
19860=>"000000000",
19861=>"001000000",
19862=>"000110000",
19863=>"011000100",
19864=>"000111111",
19865=>"111010010",
19866=>"000011000",
19867=>"000011111",
19868=>"111000000",
19869=>"000111111",
19870=>"000111000",
19871=>"000000000",
19872=>"100111011",
19873=>"011110010",
19874=>"100111000",
19875=>"100000111",
19876=>"111111101",
19877=>"000000011",
19878=>"011000001",
19879=>"000111000",
19880=>"011010000",
19881=>"000000111",
19882=>"111001111",
19883=>"000000111",
19884=>"100111000",
19885=>"000111011",
19886=>"011101101",
19887=>"011010111",
19888=>"100000000",
19889=>"011010111",
19890=>"000000000",
19891=>"000001001",
19892=>"110100100",
19893=>"100011000",
19894=>"100000110",
19895=>"011000100",
19896=>"101110110",
19897=>"010100010",
19898=>"101111011",
19899=>"101001000",
19900=>"110110011",
19901=>"000000111",
19902=>"011000100",
19903=>"111000000",
19904=>"000000110",
19905=>"000000010",
19906=>"101001100",
19907=>"011000000",
19908=>"001010000",
19909=>"100011001",
19910=>"111101000",
19911=>"000011110",
19912=>"000000110",
19913=>"000100100",
19914=>"010110010",
19915=>"000101101",
19916=>"010000011",
19917=>"011000110",
19918=>"000000010",
19919=>"111111000",
19920=>"011000010",
19921=>"010001011",
19922=>"011111101",
19923=>"101101111",
19924=>"000111111",
19925=>"000000111",
19926=>"000100111",
19927=>"000111110",
19928=>"111000000",
19929=>"111111111",
19930=>"111011110",
19931=>"000000010",
19932=>"101001000",
19933=>"000000100",
19934=>"100100010",
19935=>"110101000",
19936=>"111000000",
19937=>"111000010",
19938=>"111111011",
19939=>"001000111",
19940=>"000000111",
19941=>"101101101",
19942=>"001000111",
19943=>"110001111",
19944=>"010111111",
19945=>"000110000",
19946=>"000011011",
19947=>"001001111",
19948=>"000111100",
19949=>"000000101",
19950=>"000000000",
19951=>"111010110",
19952=>"011100100",
19953=>"000111000",
19954=>"111111000",
19955=>"100011001",
19956=>"100100010",
19957=>"000000001",
19958=>"000000111",
19959=>"011011000",
19960=>"111111000",
19961=>"010000000",
19962=>"111011111",
19963=>"010000001",
19964=>"100111111",
19965=>"000000111",
19966=>"011100100",
19967=>"100111110",
19968=>"000000100",
19969=>"110110111",
19970=>"000110111",
19971=>"110000100",
19972=>"110111111",
19973=>"001101000",
19974=>"011111111",
19975=>"110110101",
19976=>"000001011",
19977=>"111000111",
19978=>"000010000",
19979=>"000000000",
19980=>"001001111",
19981=>"111001101",
19982=>"000000000",
19983=>"001001010",
19984=>"111000000",
19985=>"001001011",
19986=>"000111111",
19987=>"011001001",
19988=>"111011000",
19989=>"000100100",
19990=>"011111011",
19991=>"000000001",
19992=>"000101111",
19993=>"000001101",
19994=>"001101001",
19995=>"111111111",
19996=>"110111111",
19997=>"000000000",
19998=>"000000000",
19999=>"110111000",
20000=>"000001000",
20001=>"000001010",
20002=>"101111111",
20003=>"110011001",
20004=>"100100100",
20005=>"011000011",
20006=>"110111001",
20007=>"111001000",
20008=>"010000010",
20009=>"000000001",
20010=>"110001000",
20011=>"111000000",
20012=>"001111101",
20013=>"010000000",
20014=>"101111001",
20015=>"111111000",
20016=>"000001000",
20017=>"001000000",
20018=>"000111110",
20019=>"111000010",
20020=>"101000010",
20021=>"111011000",
20022=>"000000010",
20023=>"101000000",
20024=>"000000111",
20025=>"111001100",
20026=>"100001010",
20027=>"000000111",
20028=>"011110100",
20029=>"010010111",
20030=>"000000000",
20031=>"100000000",
20032=>"000100111",
20033=>"000000100",
20034=>"111000001",
20035=>"001001000",
20036=>"111000000",
20037=>"010000100",
20038=>"000001011",
20039=>"000000000",
20040=>"111111111",
20041=>"110111110",
20042=>"101001111",
20043=>"000101001",
20044=>"000000101",
20045=>"011001111",
20046=>"110001001",
20047=>"110000001",
20048=>"000000000",
20049=>"000111111",
20050=>"000001001",
20051=>"001000000",
20052=>"010010000",
20053=>"110111110",
20054=>"000011010",
20055=>"100000111",
20056=>"000110111",
20057=>"110000011",
20058=>"111011000",
20059=>"000000000",
20060=>"110000001",
20061=>"111110100",
20062=>"110111111",
20063=>"001110110",
20064=>"000111111",
20065=>"010000000",
20066=>"001001111",
20067=>"101111001",
20068=>"001001001",
20069=>"000110010",
20070=>"001001110",
20071=>"110001001",
20072=>"110111100",
20073=>"000111110",
20074=>"111100011",
20075=>"100000000",
20076=>"111111110",
20077=>"111111001",
20078=>"110001011",
20079=>"001100101",
20080=>"000000001",
20081=>"010000000",
20082=>"011001000",
20083=>"111000000",
20084=>"101001001",
20085=>"000101111",
20086=>"001011100",
20087=>"000001001",
20088=>"101111000",
20089=>"111110111",
20090=>"000001001",
20091=>"000010111",
20092=>"011011110",
20093=>"100000000",
20094=>"110010110",
20095=>"001111111",
20096=>"010001001",
20097=>"001110010",
20098=>"001001001",
20099=>"111110100",
20100=>"101001000",
20101=>"001110111",
20102=>"000000100",
20103=>"011001101",
20104=>"001001111",
20105=>"000000001",
20106=>"101011001",
20107=>"010000000",
20108=>"111111000",
20109=>"000101111",
20110=>"000100101",
20111=>"100000000",
20112=>"111011000",
20113=>"000100111",
20114=>"100000100",
20115=>"111001111",
20116=>"111000000",
20117=>"001000101",
20118=>"001111111",
20119=>"011000000",
20120=>"011001001",
20121=>"100110010",
20122=>"000110111",
20123=>"110001111",
20124=>"011001011",
20125=>"111100001",
20126=>"000000111",
20127=>"101000111",
20128=>"001111111",
20129=>"110110010",
20130=>"110000000",
20131=>"101111111",
20132=>"001111000",
20133=>"000000000",
20134=>"100000000",
20135=>"001000000",
20136=>"010000111",
20137=>"000000111",
20138=>"101111111",
20139=>"000000111",
20140=>"111000001",
20141=>"000000111",
20142=>"100110011",
20143=>"111001110",
20144=>"000001001",
20145=>"011000110",
20146=>"101001001",
20147=>"101001100",
20148=>"110111000",
20149=>"111111111",
20150=>"000101111",
20151=>"101110011",
20152=>"110011001",
20153=>"110001000",
20154=>"010000010",
20155=>"111111110",
20156=>"011001011",
20157=>"111111111",
20158=>"100001011",
20159=>"000000000",
20160=>"010110001",
20161=>"111000101",
20162=>"111000000",
20163=>"010001111",
20164=>"000000011",
20165=>"100001001",
20166=>"111111000",
20167=>"010010101",
20168=>"010101101",
20169=>"000011011",
20170=>"110011111",
20171=>"000110111",
20172=>"000000111",
20173=>"100100110",
20174=>"111110000",
20175=>"001111110",
20176=>"111111111",
20177=>"111100110",
20178=>"000000101",
20179=>"101101001",
20180=>"000000111",
20181=>"111111101",
20182=>"111000001",
20183=>"001000000",
20184=>"111000000",
20185=>"011000000",
20186=>"100110111",
20187=>"001001111",
20188=>"111111100",
20189=>"010110000",
20190=>"000001001",
20191=>"000000101",
20192=>"001001011",
20193=>"000000111",
20194=>"110111111",
20195=>"000100011",
20196=>"111001001",
20197=>"011111101",
20198=>"001001000",
20199=>"111111000",
20200=>"001000000",
20201=>"111111111",
20202=>"001100100",
20203=>"000101111",
20204=>"011111111",
20205=>"000001000",
20206=>"000000111",
20207=>"111101101",
20208=>"111000100",
20209=>"001000100",
20210=>"000101001",
20211=>"110101000",
20212=>"111010000",
20213=>"111111101",
20214=>"101000010",
20215=>"100000000",
20216=>"001001111",
20217=>"001111110",
20218=>"111110010",
20219=>"000110000",
20220=>"101111100",
20221=>"010000000",
20222=>"000101011",
20223=>"001000000",
20224=>"001010111",
20225=>"010000101",
20226=>"000000101",
20227=>"000100110",
20228=>"011011110",
20229=>"011111000",
20230=>"111111001",
20231=>"111011100",
20232=>"011111000",
20233=>"111100000",
20234=>"000000000",
20235=>"111000000",
20236=>"111111010",
20237=>"110011001",
20238=>"000001001",
20239=>"111111001",
20240=>"011011111",
20241=>"101000111",
20242=>"110000000",
20243=>"110000000",
20244=>"111111111",
20245=>"011001101",
20246=>"000010111",
20247=>"101010011",
20248=>"100000000",
20249=>"011101001",
20250=>"010010100",
20251=>"010111111",
20252=>"111111111",
20253=>"000101101",
20254=>"010000000",
20255=>"001010100",
20256=>"100010000",
20257=>"111111100",
20258=>"000000100",
20259=>"111110000",
20260=>"111011011",
20261=>"010100100",
20262=>"000000101",
20263=>"011111011",
20264=>"000000111",
20265=>"000111110",
20266=>"101111101",
20267=>"000000011",
20268=>"111111111",
20269=>"111111100",
20270=>"111000100",
20271=>"000100100",
20272=>"000110111",
20273=>"111011000",
20274=>"000000000",
20275=>"001000011",
20276=>"000000111",
20277=>"000000001",
20278=>"000001011",
20279=>"001000111",
20280=>"000001111",
20281=>"000000111",
20282=>"111001000",
20283=>"000000000",
20284=>"110101000",
20285=>"111111000",
20286=>"000000000",
20287=>"010110000",
20288=>"111111110",
20289=>"101011000",
20290=>"101111111",
20291=>"010111110",
20292=>"111111111",
20293=>"011111111",
20294=>"111111010",
20295=>"010000110",
20296=>"110101111",
20297=>"111000000",
20298=>"100000001",
20299=>"000101110",
20300=>"110101000",
20301=>"111111111",
20302=>"001111001",
20303=>"111111100",
20304=>"000000000",
20305=>"111111000",
20306=>"011011010",
20307=>"000001111",
20308=>"111100000",
20309=>"000000001",
20310=>"100110111",
20311=>"001000000",
20312=>"011000000",
20313=>"000011000",
20314=>"110110110",
20315=>"111111111",
20316=>"100000100",
20317=>"100110111",
20318=>"111111111",
20319=>"000011001",
20320=>"000000000",
20321=>"001000100",
20322=>"110010000",
20323=>"011011001",
20324=>"001000111",
20325=>"000011010",
20326=>"000000110",
20327=>"011111111",
20328=>"111110111",
20329=>"111010000",
20330=>"111000000",
20331=>"111111101",
20332=>"000000000",
20333=>"011111111",
20334=>"001011000",
20335=>"011110001",
20336=>"110111100",
20337=>"000010111",
20338=>"000000100",
20339=>"000000111",
20340=>"110001111",
20341=>"001100101",
20342=>"010011111",
20343=>"000000000",
20344=>"010111110",
20345=>"010000000",
20346=>"000000101",
20347=>"111111000",
20348=>"000100000",
20349=>"000000110",
20350=>"111111111",
20351=>"000000100",
20352=>"000101110",
20353=>"111111100",
20354=>"010111000",
20355=>"001111111",
20356=>"010111111",
20357=>"000000111",
20358=>"000011011",
20359=>"110000010",
20360=>"101001100",
20361=>"011111111",
20362=>"110100111",
20363=>"111001100",
20364=>"000001111",
20365=>"111111010",
20366=>"100100000",
20367=>"000000000",
20368=>"100110111",
20369=>"110000000",
20370=>"000011111",
20371=>"100001001",
20372=>"010101111",
20373=>"010000000",
20374=>"111010111",
20375=>"001011000",
20376=>"000000000",
20377=>"111111000",
20378=>"000000000",
20379=>"100000000",
20380=>"111111100",
20381=>"101001111",
20382=>"111011111",
20383=>"000001111",
20384=>"111111110",
20385=>"000000111",
20386=>"000000101",
20387=>"000000010",
20388=>"101001000",
20389=>"000100010",
20390=>"111000101",
20391=>"111001111",
20392=>"000001000",
20393=>"100000110",
20394=>"000011111",
20395=>"010000000",
20396=>"110101100",
20397=>"000000111",
20398=>"000001010",
20399=>"001000010",
20400=>"000000000",
20401=>"100100110",
20402=>"101100010",
20403=>"100110111",
20404=>"101111010",
20405=>"001000101",
20406=>"011100000",
20407=>"010110101",
20408=>"011010000",
20409=>"001110111",
20410=>"000001001",
20411=>"111000001",
20412=>"111100011",
20413=>"011111000",
20414=>"111111000",
20415=>"101001000",
20416=>"111000010",
20417=>"000000000",
20418=>"010000110",
20419=>"011001111",
20420=>"000000101",
20421=>"000000010",
20422=>"000111111",
20423=>"111111000",
20424=>"111011000",
20425=>"000101100",
20426=>"000000111",
20427=>"000000101",
20428=>"000000100",
20429=>"000101011",
20430=>"000001111",
20431=>"111111011",
20432=>"111111010",
20433=>"110000001",
20434=>"010110100",
20435=>"011111000",
20436=>"101000000",
20437=>"011001111",
20438=>"110111110",
20439=>"110100000",
20440=>"000000101",
20441=>"011010000",
20442=>"110111111",
20443=>"100000100",
20444=>"100011111",
20445=>"111111111",
20446=>"001000100",
20447=>"010100111",
20448=>"111111111",
20449=>"011011100",
20450=>"111111000",
20451=>"011111110",
20452=>"101000000",
20453=>"111111011",
20454=>"111011010",
20455=>"011000100",
20456=>"111110111",
20457=>"010000011",
20458=>"000000000",
20459=>"100000000",
20460=>"000100000",
20461=>"111011001",
20462=>"000100000",
20463=>"000000000",
20464=>"000000000",
20465=>"001000010",
20466=>"101000110",
20467=>"000110010",
20468=>"111000011",
20469=>"101000101",
20470=>"011000000",
20471=>"000100001",
20472=>"111111000",
20473=>"111111110",
20474=>"011110011",
20475=>"000000110",
20476=>"001000111",
20477=>"000000000",
20478=>"110000101",
20479=>"101000111",
20480=>"001001100",
20481=>"000111000",
20482=>"000000101",
20483=>"000100111",
20484=>"001000001",
20485=>"111000111",
20486=>"000001000",
20487=>"101001110",
20488=>"000111111",
20489=>"001111111",
20490=>"000111011",
20491=>"000000000",
20492=>"010010000",
20493=>"011000000",
20494=>"101011001",
20495=>"001000001",
20496=>"111111010",
20497=>"111111111",
20498=>"000001000",
20499=>"001111111",
20500=>"111100000",
20501=>"101111111",
20502=>"100001111",
20503=>"001001000",
20504=>"000000000",
20505=>"111111001",
20506=>"111011111",
20507=>"100000000",
20508=>"000000001",
20509=>"011010111",
20510=>"111101111",
20511=>"111000101",
20512=>"011000001",
20513=>"110010010",
20514=>"101101100",
20515=>"111000000",
20516=>"111111001",
20517=>"111100111",
20518=>"010111111",
20519=>"111111011",
20520=>"000111110",
20521=>"101111111",
20522=>"100010000",
20523=>"010010110",
20524=>"001111111",
20525=>"000010101",
20526=>"111111111",
20527=>"110000110",
20528=>"010000111",
20529=>"001011011",
20530=>"100000111",
20531=>"011111111",
20532=>"000000000",
20533=>"101011111",
20534=>"001000100",
20535=>"101100101",
20536=>"111100010",
20537=>"000000000",
20538=>"000000001",
20539=>"111101101",
20540=>"110110010",
20541=>"001111111",
20542=>"000000000",
20543=>"000100110",
20544=>"111101111",
20545=>"001000101",
20546=>"100111111",
20547=>"000100111",
20548=>"101101111",
20549=>"000111111",
20550=>"111111101",
20551=>"110110000",
20552=>"110000000",
20553=>"000110010",
20554=>"000010111",
20555=>"000001101",
20556=>"000100110",
20557=>"100100000",
20558=>"000100110",
20559=>"110111111",
20560=>"111000000",
20561=>"000111110",
20562=>"000000101",
20563=>"001001010",
20564=>"000001111",
20565=>"111110000",
20566=>"001011001",
20567=>"000100111",
20568=>"000100111",
20569=>"100011001",
20570=>"100001011",
20571=>"010000000",
20572=>"111111111",
20573=>"001001000",
20574=>"111100000",
20575=>"001011110",
20576=>"000000011",
20577=>"010001000",
20578=>"101000000",
20579=>"000000001",
20580=>"001101000",
20581=>"111111100",
20582=>"100010000",
20583=>"100111111",
20584=>"000000110",
20585=>"000000000",
20586=>"111111001",
20587=>"111101100",
20588=>"111101000",
20589=>"010110110",
20590=>"011000000",
20591=>"110111011",
20592=>"001101010",
20593=>"111010111",
20594=>"111100000",
20595=>"110100011",
20596=>"111111000",
20597=>"100100111",
20598=>"000000011",
20599=>"101100100",
20600=>"000000010",
20601=>"101100001",
20602=>"011111101",
20603=>"000000000",
20604=>"100111110",
20605=>"100101001",
20606=>"110010011",
20607=>"000000000",
20608=>"111000000",
20609=>"000000000",
20610=>"111111111",
20611=>"111100010",
20612=>"000010111",
20613=>"111111111",
20614=>"111011110",
20615=>"111111000",
20616=>"000111011",
20617=>"111101000",
20618=>"000111111",
20619=>"111010000",
20620=>"000001101",
20621=>"111111111",
20622=>"100000001",
20623=>"001100111",
20624=>"111110000",
20625=>"000000000",
20626=>"000000000",
20627=>"010111011",
20628=>"111111010",
20629=>"111110110",
20630=>"111101000",
20631=>"010101111",
20632=>"000100000",
20633=>"000000111",
20634=>"000000010",
20635=>"000001011",
20636=>"000110110",
20637=>"010000001",
20638=>"011000000",
20639=>"010000000",
20640=>"011011000",
20641=>"111100111",
20642=>"110110000",
20643=>"000001111",
20644=>"111010001",
20645=>"110010000",
20646=>"111111111",
20647=>"101111101",
20648=>"111101111",
20649=>"110110101",
20650=>"111000000",
20651=>"000011000",
20652=>"111111101",
20653=>"000001111",
20654=>"010100001",
20655=>"101111101",
20656=>"000000000",
20657=>"111111000",
20658=>"000000001",
20659=>"000110000",
20660=>"000010011",
20661=>"101101111",
20662=>"111111100",
20663=>"110111111",
20664=>"011001000",
20665=>"111111011",
20666=>"111100111",
20667=>"111000111",
20668=>"010100010",
20669=>"011101101",
20670=>"101011101",
20671=>"000111111",
20672=>"010010000",
20673=>"001000000",
20674=>"001110111",
20675=>"000101110",
20676=>"000000000",
20677=>"111110000",
20678=>"000100000",
20679=>"110000010",
20680=>"111111000",
20681=>"110101000",
20682=>"010100000",
20683=>"101001000",
20684=>"000111111",
20685=>"001111001",
20686=>"111101000",
20687=>"000000001",
20688=>"000111111",
20689=>"011110100",
20690=>"111110110",
20691=>"100000000",
20692=>"111010000",
20693=>"111100000",
20694=>"000101101",
20695=>"000011011",
20696=>"000000001",
20697=>"111111111",
20698=>"110110110",
20699=>"000000000",
20700=>"111000011",
20701=>"000111111",
20702=>"111111111",
20703=>"110111111",
20704=>"000010111",
20705=>"111000111",
20706=>"111000001",
20707=>"111100010",
20708=>"000111000",
20709=>"111101101",
20710=>"101100110",
20711=>"110100110",
20712=>"010000111",
20713=>"110110111",
20714=>"001001000",
20715=>"001101000",
20716=>"000111100",
20717=>"110000000",
20718=>"000010010",
20719=>"000000000",
20720=>"010010110",
20721=>"110010000",
20722=>"111110111",
20723=>"000110010",
20724=>"100011001",
20725=>"101101101",
20726=>"000000000",
20727=>"000010111",
20728=>"000000000",
20729=>"000000000",
20730=>"111111001",
20731=>"111111110",
20732=>"011010000",
20733=>"110000000",
20734=>"001001000",
20735=>"110000000",
20736=>"100110100",
20737=>"000000000",
20738=>"000010000",
20739=>"110101001",
20740=>"001001000",
20741=>"010000000",
20742=>"000000000",
20743=>"101101011",
20744=>"101000000",
20745=>"111101110",
20746=>"000000111",
20747=>"111001001",
20748=>"101101111",
20749=>"100101101",
20750=>"000000010",
20751=>"000111101",
20752=>"000001000",
20753=>"111000011",
20754=>"111111010",
20755=>"011100100",
20756=>"011010000",
20757=>"011000001",
20758=>"110111011",
20759=>"101010110",
20760=>"111101110",
20761=>"010011111",
20762=>"000010010",
20763=>"000111010",
20764=>"010111000",
20765=>"111101001",
20766=>"000000100",
20767=>"111010010",
20768=>"111110000",
20769=>"100001111",
20770=>"000111111",
20771=>"100011111",
20772=>"100100110",
20773=>"011011010",
20774=>"000010110",
20775=>"111001011",
20776=>"101001011",
20777=>"100001001",
20778=>"000000000",
20779=>"100100010",
20780=>"010010000",
20781=>"000000101",
20782=>"000111110",
20783=>"011101001",
20784=>"111101100",
20785=>"100100110",
20786=>"100101111",
20787=>"010000000",
20788=>"100000101",
20789=>"111011000",
20790=>"111000010",
20791=>"000100000",
20792=>"101101101",
20793=>"101101000",
20794=>"011001010",
20795=>"101010000",
20796=>"110011110",
20797=>"001010100",
20798=>"111000100",
20799=>"000000000",
20800=>"111111000",
20801=>"010010101",
20802=>"110000000",
20803=>"100000001",
20804=>"111111011",
20805=>"101101001",
20806=>"100000001",
20807=>"111000000",
20808=>"110110110",
20809=>"100100000",
20810=>"101101101",
20811=>"000000000",
20812=>"011010000",
20813=>"001001010",
20814=>"111011011",
20815=>"111111001",
20816=>"000100101",
20817=>"111110100",
20818=>"101100100",
20819=>"110011011",
20820=>"111100111",
20821=>"000000000",
20822=>"001111010",
20823=>"000100101",
20824=>"100001000",
20825=>"011011010",
20826=>"000001000",
20827=>"100100000",
20828=>"000000110",
20829=>"000100110",
20830=>"100010000",
20831=>"001000011",
20832=>"011011010",
20833=>"011001010",
20834=>"101101111",
20835=>"100001001",
20836=>"101001011",
20837=>"000100110",
20838=>"101101110",
20839=>"100101011",
20840=>"000000010",
20841=>"111000000",
20842=>"010000111",
20843=>"111111001",
20844=>"111110010",
20845=>"111001010",
20846=>"000000101",
20847=>"000111000",
20848=>"101100111",
20849=>"000000000",
20850=>"011000000",
20851=>"000001000",
20852=>"000100011",
20853=>"010000000",
20854=>"100000010",
20855=>"001001000",
20856=>"010010111",
20857=>"000011010",
20858=>"111000111",
20859=>"111100110",
20860=>"111010100",
20861=>"011100000",
20862=>"101100111",
20863=>"101000100",
20864=>"111100000",
20865=>"010100101",
20866=>"000101101",
20867=>"011111111",
20868=>"100000111",
20869=>"001001101",
20870=>"100110111",
20871=>"001010110",
20872=>"000000011",
20873=>"101111111",
20874=>"010000000",
20875=>"100010000",
20876=>"100100101",
20877=>"000011000",
20878=>"101100000",
20879=>"100000000",
20880=>"111011001",
20881=>"000100000",
20882=>"000100111",
20883=>"101100000",
20884=>"000110000",
20885=>"000100000",
20886=>"000000000",
20887=>"100100110",
20888=>"111101000",
20889=>"110000000",
20890=>"101000100",
20891=>"000010000",
20892=>"110101101",
20893=>"111100101",
20894=>"000100101",
20895=>"011101010",
20896=>"110010110",
20897=>"001111111",
20898=>"101000000",
20899=>"000101101",
20900=>"110001111",
20901=>"010011011",
20902=>"101111111",
20903=>"111111011",
20904=>"000100000",
20905=>"000001000",
20906=>"110111000",
20907=>"010101100",
20908=>"111111100",
20909=>"100101111",
20910=>"011011001",
20911=>"000000111",
20912=>"000101110",
20913=>"110001110",
20914=>"010100010",
20915=>"011000011",
20916=>"110110110",
20917=>"111010101",
20918=>"000010011",
20919=>"110111101",
20920=>"011010011",
20921=>"100011001",
20922=>"000111110",
20923=>"000100110",
20924=>"111011011",
20925=>"010101101",
20926=>"100000000",
20927=>"101000000",
20928=>"111111111",
20929=>"000000000",
20930=>"011111000",
20931=>"110100000",
20932=>"011101111",
20933=>"111110001",
20934=>"101100000",
20935=>"101000010",
20936=>"010111010",
20937=>"000010000",
20938=>"010011110",
20939=>"010000000",
20940=>"001000000",
20941=>"111110110",
20942=>"010111000",
20943=>"011101101",
20944=>"011111001",
20945=>"000001010",
20946=>"011011111",
20947=>"000110000",
20948=>"101001000",
20949=>"001001011",
20950=>"010011001",
20951=>"100000000",
20952=>"100000101",
20953=>"011000000",
20954=>"000010001",
20955=>"111101101",
20956=>"110110110",
20957=>"000101101",
20958=>"001111111",
20959=>"000000001",
20960=>"110011111",
20961=>"000100111",
20962=>"010001011",
20963=>"110100111",
20964=>"000000000",
20965=>"111101110",
20966=>"000101000",
20967=>"010110001",
20968=>"100101100",
20969=>"101011000",
20970=>"000000001",
20971=>"001101111",
20972=>"101000111",
20973=>"111101111",
20974=>"010000011",
20975=>"010111111",
20976=>"010000001",
20977=>"100100000",
20978=>"000111011",
20979=>"001010010",
20980=>"001001011",
20981=>"100100000",
20982=>"111100101",
20983=>"010000000",
20984=>"001101101",
20985=>"001111111",
20986=>"111111110",
20987=>"111000000",
20988=>"111000000",
20989=>"010010000",
20990=>"000100100",
20991=>"110010110",
20992=>"011101010",
20993=>"000001000",
20994=>"100000111",
20995=>"000000000",
20996=>"011111111",
20997=>"010000000",
20998=>"010010110",
20999=>"000010111",
21000=>"111101110",
21001=>"000001000",
21002=>"000100100",
21003=>"111001011",
21004=>"000000000",
21005=>"011111010",
21006=>"101011010",
21007=>"001101110",
21008=>"000010110",
21009=>"101000111",
21010=>"001101000",
21011=>"111000000",
21012=>"111111111",
21013=>"001000100",
21014=>"111100011",
21015=>"011000111",
21016=>"101100111",
21017=>"111101111",
21018=>"000100100",
21019=>"000111010",
21020=>"110111101",
21021=>"101000000",
21022=>"111111000",
21023=>"011001000",
21024=>"111111111",
21025=>"010111111",
21026=>"000000000",
21027=>"000011011",
21028=>"000000100",
21029=>"111100111",
21030=>"111110101",
21031=>"001111101",
21032=>"010111001",
21033=>"010110000",
21034=>"111111101",
21035=>"111101010",
21036=>"001000000",
21037=>"110010111",
21038=>"111111011",
21039=>"000001100",
21040=>"001111111",
21041=>"000100011",
21042=>"011011111",
21043=>"110000100",
21044=>"000000000",
21045=>"111110101",
21046=>"010001011",
21047=>"000000111",
21048=>"111011000",
21049=>"000000001",
21050=>"000000011",
21051=>"111111100",
21052=>"110100111",
21053=>"000001001",
21054=>"010000001",
21055=>"111111011",
21056=>"111001000",
21057=>"101101011",
21058=>"000000000",
21059=>"001110000",
21060=>"110010010",
21061=>"000000111",
21062=>"101111111",
21063=>"001000111",
21064=>"110000000",
21065=>"111111000",
21066=>"111000000",
21067=>"000000101",
21068=>"000001000",
21069=>"001100111",
21070=>"111001111",
21071=>"111011111",
21072=>"111000111",
21073=>"010111101",
21074=>"000000010",
21075=>"001001100",
21076=>"111000000",
21077=>"010100100",
21078=>"000101001",
21079=>"000111111",
21080=>"110101000",
21081=>"111100010",
21082=>"110110111",
21083=>"111110111",
21084=>"000000000",
21085=>"111001011",
21086=>"010111100",
21087=>"101010100",
21088=>"100110000",
21089=>"000111011",
21090=>"000010100",
21091=>"001011011",
21092=>"111101101",
21093=>"001001000",
21094=>"001100000",
21095=>"111000000",
21096=>"111111111",
21097=>"011111000",
21098=>"010110111",
21099=>"111001000",
21100=>"111111110",
21101=>"000000001",
21102=>"111110000",
21103=>"000101011",
21104=>"000110100",
21105=>"001000011",
21106=>"010100110",
21107=>"001000100",
21108=>"000000111",
21109=>"101000000",
21110=>"000111111",
21111=>"111000000",
21112=>"111111111",
21113=>"000000000",
21114=>"000110111",
21115=>"000010000",
21116=>"000111000",
21117=>"110100001",
21118=>"001101111",
21119=>"111111111",
21120=>"000111000",
21121=>"111000001",
21122=>"111111110",
21123=>"111111000",
21124=>"110000000",
21125=>"111111000",
21126=>"110001110",
21127=>"000001011",
21128=>"011011111",
21129=>"111000010",
21130=>"111111111",
21131=>"001001111",
21132=>"000000001",
21133=>"000000100",
21134=>"010111111",
21135=>"000000100",
21136=>"110110100",
21137=>"001000000",
21138=>"000000101",
21139=>"000000011",
21140=>"100111111",
21141=>"000111100",
21142=>"000010000",
21143=>"001000000",
21144=>"010111100",
21145=>"111000000",
21146=>"111011000",
21147=>"001000000",
21148=>"111010100",
21149=>"111000101",
21150=>"010011111",
21151=>"101100000",
21152=>"010100000",
21153=>"010010111",
21154=>"111011010",
21155=>"010010000",
21156=>"000001010",
21157=>"111111110",
21158=>"000000010",
21159=>"100111010",
21160=>"111000110",
21161=>"000000000",
21162=>"001100101",
21163=>"110101010",
21164=>"001111000",
21165=>"100000010",
21166=>"110100000",
21167=>"000000000",
21168=>"011000000",
21169=>"011000100",
21170=>"010001000",
21171=>"101100000",
21172=>"101001000",
21173=>"111111110",
21174=>"011111111",
21175=>"011001101",
21176=>"001001011",
21177=>"001111101",
21178=>"111011001",
21179=>"110110111",
21180=>"000100100",
21181=>"111111110",
21182=>"111110011",
21183=>"101000000",
21184=>"010000000",
21185=>"011010010",
21186=>"000100011",
21187=>"011111000",
21188=>"000011000",
21189=>"110110100",
21190=>"010011101",
21191=>"111001000",
21192=>"101111111",
21193=>"000000000",
21194=>"111111111",
21195=>"111111001",
21196=>"111111111",
21197=>"110111110",
21198=>"101001110",
21199=>"010110111",
21200=>"010000000",
21201=>"110000110",
21202=>"010010111",
21203=>"000111010",
21204=>"001000101",
21205=>"010000001",
21206=>"111111000",
21207=>"010110110",
21208=>"111000111",
21209=>"000000010",
21210=>"011011011",
21211=>"000000000",
21212=>"010011111",
21213=>"011111111",
21214=>"111111000",
21215=>"010101111",
21216=>"000111011",
21217=>"000010111",
21218=>"111000001",
21219=>"011000111",
21220=>"111100101",
21221=>"000100000",
21222=>"001000010",
21223=>"011100101",
21224=>"000101010",
21225=>"000000011",
21226=>"100101001",
21227=>"000111000",
21228=>"111111010",
21229=>"111101111",
21230=>"001010001",
21231=>"000111111",
21232=>"000000000",
21233=>"011001001",
21234=>"111000000",
21235=>"110100000",
21236=>"010000111",
21237=>"101110111",
21238=>"101100111",
21239=>"100011000",
21240=>"000001010",
21241=>"000111001",
21242=>"111111111",
21243=>"000000000",
21244=>"000000110",
21245=>"111111000",
21246=>"100101010",
21247=>"010000101",
21248=>"010101101",
21249=>"110110100",
21250=>"111100100",
21251=>"111000011",
21252=>"110100100",
21253=>"111101000",
21254=>"000001010",
21255=>"010111011",
21256=>"000001011",
21257=>"110100100",
21258=>"100100110",
21259=>"000011011",
21260=>"000001001",
21261=>"100101101",
21262=>"111011001",
21263=>"001101111",
21264=>"111110110",
21265=>"011100110",
21266=>"011110000",
21267=>"001011000",
21268=>"000011010",
21269=>"111100101",
21270=>"110110010",
21271=>"100011001",
21272=>"000100110",
21273=>"001011011",
21274=>"000110100",
21275=>"111110110",
21276=>"011000000",
21277=>"011110111",
21278=>"000100000",
21279=>"100111011",
21280=>"111110100",
21281=>"100101101",
21282=>"010000000",
21283=>"001011011",
21284=>"100011011",
21285=>"001000010",
21286=>"000011011",
21287=>"000011011",
21288=>"111100111",
21289=>"000100100",
21290=>"100100001",
21291=>"111100100",
21292=>"000011000",
21293=>"010001011",
21294=>"000100100",
21295=>"001001101",
21296=>"000011000",
21297=>"100000100",
21298=>"111111011",
21299=>"000110100",
21300=>"111100100",
21301=>"111111111",
21302=>"110110110",
21303=>"100100100",
21304=>"000100000",
21305=>"000000001",
21306=>"000011011",
21307=>"100110110",
21308=>"001011011",
21309=>"001011001",
21310=>"001000000",
21311=>"000000111",
21312=>"111011000",
21313=>"000100110",
21314=>"110100110",
21315=>"111100100",
21316=>"000001000",
21317=>"010011001",
21318=>"011000011",
21319=>"110011001",
21320=>"110001000",
21321=>"011011100",
21322=>"000111011",
21323=>"111100111",
21324=>"110101000",
21325=>"000000101",
21326=>"100111111",
21327=>"111110101",
21328=>"111110101",
21329=>"011111000",
21330=>"011011011",
21331=>"001001000",
21332=>"111001111",
21333=>"001110000",
21334=>"010111111",
21335=>"011000000",
21336=>"101011011",
21337=>"000001001",
21338=>"110000001",
21339=>"100000011",
21340=>"110100100",
21341=>"011000000",
21342=>"111110110",
21343=>"111100000",
21344=>"000000001",
21345=>"111110100",
21346=>"010100100",
21347=>"111110110",
21348=>"000000011",
21349=>"000001100",
21350=>"110100001",
21351=>"111010000",
21352=>"000111111",
21353=>"011000100",
21354=>"111100111",
21355=>"011011001",
21356=>"011111100",
21357=>"001100100",
21358=>"000000001",
21359=>"010000011",
21360=>"000000000",
21361=>"000100011",
21362=>"110100100",
21363=>"001011011",
21364=>"000100100",
21365=>"001100000",
21366=>"111100001",
21367=>"000000101",
21368=>"010100000",
21369=>"010101011",
21370=>"000100001",
21371=>"000011100",
21372=>"111001001",
21373=>"000010010",
21374=>"111100110",
21375=>"100100100",
21376=>"001101100",
21377=>"000110110",
21378=>"110011000",
21379=>"010011011",
21380=>"000010001",
21381=>"111010110",
21382=>"000000001",
21383=>"010110010",
21384=>"101011011",
21385=>"000100111",
21386=>"110110110",
21387=>"011011100",
21388=>"110110110",
21389=>"111100100",
21390=>"011011000",
21391=>"111100111",
21392=>"110010010",
21393=>"101110110",
21394=>"111110011",
21395=>"111111000",
21396=>"001011010",
21397=>"111100100",
21398=>"100001111",
21399=>"011100110",
21400=>"110011001",
21401=>"000011011",
21402=>"000001001",
21403=>"111100100",
21404=>"000001001",
21405=>"110100100",
21406=>"111100010",
21407=>"011111001",
21408=>"100100010",
21409=>"111110100",
21410=>"110110110",
21411=>"011001011",
21412=>"000100001",
21413=>"010011011",
21414=>"011011010",
21415=>"010100000",
21416=>"011000000",
21417=>"111110111",
21418=>"111100100",
21419=>"000100100",
21420=>"110011000",
21421=>"000001001",
21422=>"000111110",
21423=>"100110010",
21424=>"000000000",
21425=>"111100100",
21426=>"001111110",
21427=>"000001010",
21428=>"101001011",
21429=>"110101110",
21430=>"000001000",
21431=>"110000001",
21432=>"110001011",
21433=>"000010000",
21434=>"001011011",
21435=>"000011100",
21436=>"100001001",
21437=>"000111110",
21438=>"011010000",
21439=>"001001001",
21440=>"100000000",
21441=>"000100111",
21442=>"111110110",
21443=>"100100111",
21444=>"000010001",
21445=>"110100000",
21446=>"011011011",
21447=>"111100100",
21448=>"000011111",
21449=>"110100100",
21450=>"011011110",
21451=>"111100100",
21452=>"100100110",
21453=>"011100001",
21454=>"100100001",
21455=>"110111011",
21456=>"000001001",
21457=>"000000001",
21458=>"111000001",
21459=>"000000010",
21460=>"011100100",
21461=>"101000000",
21462=>"010011011",
21463=>"001011110",
21464=>"001011111",
21465=>"100001000",
21466=>"000010110",
21467=>"111100110",
21468=>"101010001",
21469=>"000011011",
21470=>"001001011",
21471=>"000110100",
21472=>"100000100",
21473=>"001011010",
21474=>"110001000",
21475=>"011110000",
21476=>"011000100",
21477=>"111100100",
21478=>"000011011",
21479=>"100011001",
21480=>"100000001",
21481=>"011000000",
21482=>"111001001",
21483=>"011110110",
21484=>"100100100",
21485=>"000001001",
21486=>"000000010",
21487=>"111101000",
21488=>"001011010",
21489=>"000010010",
21490=>"000000000",
21491=>"011011111",
21492=>"001010110",
21493=>"001100000",
21494=>"001000001",
21495=>"011100000",
21496=>"010110111",
21497=>"000111111",
21498=>"001011011",
21499=>"000011000",
21500=>"000000000",
21501=>"111110110",
21502=>"100111100",
21503=>"111100000",
21504=>"001011001",
21505=>"101001011",
21506=>"101111111",
21507=>"001000000",
21508=>"110111000",
21509=>"000000101",
21510=>"011011010",
21511=>"111110110",
21512=>"001000100",
21513=>"000000000",
21514=>"000000100",
21515=>"111111001",
21516=>"111111101",
21517=>"000000000",
21518=>"111110011",
21519=>"111111111",
21520=>"101101110",
21521=>"000000000",
21522=>"000000000",
21523=>"011111111",
21524=>"000111011",
21525=>"000000010",
21526=>"011011000",
21527=>"111111010",
21528=>"000000000",
21529=>"000011000",
21530=>"101111111",
21531=>"111011100",
21532=>"111111110",
21533=>"111111111",
21534=>"000000111",
21535=>"001001111",
21536=>"100001000",
21537=>"001000001",
21538=>"101100000",
21539=>"111111111",
21540=>"110111000",
21541=>"111111110",
21542=>"000010111",
21543=>"111111100",
21544=>"000101111",
21545=>"000001010",
21546=>"100100100",
21547=>"101111001",
21548=>"111111111",
21549=>"000000000",
21550=>"111100101",
21551=>"000001001",
21552=>"101101111",
21553=>"100100101",
21554=>"100000010",
21555=>"000100000",
21556=>"000000101",
21557=>"000111110",
21558=>"100000100",
21559=>"111110000",
21560=>"000000000",
21561=>"111000001",
21562=>"111111111",
21563=>"111111100",
21564=>"111111111",
21565=>"011111111",
21566=>"000000000",
21567=>"011010110",
21568=>"101100100",
21569=>"000001111",
21570=>"010000000",
21571=>"011000001",
21572=>"111011001",
21573=>"000000010",
21574=>"111111111",
21575=>"000000000",
21576=>"111011110",
21577=>"101101011",
21578=>"101000111",
21579=>"111111111",
21580=>"000000100",
21581=>"111111110",
21582=>"111100010",
21583=>"111111110",
21584=>"000000111",
21585=>"111111111",
21586=>"001101001",
21587=>"001111001",
21588=>"000000001",
21589=>"110111111",
21590=>"111100000",
21591=>"000000100",
21592=>"100111100",
21593=>"111111101",
21594=>"000011011",
21595=>"101111011",
21596=>"000000001",
21597=>"001001001",
21598=>"011000100",
21599=>"100000001",
21600=>"000010111",
21601=>"101101101",
21602=>"000110111",
21603=>"000100100",
21604=>"110010000",
21605=>"111111100",
21606=>"111000000",
21607=>"000000000",
21608=>"110001001",
21609=>"000110000",
21610=>"001000000",
21611=>"010011111",
21612=>"111001000",
21613=>"000000010",
21614=>"111101000",
21615=>"111011000",
21616=>"011011010",
21617=>"111100000",
21618=>"011000001",
21619=>"000000111",
21620=>"000000111",
21621=>"000000001",
21622=>"100110111",
21623=>"100000000",
21624=>"111011000",
21625=>"000011000",
21626=>"001110110",
21627=>"001111010",
21628=>"110100010",
21629=>"100100110",
21630=>"111011010",
21631=>"000010111",
21632=>"111001001",
21633=>"100100000",
21634=>"000111111",
21635=>"111111111",
21636=>"000000110",
21637=>"111111011",
21638=>"101001001",
21639=>"001100110",
21640=>"100100101",
21641=>"111110011",
21642=>"000000001",
21643=>"000000000",
21644=>"100000001",
21645=>"000111000",
21646=>"111111001",
21647=>"000001010",
21648=>"100100000",
21649=>"000000001",
21650=>"110000101",
21651=>"111101111",
21652=>"111101101",
21653=>"000000100",
21654=>"111111101",
21655=>"100000000",
21656=>"111111000",
21657=>"111111111",
21658=>"000111111",
21659=>"000010000",
21660=>"011001101",
21661=>"100000111",
21662=>"111000010",
21663=>"111111000",
21664=>"001110100",
21665=>"001001011",
21666=>"101100101",
21667=>"111111011",
21668=>"001111111",
21669=>"001011101",
21670=>"111010010",
21671=>"101110000",
21672=>"000111001",
21673=>"000000000",
21674=>"000101010",
21675=>"000000000",
21676=>"101111011",
21677=>"000110111",
21678=>"110110110",
21679=>"010000000",
21680=>"101000111",
21681=>"011001001",
21682=>"000111111",
21683=>"000100000",
21684=>"111111000",
21685=>"000000000",
21686=>"111100111",
21687=>"111111011",
21688=>"111110111",
21689=>"111100110",
21690=>"010111111",
21691=>"110001111",
21692=>"000011010",
21693=>"000000010",
21694=>"000011011",
21695=>"000000000",
21696=>"000001000",
21697=>"110110100",
21698=>"000001001",
21699=>"001011011",
21700=>"110110010",
21701=>"111011001",
21702=>"111111111",
21703=>"000110111",
21704=>"111111010",
21705=>"111010000",
21706=>"000000111",
21707=>"101000000",
21708=>"000110111",
21709=>"001111011",
21710=>"000000110",
21711=>"000100000",
21712=>"011011010",
21713=>"011000001",
21714=>"000100101",
21715=>"111111101",
21716=>"010111101",
21717=>"000100100",
21718=>"000000101",
21719=>"111000000",
21720=>"111111010",
21721=>"011000000",
21722=>"100100001",
21723=>"000000000",
21724=>"111111000",
21725=>"011100000",
21726=>"011111100",
21727=>"111100110",
21728=>"000011001",
21729=>"001000101",
21730=>"111111111",
21731=>"000111110",
21732=>"000000000",
21733=>"000111111",
21734=>"111110100",
21735=>"011011011",
21736=>"000000000",
21737=>"011000111",
21738=>"000000001",
21739=>"101111111",
21740=>"100111111",
21741=>"010000000",
21742=>"010010010",
21743=>"010111111",
21744=>"111111111",
21745=>"000100100",
21746=>"011001001",
21747=>"111111101",
21748=>"110100100",
21749=>"000000000",
21750=>"000000111",
21751=>"111111111",
21752=>"111000000",
21753=>"101001110",
21754=>"000101000",
21755=>"111111111",
21756=>"000111111",
21757=>"011101111",
21758=>"001011101",
21759=>"010010010",
21760=>"000001001",
21761=>"011111111",
21762=>"000000000",
21763=>"100111111",
21764=>"001100101",
21765=>"111101111",
21766=>"110000100",
21767=>"101000111",
21768=>"000100111",
21769=>"010000000",
21770=>"110011001",
21771=>"001000011",
21772=>"011001101",
21773=>"011010000",
21774=>"100000100",
21775=>"111000000",
21776=>"111111000",
21777=>"010010000",
21778=>"000000000",
21779=>"111111111",
21780=>"000111101",
21781=>"101111010",
21782=>"000000100",
21783=>"111111000",
21784=>"111111101",
21785=>"101111110",
21786=>"111110010",
21787=>"000111111",
21788=>"000011000",
21789=>"010010000",
21790=>"110101101",
21791=>"001000011",
21792=>"000000000",
21793=>"010101111",
21794=>"010010100",
21795=>"000010110",
21796=>"110110111",
21797=>"000010111",
21798=>"111110010",
21799=>"111101000",
21800=>"101000101",
21801=>"001101111",
21802=>"000000000",
21803=>"101111111",
21804=>"100000110",
21805=>"111111011",
21806=>"000000001",
21807=>"101101001",
21808=>"110111000",
21809=>"011101000",
21810=>"101110111",
21811=>"101000000",
21812=>"111111000",
21813=>"111001000",
21814=>"111111110",
21815=>"000111111",
21816=>"000111100",
21817=>"000000111",
21818=>"000000110",
21819=>"111110000",
21820=>"001000110",
21821=>"000101011",
21822=>"000000100",
21823=>"111111111",
21824=>"111010000",
21825=>"011101111",
21826=>"000111000",
21827=>"001100001",
21828=>"111000000",
21829=>"000000000",
21830=>"010000001",
21831=>"111000000",
21832=>"001111111",
21833=>"101001010",
21834=>"100111101",
21835=>"101111000",
21836=>"000010111",
21837=>"001001110",
21838=>"100100000",
21839=>"111111111",
21840=>"001000111",
21841=>"011111000",
21842=>"011100010",
21843=>"001000001",
21844=>"110110000",
21845=>"000101100",
21846=>"011011001",
21847=>"000000000",
21848=>"000001111",
21849=>"001001011",
21850=>"100100011",
21851=>"111110011",
21852=>"000001111",
21853=>"000000111",
21854=>"111010000",
21855=>"000100110",
21856=>"111101000",
21857=>"001000000",
21858=>"000111111",
21859=>"001001110",
21860=>"001100111",
21861=>"000000000",
21862=>"100111101",
21863=>"000111010",
21864=>"111000000",
21865=>"000000101",
21866=>"100000111",
21867=>"000101111",
21868=>"111100111",
21869=>"110110010",
21870=>"000100001",
21871=>"001110110",
21872=>"100101111",
21873=>"101100000",
21874=>"111011001",
21875=>"111000000",
21876=>"111111000",
21877=>"101111010",
21878=>"111000000",
21879=>"111111000",
21880=>"111101010",
21881=>"110001101",
21882=>"000001000",
21883=>"111101000",
21884=>"000001111",
21885=>"100000100",
21886=>"100000000",
21887=>"000000101",
21888=>"000000000",
21889=>"000001011",
21890=>"111111111",
21891=>"011111110",
21892=>"000000100",
21893=>"000010000",
21894=>"000110011",
21895=>"100000011",
21896=>"001100110",
21897=>"010111101",
21898=>"010011111",
21899=>"101100000",
21900=>"000000111",
21901=>"000000111",
21902=>"000001111",
21903=>"001001000",
21904=>"001001011",
21905=>"101001100",
21906=>"111000010",
21907=>"010010010",
21908=>"000010101",
21909=>"000101001",
21910=>"000101111",
21911=>"000001011",
21912=>"111111111",
21913=>"000001111",
21914=>"111000000",
21915=>"111000000",
21916=>"000000101",
21917=>"111001111",
21918=>"111111011",
21919=>"000000000",
21920=>"101111011",
21921=>"000000000",
21922=>"100101110",
21923=>"111111111",
21924=>"110000100",
21925=>"111110100",
21926=>"100000000",
21927=>"101000011",
21928=>"001111110",
21929=>"000000111",
21930=>"100000101",
21931=>"111000000",
21932=>"010111110",
21933=>"000000101",
21934=>"000000110",
21935=>"011000001",
21936=>"101111101",
21937=>"001001111",
21938=>"111111110",
21939=>"000110111",
21940=>"111111000",
21941=>"111000000",
21942=>"111111000",
21943=>"101000100",
21944=>"100100111",
21945=>"000000110",
21946=>"000000110",
21947=>"111010000",
21948=>"000110111",
21949=>"111110010",
21950=>"101111011",
21951=>"000101100",
21952=>"111111000",
21953=>"011111111",
21954=>"100111001",
21955=>"100100110",
21956=>"111111001",
21957=>"100000111",
21958=>"010010110",
21959=>"111000000",
21960=>"000000000",
21961=>"100000000",
21962=>"101000110",
21963=>"111111001",
21964=>"011111101",
21965=>"000100011",
21966=>"111001101",
21967=>"000011111",
21968=>"111010000",
21969=>"000100111",
21970=>"000000111",
21971=>"100100001",
21972=>"000000111",
21973=>"000110111",
21974=>"000001111",
21975=>"111111111",
21976=>"111111000",
21977=>"000010010",
21978=>"111100100",
21979=>"111000000",
21980=>"000111001",
21981=>"000000111",
21982=>"111111100",
21983=>"110111100",
21984=>"111101000",
21985=>"000101111",
21986=>"111011000",
21987=>"000000001",
21988=>"000001010",
21989=>"101111101",
21990=>"000000111",
21991=>"000000111",
21992=>"111100000",
21993=>"000000000",
21994=>"110110100",
21995=>"111111000",
21996=>"111111111",
21997=>"111010000",
21998=>"000000000",
21999=>"000111110",
22000=>"000000011",
22001=>"011001111",
22002=>"010111111",
22003=>"111100110",
22004=>"100111011",
22005=>"101100100",
22006=>"000100111",
22007=>"000100100",
22008=>"111001101",
22009=>"101000110",
22010=>"111111111",
22011=>"111000011",
22012=>"011111000",
22013=>"000000000",
22014=>"100111011",
22015=>"000000101",
22016=>"001111011",
22017=>"011000011",
22018=>"100000000",
22019=>"111010000",
22020=>"000111100",
22021=>"101001000",
22022=>"111001000",
22023=>"100000101",
22024=>"000010010",
22025=>"000000101",
22026=>"000000101",
22027=>"010111000",
22028=>"000010111",
22029=>"000111111",
22030=>"100100100",
22031=>"110100010",
22032=>"110010000",
22033=>"100000001",
22034=>"111000100",
22035=>"001000101",
22036=>"111110101",
22037=>"100100101",
22038=>"011010110",
22039=>"000000000",
22040=>"001000001",
22041=>"000100010",
22042=>"010111110",
22043=>"000011111",
22044=>"110001111",
22045=>"000000100",
22046=>"000100000",
22047=>"000111010",
22048=>"111111110",
22049=>"011111000",
22050=>"000110111",
22051=>"011000000",
22052=>"001111111",
22053=>"000010011",
22054=>"000110111",
22055=>"101000000",
22056=>"110110000",
22057=>"000101001",
22058=>"111111101",
22059=>"001000000",
22060=>"100100000",
22061=>"111000101",
22062=>"111010100",
22063=>"000101101",
22064=>"000101011",
22065=>"000001101",
22066=>"010011010",
22067=>"111101000",
22068=>"001001000",
22069=>"001010110",
22070=>"100000101",
22071=>"010010100",
22072=>"111001111",
22073=>"001001101",
22074=>"011000000",
22075=>"101101001",
22076=>"010011111",
22077=>"111011000",
22078=>"000000000",
22079=>"011011001",
22080=>"000111111",
22081=>"000001110",
22082=>"101000000",
22083=>"001100011",
22084=>"011010011",
22085=>"011000000",
22086=>"101101101",
22087=>"110110000",
22088=>"100001101",
22089=>"100000100",
22090=>"000000000",
22091=>"111010000",
22092=>"111000110",
22093=>"101111110",
22094=>"001110011",
22095=>"010000101",
22096=>"101100000",
22097=>"011011000",
22098=>"110001111",
22099=>"011001001",
22100=>"010000110",
22101=>"111100000",
22102=>"001101011",
22103=>"101000101",
22104=>"001101111",
22105=>"000100110",
22106=>"000001111",
22107=>"010011011",
22108=>"000110110",
22109=>"000001000",
22110=>"111011000",
22111=>"100111010",
22112=>"001101111",
22113=>"110111101",
22114=>"101000101",
22115=>"111100111",
22116=>"011111100",
22117=>"001101000",
22118=>"000001000",
22119=>"000010001",
22120=>"111110110",
22121=>"111100101",
22122=>"110111000",
22123=>"111000010",
22124=>"000110110",
22125=>"001001000",
22126=>"000000011",
22127=>"110000000",
22128=>"100110100",
22129=>"000000111",
22130=>"001001101",
22131=>"000010111",
22132=>"111100000",
22133=>"111101000",
22134=>"011101000",
22135=>"000111111",
22136=>"000000111",
22137=>"111011111",
22138=>"000110011",
22139=>"000111110",
22140=>"001001001",
22141=>"011101000",
22142=>"000100000",
22143=>"000110000",
22144=>"000111111",
22145=>"111000000",
22146=>"000011111",
22147=>"000000000",
22148=>"111001101",
22149=>"111001000",
22150=>"000000000",
22151=>"000011011",
22152=>"000111110",
22153=>"000000010",
22154=>"000000100",
22155=>"111010000",
22156=>"010111010",
22157=>"101111110",
22158=>"010110111",
22159=>"000000110",
22160=>"101111111",
22161=>"000111111",
22162=>"000001000",
22163=>"111001000",
22164=>"110101010",
22165=>"101001111",
22166=>"111101111",
22167=>"000011010",
22168=>"111000000",
22169=>"000000000",
22170=>"000111011",
22171=>"111001000",
22172=>"111101111",
22173=>"000000000",
22174=>"010111000",
22175=>"111000000",
22176=>"011111111",
22177=>"110110111",
22178=>"000111110",
22179=>"000100111",
22180=>"110011100",
22181=>"100110111",
22182=>"110110000",
22183=>"001001100",
22184=>"101000000",
22185=>"011111010",
22186=>"001101111",
22187=>"101000011",
22188=>"101110010",
22189=>"101001101",
22190=>"111111000",
22191=>"110110000",
22192=>"000110100",
22193=>"001011111",
22194=>"111000010",
22195=>"001101010",
22196=>"011011000",
22197=>"111111110",
22198=>"000010100",
22199=>"001010010",
22200=>"001011111",
22201=>"000000000",
22202=>"000110001",
22203=>"010010010",
22204=>"100000000",
22205=>"101111010",
22206=>"010011010",
22207=>"111111101",
22208=>"101000000",
22209=>"101001101",
22210=>"101101111",
22211=>"001011011",
22212=>"011001001",
22213=>"110110001",
22214=>"000100100",
22215=>"001001101",
22216=>"001001000",
22217=>"000110110",
22218=>"101100111",
22219=>"100111010",
22220=>"010111110",
22221=>"100100000",
22222=>"000110000",
22223=>"100111000",
22224=>"001001001",
22225=>"000111111",
22226=>"000000100",
22227=>"001001010",
22228=>"111100000",
22229=>"000100100",
22230=>"101001111",
22231=>"101101110",
22232=>"110000000",
22233=>"010010111",
22234=>"001101111",
22235=>"101000010",
22236=>"001111001",
22237=>"000000100",
22238=>"110000110",
22239=>"110001101",
22240=>"000010110",
22241=>"111101001",
22242=>"111000000",
22243=>"001111111",
22244=>"000000001",
22245=>"010111100",
22246=>"111010010",
22247=>"010110111",
22248=>"111101000",
22249=>"110111101",
22250=>"000000000",
22251=>"000111001",
22252=>"000010101",
22253=>"010110111",
22254=>"101000000",
22255=>"000111100",
22256=>"110010000",
22257=>"111011001",
22258=>"111001000",
22259=>"101000011",
22260=>"110101100",
22261=>"101011001",
22262=>"000000111",
22263=>"000110000",
22264=>"111000000",
22265=>"111001011",
22266=>"010000110",
22267=>"111111101",
22268=>"111000100",
22269=>"010010010",
22270=>"000111011",
22271=>"111001101",
22272=>"010001001",
22273=>"000000000",
22274=>"010110010",
22275=>"000000000",
22276=>"000101001",
22277=>"000000010",
22278=>"010010000",
22279=>"000001010",
22280=>"111110110",
22281=>"000000000",
22282=>"001111111",
22283=>"101010000",
22284=>"111000100",
22285=>"011011001",
22286=>"101000011",
22287=>"111000111",
22288=>"001000000",
22289=>"000000001",
22290=>"100000110",
22291=>"000000010",
22292=>"000000001",
22293=>"000000000",
22294=>"001011010",
22295=>"000000100",
22296=>"000000001",
22297=>"000001001",
22298=>"010111111",
22299=>"011111011",
22300=>"011111111",
22301=>"111110010",
22302=>"000000000",
22303=>"111101110",
22304=>"000101011",
22305=>"000101001",
22306=>"110000111",
22307=>"110000111",
22308=>"011111011",
22309=>"010000010",
22310=>"000000100",
22311=>"001111011",
22312=>"111111111",
22313=>"111111010",
22314=>"001000001",
22315=>"101101000",
22316=>"111111001",
22317=>"000000000",
22318=>"110000010",
22319=>"011000000",
22320=>"000000000",
22321=>"111111111",
22322=>"111111010",
22323=>"000000000",
22324=>"000010000",
22325=>"001111000",
22326=>"000100100",
22327=>"001000000",
22328=>"000000000",
22329=>"100000000",
22330=>"100101111",
22331=>"111110111",
22332=>"100000000",
22333=>"111111111",
22334=>"000000010",
22335=>"000011110",
22336=>"001001000",
22337=>"111111111",
22338=>"111101001",
22339=>"000111011",
22340=>"111111000",
22341=>"000000000",
22342=>"010000000",
22343=>"110111100",
22344=>"000000000",
22345=>"101111011",
22346=>"111111001",
22347=>"001111001",
22348=>"000000011",
22349=>"111111110",
22350=>"111111111",
22351=>"111111011",
22352=>"000110111",
22353=>"000010010",
22354=>"000000000",
22355=>"011001000",
22356=>"010110110",
22357=>"000000000",
22358=>"111111111",
22359=>"000000000",
22360=>"111111010",
22361=>"000111111",
22362=>"101100101",
22363=>"000100111",
22364=>"111000000",
22365=>"001000011",
22366=>"011010110",
22367=>"101111000",
22368=>"010111111",
22369=>"101111000",
22370=>"101111000",
22371=>"100101111",
22372=>"110110110",
22373=>"111111011",
22374=>"101111111",
22375=>"110111111",
22376=>"010000000",
22377=>"000000000",
22378=>"000000000",
22379=>"111111110",
22380=>"110111111",
22381=>"111111111",
22382=>"001000000",
22383=>"000000010",
22384=>"000110011",
22385=>"000000000",
22386=>"000010010",
22387=>"111111111",
22388=>"000000000",
22389=>"000000001",
22390=>"000000000",
22391=>"111111111",
22392=>"010000111",
22393=>"010000000",
22394=>"001000001",
22395=>"100100100",
22396=>"000100010",
22397=>"100100000",
22398=>"010000000",
22399=>"110111111",
22400=>"000001111",
22401=>"000100000",
22402=>"000010010",
22403=>"111110111",
22404=>"000100101",
22405=>"000100101",
22406=>"011010111",
22407=>"011001000",
22408=>"001111111",
22409=>"101111111",
22410=>"101011111",
22411=>"110000000",
22412=>"111111000",
22413=>"000000001",
22414=>"010110110",
22415=>"101000000",
22416=>"100101111",
22417=>"111111111",
22418=>"000000000",
22419=>"011010000",
22420=>"111111111",
22421=>"000000000",
22422=>"111111111",
22423=>"001000011",
22424=>"010010100",
22425=>"000001110",
22426=>"001001011",
22427=>"000010010",
22428=>"000010010",
22429=>"100111101",
22430=>"000000000",
22431=>"000001000",
22432=>"001111101",
22433=>"001000000",
22434=>"111111111",
22435=>"111000100",
22436=>"000000000",
22437=>"110110110",
22438=>"111010000",
22439=>"111111011",
22440=>"000000101",
22441=>"000000010",
22442=>"111111110",
22443=>"000101111",
22444=>"111000100",
22445=>"110110010",
22446=>"110101111",
22447=>"010010110",
22448=>"010010010",
22449=>"101001001",
22450=>"111100000",
22451=>"000000110",
22452=>"111111111",
22453=>"111110101",
22454=>"000000000",
22455=>"010010010",
22456=>"011000000",
22457=>"111110100",
22458=>"110111110",
22459=>"000110010",
22460=>"001110110",
22461=>"101111000",
22462=>"011011011",
22463=>"010000000",
22464=>"010000000",
22465=>"000010100",
22466=>"000000010",
22467=>"111111100",
22468=>"010010011",
22469=>"100001101",
22470=>"000000000",
22471=>"111111011",
22472=>"111101111",
22473=>"011001111",
22474=>"111000000",
22475=>"000100111",
22476=>"001110000",
22477=>"000000000",
22478=>"000000000",
22479=>"000000000",
22480=>"000000010",
22481=>"111111110",
22482=>"110111111",
22483=>"110100110",
22484=>"010000000",
22485=>"100000000",
22486=>"010100100",
22487=>"000000000",
22488=>"111110110",
22489=>"000000111",
22490=>"110111111",
22491=>"000000000",
22492=>"000000000",
22493=>"000000010",
22494=>"010010001",
22495=>"000000000",
22496=>"011000001",
22497=>"000111000",
22498=>"111010110",
22499=>"101101111",
22500=>"001000001",
22501=>"101111000",
22502=>"100110000",
22503=>"111111101",
22504=>"000000000",
22505=>"110111111",
22506=>"101111110",
22507=>"000010000",
22508=>"000000010",
22509=>"001001100",
22510=>"010010010",
22511=>"111010110",
22512=>"010000010",
22513=>"111000011",
22514=>"000001100",
22515=>"101001100",
22516=>"110000000",
22517=>"111111111",
22518=>"000000010",
22519=>"000000000",
22520=>"000000000",
22521=>"000000010",
22522=>"011011000",
22523=>"111011111",
22524=>"111101111",
22525=>"110000111",
22526=>"111111101",
22527=>"000000111",
22528=>"001001000",
22529=>"111101101",
22530=>"011000111",
22531=>"001000000",
22532=>"000110110",
22533=>"000100011",
22534=>"111101101",
22535=>"110111011",
22536=>"000111010",
22537=>"101100000",
22538=>"000000000",
22539=>"111101000",
22540=>"001111011",
22541=>"101000000",
22542=>"000001100",
22543=>"010110000",
22544=>"011000010",
22545=>"100000010",
22546=>"011000100",
22547=>"011011000",
22548=>"111001001",
22549=>"101100100",
22550=>"110111001",
22551=>"111101011",
22552=>"101000000",
22553=>"000001110",
22554=>"010010000",
22555=>"011000100",
22556=>"000111011",
22557=>"000100100",
22558=>"101101111",
22559=>"001111010",
22560=>"000000000",
22561=>"011101111",
22562=>"100111000",
22563=>"000011111",
22564=>"000100110",
22565=>"110100111",
22566=>"111111111",
22567=>"101011000",
22568=>"111100111",
22569=>"111101101",
22570=>"101100100",
22571=>"010100100",
22572=>"101101111",
22573=>"000110111",
22574=>"100000110",
22575=>"110111011",
22576=>"000111111",
22577=>"001111111",
22578=>"001011011",
22579=>"110111100",
22580=>"000000000",
22581=>"111111010",
22582=>"110100100",
22583=>"000000010",
22584=>"010010000",
22585=>"101100101",
22586=>"001111111",
22587=>"110011010",
22588=>"101111011",
22589=>"011111010",
22590=>"100000100",
22591=>"100111111",
22592=>"111111111",
22593=>"010000001",
22594=>"000000010",
22595=>"001000110",
22596=>"111111010",
22597=>"111111101",
22598=>"000000000",
22599=>"111011100",
22600=>"000010111",
22601=>"000000010",
22602=>"111101101",
22603=>"111000001",
22604=>"111101101",
22605=>"000010010",
22606=>"000001111",
22607=>"011111111",
22608=>"001001001",
22609=>"111000111",
22610=>"111101101",
22611=>"111101101",
22612=>"101100100",
22613=>"000000010",
22614=>"101111010",
22615=>"110100100",
22616=>"111000000",
22617=>"101100101",
22618=>"100110111",
22619=>"000000000",
22620=>"000010111",
22621=>"000000000",
22622=>"111000010",
22623=>"100000111",
22624=>"111010011",
22625=>"110101010",
22626=>"000000010",
22627=>"001001000",
22628=>"100100010",
22629=>"000100100",
22630=>"111111111",
22631=>"011011001",
22632=>"111110010",
22633=>"000000000",
22634=>"000010011",
22635=>"100011111",
22636=>"000010101",
22637=>"000000111",
22638=>"010111011",
22639=>"111101111",
22640=>"111111101",
22641=>"000000111",
22642=>"111001000",
22643=>"000011000",
22644=>"000000000",
22645=>"001100101",
22646=>"010010111",
22647=>"111100101",
22648=>"010000000",
22649=>"011010000",
22650=>"100100000",
22651=>"000101010",
22652=>"010100111",
22653=>"100100100",
22654=>"101000011",
22655=>"101000100",
22656=>"111101000",
22657=>"000000011",
22658=>"000000011",
22659=>"011111101",
22660=>"111100100",
22661=>"111111101",
22662=>"001111111",
22663=>"001001000",
22664=>"001110100",
22665=>"001000101",
22666=>"111000101",
22667=>"111111001",
22668=>"000100000",
22669=>"101000000",
22670=>"000010001",
22671=>"111100110",
22672=>"100100100",
22673=>"010011011",
22674=>"001000010",
22675=>"000101000",
22676=>"000001010",
22677=>"011100101",
22678=>"001111011",
22679=>"001001011",
22680=>"000011111",
22681=>"000010000",
22682=>"110000001",
22683=>"111100101",
22684=>"011101100",
22685=>"100001000",
22686=>"010010110",
22687=>"000010101",
22688=>"000001001",
22689=>"111101000",
22690=>"000011010",
22691=>"100101101",
22692=>"010111101",
22693=>"010101100",
22694=>"010111000",
22695=>"001000001",
22696=>"111010000",
22697=>"010010000",
22698=>"111001011",
22699=>"111100000",
22700=>"110010000",
22701=>"101101100",
22702=>"101100001",
22703=>"000100110",
22704=>"010100010",
22705=>"000000011",
22706=>"011100100",
22707=>"001000000",
22708=>"000001010",
22709=>"111111000",
22710=>"011100100",
22711=>"000011000",
22712=>"000000010",
22713=>"100010010",
22714=>"111011001",
22715=>"110011000",
22716=>"000001011",
22717=>"000000011",
22718=>"100000100",
22719=>"110000010",
22720=>"011000000",
22721=>"111000100",
22722=>"010100011",
22723=>"001100011",
22724=>"101111010",
22725=>"110000110",
22726=>"111111010",
22727=>"100100111",
22728=>"000000101",
22729=>"111101000",
22730=>"000001100",
22731=>"000011011",
22732=>"011000110",
22733=>"110111111",
22734=>"101011000",
22735=>"110111010",
22736=>"010100111",
22737=>"000110110",
22738=>"010101110",
22739=>"000101000",
22740=>"010010010",
22741=>"000000111",
22742=>"011010111",
22743=>"000000011",
22744=>"011011011",
22745=>"110000000",
22746=>"111110110",
22747=>"100000100",
22748=>"101001001",
22749=>"110000000",
22750=>"011111000",
22751=>"000000000",
22752=>"111100000",
22753=>"101100000",
22754=>"010101100",
22755=>"100000000",
22756=>"111100101",
22757=>"111111101",
22758=>"000000000",
22759=>"101111110",
22760=>"000101011",
22761=>"010010000",
22762=>"000000000",
22763=>"100000111",
22764=>"111100000",
22765=>"000101110",
22766=>"000000001",
22767=>"000011010",
22768=>"000110010",
22769=>"001000001",
22770=>"111101101",
22771=>"001101100",
22772=>"111100100",
22773=>"101000000",
22774=>"000000010",
22775=>"110000100",
22776=>"011111111",
22777=>"010100011",
22778=>"000000000",
22779=>"101100010",
22780=>"000011011",
22781=>"000011011",
22782=>"000011011",
22783=>"101001101",
22784=>"000100100",
22785=>"001000000",
22786=>"110111010",
22787=>"000000000",
22788=>"001000101",
22789=>"101101001",
22790=>"111100101",
22791=>"000000000",
22792=>"000001000",
22793=>"111111101",
22794=>"111111111",
22795=>"000000000",
22796=>"111110110",
22797=>"000100111",
22798=>"000000000",
22799=>"111111111",
22800=>"010010000",
22801=>"000000000",
22802=>"111000000",
22803=>"000000000",
22804=>"111111111",
22805=>"110110111",
22806=>"010100101",
22807=>"111111101",
22808=>"000111111",
22809=>"100010000",
22810=>"111000111",
22811=>"111111111",
22812=>"111111111",
22813=>"111001111",
22814=>"000001111",
22815=>"100100100",
22816=>"111101111",
22817=>"111101111",
22818=>"111110000",
22819=>"111111110",
22820=>"000000100",
22821=>"000000001",
22822=>"110111110",
22823=>"000000111",
22824=>"111111001",
22825=>"000000101",
22826=>"000000101",
22827=>"100110000",
22828=>"000000000",
22829=>"000110111",
22830=>"000000000",
22831=>"101110001",
22832=>"000000000",
22833=>"001101100",
22834=>"011011011",
22835=>"000000000",
22836=>"100000100",
22837=>"111111111",
22838=>"111111111",
22839=>"000000111",
22840=>"101101000",
22841=>"000011001",
22842=>"011000101",
22843=>"000000000",
22844=>"000000000",
22845=>"111111101",
22846=>"111111111",
22847=>"000000000",
22848=>"010010001",
22849=>"000000001",
22850=>"111101001",
22851=>"110111111",
22852=>"111100111",
22853=>"000000101",
22854=>"001000101",
22855=>"001000111",
22856=>"010111111",
22857=>"111111101",
22858=>"000000001",
22859=>"110111111",
22860=>"000000000",
22861=>"100000011",
22862=>"011000001",
22863=>"000011111",
22864=>"111111111",
22865=>"111111111",
22866=>"000001000",
22867=>"000000110",
22868=>"110111000",
22869=>"000000000",
22870=>"000000000",
22871=>"111111111",
22872=>"001001100",
22873=>"000000000",
22874=>"000000000",
22875=>"000000000",
22876=>"000000100",
22877=>"100000100",
22878=>"111111110",
22879=>"000100001",
22880=>"000000000",
22881=>"000000100",
22882=>"111111100",
22883=>"000000000",
22884=>"001001001",
22885=>"001010000",
22886=>"000000111",
22887=>"011101101",
22888=>"000000000",
22889=>"000000000",
22890=>"000000111",
22891=>"011110111",
22892=>"000000001",
22893=>"111111111",
22894=>"111110000",
22895=>"000000000",
22896=>"000000000",
22897=>"000000001",
22898=>"111001001",
22899=>"101011100",
22900=>"000000101",
22901=>"010010000",
22902=>"000000001",
22903=>"011111011",
22904=>"111100111",
22905=>"001000000",
22906=>"000000101",
22907=>"111111111",
22908=>"000111000",
22909=>"000000001",
22910=>"111111111",
22911=>"111111010",
22912=>"000000000",
22913=>"111111111",
22914=>"000000000",
22915=>"001000101",
22916=>"100000101",
22917=>"000111011",
22918=>"000000010",
22919=>"000000000",
22920=>"000000001",
22921=>"000000111",
22922=>"000001001",
22923=>"000000000",
22924=>"111111110",
22925=>"111101101",
22926=>"111111011",
22927=>"000011000",
22928=>"000000100",
22929=>"000000000",
22930=>"001000000",
22931=>"000000101",
22932=>"000000000",
22933=>"111111000",
22934=>"110100100",
22935=>"000000001",
22936=>"000100001",
22937=>"000010001",
22938=>"111111110",
22939=>"000101100",
22940=>"000110111",
22941=>"100110111",
22942=>"010001110",
22943=>"111111001",
22944=>"111111010",
22945=>"000000000",
22946=>"001000101",
22947=>"111011111",
22948=>"001010101",
22949=>"000000100",
22950=>"000000100",
22951=>"111111111",
22952=>"000000000",
22953=>"000001111",
22954=>"111111111",
22955=>"110000000",
22956=>"001001111",
22957=>"000000000",
22958=>"111101101",
22959=>"100111110",
22960=>"000101001",
22961=>"000000010",
22962=>"111000111",
22963=>"010000000",
22964=>"000000001",
22965=>"111101111",
22966=>"000000000",
22967=>"000000000",
22968=>"000000000",
22969=>"000000001",
22970=>"000000000",
22971=>"000000000",
22972=>"000101111",
22973=>"111110110",
22974=>"000000000",
22975=>"111011101",
22976=>"110111111",
22977=>"111111111",
22978=>"000000010",
22979=>"101100101",
22980=>"000110010",
22981=>"010010111",
22982=>"001000000",
22983=>"111111111",
22984=>"000000001",
22985=>"111110000",
22986=>"000000010",
22987=>"100111000",
22988=>"000010110",
22989=>"000010000",
22990=>"111000000",
22991=>"000001101",
22992=>"110000000",
22993=>"000000000",
22994=>"001000000",
22995=>"111110100",
22996=>"000100000",
22997=>"000000001",
22998=>"111111110",
22999=>"001000000",
23000=>"111111111",
23001=>"101110110",
23002=>"001011011",
23003=>"111110000",
23004=>"000000001",
23005=>"100000111",
23006=>"111111111",
23007=>"010000010",
23008=>"111111010",
23009=>"000101111",
23010=>"111111111",
23011=>"000000000",
23012=>"000011000",
23013=>"110110111",
23014=>"000000000",
23015=>"000001000",
23016=>"010000101",
23017=>"111111000",
23018=>"101111111",
23019=>"111101111",
23020=>"111111000",
23021=>"111111000",
23022=>"110111000",
23023=>"111101101",
23024=>"111110000",
23025=>"100100111",
23026=>"001101111",
23027=>"000000000",
23028=>"000001011",
23029=>"110110111",
23030=>"101111111",
23031=>"001001101",
23032=>"111111111",
23033=>"000001000",
23034=>"111100101",
23035=>"000000000",
23036=>"111000111",
23037=>"111000111",
23038=>"000000100",
23039=>"110111000",
23040=>"110111011",
23041=>"000000000",
23042=>"000110111",
23043=>"001000100",
23044=>"001010010",
23045=>"101000000",
23046=>"111011110",
23047=>"000000000",
23048=>"000011010",
23049=>"000110110",
23050=>"001011011",
23051=>"101100111",
23052=>"100000101",
23053=>"001100110",
23054=>"000100110",
23055=>"111011011",
23056=>"111111001",
23057=>"000000111",
23058=>"111011100",
23059=>"000000000",
23060=>"111011001",
23061=>"000111111",
23062=>"111001100",
23063=>"111111110",
23064=>"101001110",
23065=>"010000000",
23066=>"001101011",
23067=>"000000101",
23068=>"000000000",
23069=>"111000000",
23070=>"010111111",
23071=>"000000000",
23072=>"000011000",
23073=>"100111111",
23074=>"110101101",
23075=>"000101101",
23076=>"111011001",
23077=>"001011000",
23078=>"000010010",
23079=>"001101111",
23080=>"011111111",
23081=>"001010010",
23082=>"101100110",
23083=>"110000000",
23084=>"000100011",
23085=>"111011100",
23086=>"111101110",
23087=>"000111000",
23088=>"001001000",
23089=>"011100101",
23090=>"001101101",
23091=>"000000000",
23092=>"000010010",
23093=>"110111110",
23094=>"011111110",
23095=>"010010010",
23096=>"111111100",
23097=>"000010000",
23098=>"000001100",
23099=>"000000000",
23100=>"001000000",
23101=>"100111111",
23102=>"110000010",
23103=>"000001100",
23104=>"111111000",
23105=>"010001001",
23106=>"101111111",
23107=>"001000000",
23108=>"111110000",
23109=>"000100111",
23110=>"000111111",
23111=>"111111111",
23112=>"101110000",
23113=>"011001101",
23114=>"000000111",
23115=>"010010010",
23116=>"111111010",
23117=>"010100010",
23118=>"011011111",
23119=>"000000011",
23120=>"000011111",
23121=>"100111011",
23122=>"000000110",
23123=>"111100000",
23124=>"000000001",
23125=>"111111111",
23126=>"000101110",
23127=>"000000010",
23128=>"111101100",
23129=>"000110000",
23130=>"000001101",
23131=>"111110000",
23132=>"000110000",
23133=>"110101000",
23134=>"101000000",
23135=>"000000100",
23136=>"010110010",
23137=>"000000000",
23138=>"011011011",
23139=>"111111111",
23140=>"000000100",
23141=>"000000000",
23142=>"000100111",
23143=>"000000111",
23144=>"100000000",
23145=>"111111101",
23146=>"010111111",
23147=>"000000100",
23148=>"100000111",
23149=>"101000101",
23150=>"000000000",
23151=>"000000101",
23152=>"011001011",
23153=>"010000101",
23154=>"111111011",
23155=>"001001001",
23156=>"111111111",
23157=>"000000000",
23158=>"001000000",
23159=>"010111011",
23160=>"101100111",
23161=>"111100000",
23162=>"111100100",
23163=>"111000100",
23164=>"000111111",
23165=>"111100000",
23166=>"101111011",
23167=>"000100000",
23168=>"111001000",
23169=>"000000000",
23170=>"101010000",
23171=>"111111111",
23172=>"000000000",
23173=>"111101000",
23174=>"101110000",
23175=>"000100000",
23176=>"000000000",
23177=>"000010000",
23178=>"000101111",
23179=>"111101101",
23180=>"010000000",
23181=>"101101100",
23182=>"111010000",
23183=>"000010010",
23184=>"001001001",
23185=>"000000000",
23186=>"000000000",
23187=>"000000101",
23188=>"100000000",
23189=>"000010010",
23190=>"111111100",
23191=>"000100001",
23192=>"001000000",
23193=>"000001000",
23194=>"010010010",
23195=>"111100011",
23196=>"000000111",
23197=>"010110110",
23198=>"001111111",
23199=>"000010000",
23200=>"101110000",
23201=>"000111111",
23202=>"101000000",
23203=>"111111010",
23204=>"011000000",
23205=>"011011011",
23206=>"111110100",
23207=>"001111111",
23208=>"001000101",
23209=>"000000101",
23210=>"011001101",
23211=>"000001000",
23212=>"111100000",
23213=>"000000111",
23214=>"001111111",
23215=>"100100101",
23216=>"110000001",
23217=>"000001001",
23218=>"111000000",
23219=>"000001100",
23220=>"101100111",
23221=>"101010000",
23222=>"010111111",
23223=>"100101101",
23224=>"000000000",
23225=>"000000000",
23226=>"000011111",
23227=>"111100111",
23228=>"000000101",
23229=>"111011011",
23230=>"110110000",
23231=>"011011111",
23232=>"001010010",
23233=>"000000000",
23234=>"111011111",
23235=>"100000010",
23236=>"110101101",
23237=>"111111111",
23238=>"010000011",
23239=>"111001000",
23240=>"111101111",
23241=>"000000000",
23242=>"111111101",
23243=>"001000000",
23244=>"000001000",
23245=>"000000111",
23246=>"010111010",
23247=>"110010101",
23248=>"000000000",
23249=>"011011001",
23250=>"110000101",
23251=>"111111111",
23252=>"000001111",
23253=>"000110100",
23254=>"000111011",
23255=>"000111001",
23256=>"111101111",
23257=>"000000111",
23258=>"101001000",
23259=>"101000101",
23260=>"111111001",
23261=>"100101111",
23262=>"010111011",
23263=>"111010111",
23264=>"000000111",
23265=>"111000110",
23266=>"110101001",
23267=>"001011000",
23268=>"000000000",
23269=>"101111101",
23270=>"100000000",
23271=>"100110110",
23272=>"000101111",
23273=>"000100000",
23274=>"110110010",
23275=>"011101111",
23276=>"000000111",
23277=>"110111111",
23278=>"000000000",
23279=>"110000000",
23280=>"000000000",
23281=>"011111110",
23282=>"111001101",
23283=>"001011000",
23284=>"101111011",
23285=>"101001000",
23286=>"001000011",
23287=>"110000011",
23288=>"111111000",
23289=>"111111111",
23290=>"100000000",
23291=>"000000110",
23292=>"111111000",
23293=>"101000000",
23294=>"110111011",
23295=>"101000010",
23296=>"100000010",
23297=>"000000000",
23298=>"100000100",
23299=>"011011111",
23300=>"110001001",
23301=>"101000011",
23302=>"110001010",
23303=>"000111000",
23304=>"100010000",
23305=>"110000010",
23306=>"010001011",
23307=>"010000100",
23308=>"110100000",
23309=>"011011000",
23310=>"010000000",
23311=>"000001000",
23312=>"000100000",
23313=>"000101111",
23314=>"101100001",
23315=>"111100110",
23316=>"100000000",
23317=>"001011111",
23318=>"111011001",
23319=>"111101011",
23320=>"000001110",
23321=>"111110110",
23322=>"001000000",
23323=>"111111110",
23324=>"110000000",
23325=>"001000000",
23326=>"111000000",
23327=>"000100000",
23328=>"001011110",
23329=>"001111100",
23330=>"000110101",
23331=>"011011011",
23332=>"110111110",
23333=>"111100100",
23334=>"000011110",
23335=>"111110001",
23336=>"110111100",
23337=>"110110011",
23338=>"100100100",
23339=>"110001010",
23340=>"110110110",
23341=>"000000000",
23342=>"110100110",
23343=>"111100101",
23344=>"111100110",
23345=>"110100010",
23346=>"000000000",
23347=>"111000000",
23348=>"010001110",
23349=>"000111011",
23350=>"111100000",
23351=>"011111110",
23352=>"100000011",
23353=>"001001000",
23354=>"000100010",
23355=>"111111111",
23356=>"111111111",
23357=>"010110001",
23358=>"000001001",
23359=>"001001011",
23360=>"110001000",
23361=>"110101010",
23362=>"110111111",
23363=>"000011011",
23364=>"111111111",
23365=>"000101100",
23366=>"010010011",
23367=>"101011111",
23368=>"000001011",
23369=>"011011010",
23370=>"000000000",
23371=>"010001100",
23372=>"100100010",
23373=>"011111111",
23374=>"001111000",
23375=>"001000001",
23376=>"011110100",
23377=>"111100101",
23378=>"110000000",
23379=>"000000011",
23380=>"111011000",
23381=>"011100001",
23382=>"110111110",
23383=>"001010001",
23384=>"110110111",
23385=>"110110100",
23386=>"001110110",
23387=>"100111100",
23388=>"100110001",
23389=>"000000000",
23390=>"111111111",
23391=>"010011101",
23392=>"011000001",
23393=>"000010001",
23394=>"110110010",
23395=>"000110100",
23396=>"000111100",
23397=>"111100010",
23398=>"111010010",
23399=>"000010110",
23400=>"000000010",
23401=>"011101001",
23402=>"010110110",
23403=>"000001001",
23404=>"100001111",
23405=>"000001001",
23406=>"011011011",
23407=>"000000000",
23408=>"110110110",
23409=>"000101111",
23410=>"000000111",
23411=>"100100100",
23412=>"011000011",
23413=>"100100110",
23414=>"001010010",
23415=>"111110000",
23416=>"000111111",
23417=>"010010100",
23418=>"000100100",
23419=>"101001101",
23420=>"001111111",
23421=>"110100001",
23422=>"110100100",
23423=>"011111001",
23424=>"111001000",
23425=>"110100100",
23426=>"111001011",
23427=>"000000011",
23428=>"001101001",
23429=>"101011101",
23430=>"000000000",
23431=>"000000000",
23432=>"110001001",
23433=>"000001101",
23434=>"100110101",
23435=>"101001100",
23436=>"100011111",
23437=>"001001011",
23438=>"111111111",
23439=>"101000100",
23440=>"010100000",
23441=>"100100000",
23442=>"100011010",
23443=>"000100000",
23444=>"000010000",
23445=>"000000001",
23446=>"011010110",
23447=>"100000000",
23448=>"011000101",
23449=>"101010010",
23450=>"011111110",
23451=>"000100110",
23452=>"111100001",
23453=>"000111111",
23454=>"010011001",
23455=>"100101101",
23456=>"100001000",
23457=>"110110001",
23458=>"011011000",
23459=>"010010100",
23460=>"011000010",
23461=>"011111111",
23462=>"111111010",
23463=>"111011001",
23464=>"011000000",
23465=>"000000110",
23466=>"001000000",
23467=>"101101000",
23468=>"011111110",
23469=>"010011010",
23470=>"111100000",
23471=>"001010110",
23472=>"000010000",
23473=>"111111001",
23474=>"011100000",
23475=>"000001111",
23476=>"001011111",
23477=>"000010010",
23478=>"110000011",
23479=>"000000000",
23480=>"000000000",
23481=>"111111111",
23482=>"111110100",
23483=>"100100111",
23484=>"001000000",
23485=>"001001111",
23486=>"000011000",
23487=>"000111110",
23488=>"000001000",
23489=>"001000011",
23490=>"001101111",
23491=>"110010100",
23492=>"000000001",
23493=>"000001011",
23494=>"110100011",
23495=>"111111111",
23496=>"101101110",
23497=>"110110100",
23498=>"101101100",
23499=>"100001110",
23500=>"000011100",
23501=>"000000000",
23502=>"101001000",
23503=>"111100100",
23504=>"000110110",
23505=>"111111101",
23506=>"000001000",
23507=>"100000001",
23508=>"011010000",
23509=>"001111001",
23510=>"100100001",
23511=>"110100011",
23512=>"110110000",
23513=>"000100100",
23514=>"000001111",
23515=>"000001101",
23516=>"110111000",
23517=>"000000110",
23518=>"001000100",
23519=>"011101001",
23520=>"000011011",
23521=>"100100100",
23522=>"000110110",
23523=>"100110110",
23524=>"000000011",
23525=>"111110110",
23526=>"101111100",
23527=>"000000110",
23528=>"011110100",
23529=>"001111111",
23530=>"001001010",
23531=>"111110110",
23532=>"011001000",
23533=>"101111001",
23534=>"101000000",
23535=>"011100111",
23536=>"110001011",
23537=>"110111110",
23538=>"011100100",
23539=>"110101011",
23540=>"111100000",
23541=>"001111101",
23542=>"000001011",
23543=>"000000100",
23544=>"000001001",
23545=>"011001011",
23546=>"000011011",
23547=>"000111110",
23548=>"110111011",
23549=>"000000110",
23550=>"100001000",
23551=>"011001010",
23552=>"000001100",
23553=>"111011000",
23554=>"000000111",
23555=>"011000000",
23556=>"110100100",
23557=>"000000111",
23558=>"110111001",
23559=>"100000100",
23560=>"000000000",
23561=>"000000000",
23562=>"011111000",
23563=>"001000111",
23564=>"110111000",
23565=>"111011001",
23566=>"001000000",
23567=>"110101000",
23568=>"100001001",
23569=>"000000111",
23570=>"111111011",
23571=>"111010000",
23572=>"010111110",
23573=>"101000000",
23574=>"000011000",
23575=>"111000000",
23576=>"111000001",
23577=>"110111001",
23578=>"000000001",
23579=>"000000110",
23580=>"111110011",
23581=>"111111001",
23582=>"111111111",
23583=>"001001101",
23584=>"000000000",
23585=>"101111111",
23586=>"100010010",
23587=>"100000000",
23588=>"101111001",
23589=>"100000010",
23590=>"000000011",
23591=>"000000011",
23592=>"000001111",
23593=>"111111110",
23594=>"000000011",
23595=>"111000000",
23596=>"011001010",
23597=>"010101101",
23598=>"111000111",
23599=>"011111011",
23600=>"000000000",
23601=>"100100110",
23602=>"111111111",
23603=>"110000110",
23604=>"000110000",
23605=>"111111111",
23606=>"101011011",
23607=>"101001000",
23608=>"111101000",
23609=>"111111111",
23610=>"000000000",
23611=>"000000010",
23612=>"000001001",
23613=>"111111111",
23614=>"000000000",
23615=>"110110010",
23616=>"111111110",
23617=>"100000110",
23618=>"011010000",
23619=>"001000000",
23620=>"111111111",
23621=>"110000000",
23622=>"010110010",
23623=>"110111101",
23624=>"001001001",
23625=>"000000000",
23626=>"101001011",
23627=>"111111110",
23628=>"001000110",
23629=>"101111100",
23630=>"001001011",
23631=>"000000010",
23632=>"000011101",
23633=>"101111111",
23634=>"000001000",
23635=>"001000000",
23636=>"111111110",
23637=>"101111100",
23638=>"110111011",
23639=>"001011111",
23640=>"001111111",
23641=>"000111110",
23642=>"101001000",
23643=>"011000000",
23644=>"010110100",
23645=>"001000000",
23646=>"111111111",
23647=>"001000000",
23648=>"010001110",
23649=>"011111111",
23650=>"000000111",
23651=>"000000000",
23652=>"000110100",
23653=>"111111111",
23654=>"001001001",
23655=>"000100000",
23656=>"111011111",
23657=>"001010111",
23658=>"101111111",
23659=>"000010101",
23660=>"111000100",
23661=>"010000101",
23662=>"011000000",
23663=>"111001110",
23664=>"000000000",
23665=>"111111011",
23666=>"111101111",
23667=>"010011000",
23668=>"000000000",
23669=>"101100110",
23670=>"110000001",
23671=>"111011100",
23672=>"000000000",
23673=>"000110101",
23674=>"000000000",
23675=>"010001000",
23676=>"100100011",
23677=>"000000000",
23678=>"000000000",
23679=>"000000000",
23680=>"010000110",
23681=>"000011010",
23682=>"000000111",
23683=>"000111101",
23684=>"111111100",
23685=>"100010010",
23686=>"001101001",
23687=>"011000110",
23688=>"001011000",
23689=>"011100000",
23690=>"011011000",
23691=>"010111111",
23692=>"111001000",
23693=>"000000011",
23694=>"000110111",
23695=>"111000001",
23696=>"101111111",
23697=>"000111101",
23698=>"010000000",
23699=>"001101000",
23700=>"011010101",
23701=>"000000000",
23702=>"110111111",
23703=>"011101100",
23704=>"111000111",
23705=>"000000001",
23706=>"000100010",
23707=>"000000000",
23708=>"111101001",
23709=>"101100111",
23710=>"101111111",
23711=>"000000000",
23712=>"000010001",
23713=>"000011111",
23714=>"010100000",
23715=>"000010101",
23716=>"111111111",
23717=>"110111011",
23718=>"110111110",
23719=>"001000001",
23720=>"111000111",
23721=>"111001001",
23722=>"000000110",
23723=>"101111111",
23724=>"111100000",
23725=>"001001111",
23726=>"001111011",
23727=>"000000110",
23728=>"000000001",
23729=>"100100101",
23730=>"000010111",
23731=>"001000010",
23732=>"011111000",
23733=>"110100100",
23734=>"011111110",
23735=>"010000000",
23736=>"001000100",
23737=>"111100001",
23738=>"110010111",
23739=>"010111111",
23740=>"111111101",
23741=>"111111111",
23742=>"001000110",
23743=>"000111111",
23744=>"110111000",
23745=>"000000100",
23746=>"111111110",
23747=>"000011100",
23748=>"110111111",
23749=>"000001000",
23750=>"111010100",
23751=>"100000000",
23752=>"000000000",
23753=>"101000000",
23754=>"110011111",
23755=>"111001010",
23756=>"101000000",
23757=>"011011100",
23758=>"111111111",
23759=>"000000111",
23760=>"111000001",
23761=>"100110110",
23762=>"110110110",
23763=>"111111011",
23764=>"000000111",
23765=>"111111001",
23766=>"101100000",
23767=>"110111001",
23768=>"000001000",
23769=>"000000000",
23770=>"000000000",
23771=>"000010111",
23772=>"001000011",
23773=>"110111101",
23774=>"111110111",
23775=>"111111101",
23776=>"001000011",
23777=>"000001011",
23778=>"000000000",
23779=>"000000000",
23780=>"000000000",
23781=>"000001000",
23782=>"000000000",
23783=>"001011010",
23784=>"000000010",
23785=>"111110001",
23786=>"110111111",
23787=>"110010000",
23788=>"001000010",
23789=>"111011000",
23790=>"000000000",
23791=>"000000101",
23792=>"101101111",
23793=>"001000011",
23794=>"111000101",
23795=>"101000000",
23796=>"100001011",
23797=>"000000001",
23798=>"010010111",
23799=>"000000100",
23800=>"000000000",
23801=>"101001000",
23802=>"110111111",
23803=>"111010000",
23804=>"111111011",
23805=>"010000111",
23806=>"101011011",
23807=>"000000000",
23808=>"011001001",
23809=>"000001110",
23810=>"001000001",
23811=>"000000001",
23812=>"011111111",
23813=>"000100110",
23814=>"000010010",
23815=>"111000000",
23816=>"000000000",
23817=>"010000010",
23818=>"111111111",
23819=>"000000000",
23820=>"000011011",
23821=>"010001001",
23822=>"011111001",
23823=>"000110011",
23824=>"001101000",
23825=>"000110000",
23826=>"110111100",
23827=>"111111111",
23828=>"111100100",
23829=>"111111111",
23830=>"111111111",
23831=>"000001000",
23832=>"000000000",
23833=>"111001101",
23834=>"000000101",
23835=>"010000000",
23836=>"111111111",
23837=>"001101111",
23838=>"111110010",
23839=>"000000000",
23840=>"000110000",
23841=>"111111111",
23842=>"001000000",
23843=>"000000000",
23844=>"011111000",
23845=>"110110010",
23846=>"000101111",
23847=>"000001101",
23848=>"110110000",
23849=>"111110110",
23850=>"001111000",
23851=>"111101010",
23852=>"111111111",
23853=>"100000000",
23854=>"000001000",
23855=>"011001111",
23856=>"000000000",
23857=>"011111000",
23858=>"000000000",
23859=>"111110010",
23860=>"111111111",
23861=>"111111111",
23862=>"110110101",
23863=>"101000010",
23864=>"111101111",
23865=>"000000000",
23866=>"000000001",
23867=>"010001000",
23868=>"001110000",
23869=>"111111111",
23870=>"001000100",
23871=>"101001100",
23872=>"011000111",
23873=>"011111011",
23874=>"111110000",
23875=>"001000100",
23876=>"111111111",
23877=>"000000000",
23878=>"010010010",
23879=>"111110010",
23880=>"000101001",
23881=>"000000000",
23882=>"000000001",
23883=>"001000001",
23884=>"001000001",
23885=>"111011000",
23886=>"110111110",
23887=>"110110110",
23888=>"111011100",
23889=>"110010100",
23890=>"000001111",
23891=>"001000111",
23892=>"000000001",
23893=>"111111101",
23894=>"111111000",
23895=>"001000001",
23896=>"010000000",
23897=>"111110111",
23898=>"111111111",
23899=>"111100111",
23900=>"111000000",
23901=>"001001001",
23902=>"110111010",
23903=>"100000000",
23904=>"001000000",
23905=>"000001001",
23906=>"111110010",
23907=>"000110011",
23908=>"000110100",
23909=>"111000000",
23910=>"000000001",
23911=>"000100100",
23912=>"001001111",
23913=>"011101000",
23914=>"111111110",
23915=>"000000111",
23916=>"011000100",
23917=>"010111000",
23918=>"001000010",
23919=>"010011000",
23920=>"110110111",
23921=>"011111110",
23922=>"011111111",
23923=>"000000101",
23924=>"000001111",
23925=>"100000100",
23926=>"111111111",
23927=>"100110110",
23928=>"000000000",
23929=>"111111000",
23930=>"111111100",
23931=>"000001001",
23932=>"111111111",
23933=>"100110101",
23934=>"011111111",
23935=>"001000001",
23936=>"001111111",
23937=>"111111111",
23938=>"010011010",
23939=>"111111110",
23940=>"001000110",
23941=>"111101000",
23942=>"100111100",
23943=>"000100000",
23944=>"011011001",
23945=>"010010001",
23946=>"000000000",
23947=>"000000000",
23948=>"000000000",
23949=>"110010111",
23950=>"001000011",
23951=>"000001000",
23952=>"101111001",
23953=>"000111111",
23954=>"000000111",
23955=>"000000110",
23956=>"011111110",
23957=>"000110011",
23958=>"110110000",
23959=>"000001000",
23960=>"111111111",
23961=>"000110111",
23962=>"010010010",
23963=>"100000010",
23964=>"000010011",
23965=>"000110010",
23966=>"000111010",
23967=>"001000001",
23968=>"001101000",
23969=>"010111101",
23970=>"000000101",
23971=>"000000000",
23972=>"001001111",
23973=>"000011011",
23974=>"101101001",
23975=>"011111101",
23976=>"110111111",
23977=>"100110100",
23978=>"000110100",
23979=>"011011111",
23980=>"011100000",
23981=>"100100110",
23982=>"100100101",
23983=>"111111010",
23984=>"000000000",
23985=>"011101000",
23986=>"000111011",
23987=>"001101000",
23988=>"001000100",
23989=>"111111111",
23990=>"011000000",
23991=>"010110000",
23992=>"110111011",
23993=>"011010011",
23994=>"101101010",
23995=>"000000000",
23996=>"000011000",
23997=>"111111010",
23998=>"100000000",
23999=>"000000000",
24000=>"000000000",
24001=>"011000011",
24002=>"000111111",
24003=>"011111111",
24004=>"000000000",
24005=>"110111110",
24006=>"010110110",
24007=>"111001111",
24008=>"000000000",
24009=>"000000100",
24010=>"001000000",
24011=>"111111111",
24012=>"001000000",
24013=>"111111111",
24014=>"111011111",
24015=>"110010011",
24016=>"000000110",
24017=>"100110000",
24018=>"000000000",
24019=>"001000011",
24020=>"000101111",
24021=>"000100000",
24022=>"000000000",
24023=>"111111111",
24024=>"000000100",
24025=>"010101101",
24026=>"111101100",
24027=>"000111111",
24028=>"111111110",
24029=>"000000001",
24030=>"100000011",
24031=>"110010000",
24032=>"010000010",
24033=>"000000000",
24034=>"000110000",
24035=>"010000000",
24036=>"000000100",
24037=>"001110111",
24038=>"001111111",
24039=>"111011001",
24040=>"101101110",
24041=>"000101111",
24042=>"111111111",
24043=>"101111111",
24044=>"000000000",
24045=>"100101000",
24046=>"110001010",
24047=>"000000000",
24048=>"111000010",
24049=>"111111111",
24050=>"001000010",
24051=>"001111111",
24052=>"100110100",
24053=>"111011101",
24054=>"000000111",
24055=>"101100101",
24056=>"000001000",
24057=>"111000111",
24058=>"010010000",
24059=>"000111011",
24060=>"110111111",
24061=>"111111111",
24062=>"110110010",
24063=>"101111101",
24064=>"001001110",
24065=>"011011010",
24066=>"111101101",
24067=>"011010100",
24068=>"000011111",
24069=>"101010011",
24070=>"000000010",
24071=>"000000000",
24072=>"000100010",
24073=>"111011000",
24074=>"001000100",
24075=>"100100000",
24076=>"101100011",
24077=>"001111101",
24078=>"110100000",
24079=>"100111000",
24080=>"010011011",
24081=>"100000100",
24082=>"100010000",
24083=>"000000010",
24084=>"111111001",
24085=>"011100111",
24086=>"111110111",
24087=>"111001011",
24088=>"100100110",
24089=>"000010011",
24090=>"000101100",
24091=>"111101000",
24092=>"100100100",
24093=>"100100001",
24094=>"111010000",
24095=>"000100111",
24096=>"001111111",
24097=>"011000000",
24098=>"111101101",
24099=>"000100011",
24100=>"000000110",
24101=>"110110111",
24102=>"000000111",
24103=>"000101101",
24104=>"010011011",
24105=>"000011111",
24106=>"010010111",
24107=>"001011001",
24108=>"000100000",
24109=>"001101011",
24110=>"111011111",
24111=>"000000000",
24112=>"000010010",
24113=>"000000001",
24114=>"011011101",
24115=>"101111100",
24116=>"100101000",
24117=>"101101000",
24118=>"000000001",
24119=>"000000000",
24120=>"000010010",
24121=>"011000101",
24122=>"111100100",
24123=>"001000111",
24124=>"011110110",
24125=>"111111011",
24126=>"000100100",
24127=>"001110010",
24128=>"111111000",
24129=>"011111101",
24130=>"111000000",
24131=>"001011010",
24132=>"011000000",
24133=>"000011011",
24134=>"000000010",
24135=>"111000000",
24136=>"000011011",
24137=>"011000000",
24138=>"000001111",
24139=>"010011011",
24140=>"111111011",
24141=>"001111111",
24142=>"000001100",
24143=>"111101000",
24144=>"000100111",
24145=>"111011000",
24146=>"011010011",
24147=>"011001000",
24148=>"111111100",
24149=>"001001001",
24150=>"111100111",
24151=>"111011000",
24152=>"101100110",
24153=>"000100101",
24154=>"011011101",
24155=>"001101100",
24156=>"010010010",
24157=>"000000001",
24158=>"011111001",
24159=>"100110010",
24160=>"000011111",
24161=>"011011111",
24162=>"100100110",
24163=>"110010010",
24164=>"000000010",
24165=>"110111101",
24166=>"111111000",
24167=>"010011101",
24168=>"100111111",
24169=>"011000100",
24170=>"101000000",
24171=>"100010111",
24172=>"000010011",
24173=>"000000000",
24174=>"001010000",
24175=>"010001000",
24176=>"000101001",
24177=>"000110000",
24178=>"000000010",
24179=>"100111111",
24180=>"110111100",
24181=>"000000100",
24182=>"111111011",
24183=>"000101101",
24184=>"111000100",
24185=>"111000110",
24186=>"000001111",
24187=>"000000001",
24188=>"110110110",
24189=>"110100000",
24190=>"011011011",
24191=>"100100101",
24192=>"011010100",
24193=>"011100000",
24194=>"001000000",
24195=>"100000011",
24196=>"101100010",
24197=>"000111111",
24198=>"011011011",
24199=>"000001111",
24200=>"000110111",
24201=>"011010001",
24202=>"011000100",
24203=>"000110101",
24204=>"000000100",
24205=>"101101111",
24206=>"100100100",
24207=>"000000001",
24208=>"001101101",
24209=>"111111110",
24210=>"000000100",
24211=>"101000000",
24212=>"000000000",
24213=>"111011000",
24214=>"110000000",
24215=>"010100011",
24216=>"111101100",
24217=>"010001000",
24218=>"100111111",
24219=>"000000000",
24220=>"111110000",
24221=>"111011111",
24222=>"011101100",
24223=>"000000000",
24224=>"100001010",
24225=>"100101111",
24226=>"000000111",
24227=>"111000011",
24228=>"100100111",
24229=>"000111011",
24230=>"111010111",
24231=>"001111111",
24232=>"111000111",
24233=>"101001111",
24234=>"101000000",
24235=>"000010110",
24236=>"111000100",
24237=>"101000100",
24238=>"001001000",
24239=>"011011011",
24240=>"000011000",
24241=>"100111011",
24242=>"000001011",
24243=>"000001100",
24244=>"100100111",
24245=>"110111011",
24246=>"101000111",
24247=>"111011101",
24248=>"110001011",
24249=>"000100011",
24250=>"000111111",
24251=>"111000000",
24252=>"011111000",
24253=>"111111111",
24254=>"000001001",
24255=>"000111111",
24256=>"100010010",
24257=>"000000000",
24258=>"011011011",
24259=>"000000111",
24260=>"000000001",
24261=>"110000000",
24262=>"010010011",
24263=>"101000100",
24264=>"000100000",
24265=>"000000011",
24266=>"100011011",
24267=>"100110110",
24268=>"000011011",
24269=>"011000001",
24270=>"111110000",
24271=>"111111101",
24272=>"011000101",
24273=>"001001110",
24274=>"000100111",
24275=>"100100100",
24276=>"100111101",
24277=>"000100110",
24278=>"111000000",
24279=>"011010000",
24280=>"000111000",
24281=>"100111000",
24282=>"001000100",
24283=>"111000000",
24284=>"001001110",
24285=>"000001001",
24286=>"100000000",
24287=>"111011000",
24288=>"000000001",
24289=>"001001001",
24290=>"101000111",
24291=>"001001001",
24292=>"000011111",
24293=>"000010111",
24294=>"000010011",
24295=>"100100100",
24296=>"011101000",
24297=>"111000101",
24298=>"110000001",
24299=>"111111100",
24300=>"010011010",
24301=>"100100000",
24302=>"111000000",
24303=>"000000010",
24304=>"000000000",
24305=>"000100000",
24306=>"111111101",
24307=>"001101100",
24308=>"100110101",
24309=>"111000000",
24310=>"000000000",
24311=>"000100000",
24312=>"000000110",
24313=>"111111000",
24314=>"111101101",
24315=>"100000111",
24316=>"111000000",
24317=>"001111111",
24318=>"110100111",
24319=>"101011010",
24320=>"100011100",
24321=>"001000001",
24322=>"011010010",
24323=>"111101111",
24324=>"011111111",
24325=>"110101110",
24326=>"000000111",
24327=>"000000011",
24328=>"110100000",
24329=>"110110011",
24330=>"111000000",
24331=>"111011111",
24332=>"111111001",
24333=>"100000000",
24334=>"101011011",
24335=>"100011010",
24336=>"011111100",
24337=>"001111110",
24338=>"111101100",
24339=>"000000101",
24340=>"010011000",
24341=>"101100100",
24342=>"000000011",
24343=>"110111110",
24344=>"000100001",
24345=>"101101011",
24346=>"011100111",
24347=>"100000111",
24348=>"111110111",
24349=>"000100001",
24350=>"011110110",
24351=>"001001000",
24352=>"011111000",
24353=>"010111100",
24354=>"111000001",
24355=>"111000110",
24356=>"010111001",
24357=>"000100000",
24358=>"000000000",
24359=>"110001111",
24360=>"001101000",
24361=>"110100000",
24362=>"010010110",
24363=>"011111011",
24364=>"100111001",
24365=>"100000000",
24366=>"011111000",
24367=>"000000001",
24368=>"111011011",
24369=>"000001001",
24370=>"011111110",
24371=>"010110110",
24372=>"001001001",
24373=>"111110110",
24374=>"011001011",
24375=>"100000100",
24376=>"010111010",
24377=>"100000110",
24378=>"111000000",
24379=>"111001011",
24380=>"000110000",
24381=>"001001000",
24382=>"110100000",
24383=>"001011010",
24384=>"101011000",
24385=>"001000000",
24386=>"101011000",
24387=>"000011100",
24388=>"111000011",
24389=>"000111111",
24390=>"110000001",
24391=>"011111011",
24392=>"111110000",
24393=>"111110000",
24394=>"010100100",
24395=>"001001101",
24396=>"000100101",
24397=>"001011011",
24398=>"010001000",
24399=>"110001011",
24400=>"001000000",
24401=>"100111111",
24402=>"111100010",
24403=>"111000000",
24404=>"001000000",
24405=>"011000001",
24406=>"101001001",
24407=>"111110100",
24408=>"111100101",
24409=>"001011011",
24410=>"001000001",
24411=>"000001110",
24412=>"111111111",
24413=>"100000101",
24414=>"110111010",
24415=>"001011000",
24416=>"111111011",
24417=>"011001000",
24418=>"011110011",
24419=>"000000000",
24420=>"110000000",
24421=>"001111000",
24422=>"001100001",
24423=>"101000000",
24424=>"001101000",
24425=>"000010010",
24426=>"010010111",
24427=>"100100111",
24428=>"111011111",
24429=>"100100110",
24430=>"110100000",
24431=>"110000011",
24432=>"001011011",
24433=>"011111110",
24434=>"111000001",
24435=>"011000000",
24436=>"111001111",
24437=>"100100101",
24438=>"000100110",
24439=>"111000100",
24440=>"011110000",
24441=>"110001110",
24442=>"000001111",
24443=>"100100000",
24444=>"000000001",
24445=>"110000000",
24446=>"111000100",
24447=>"011000000",
24448=>"000110110",
24449=>"111000100",
24450=>"110000001",
24451=>"011000001",
24452=>"110100001",
24453=>"110100111",
24454=>"010111000",
24455=>"000001010",
24456=>"001001001",
24457=>"011000000",
24458=>"000000100",
24459=>"101100110",
24460=>"111110100",
24461=>"101100011",
24462=>"110000001",
24463=>"011011000",
24464=>"010011011",
24465=>"011110000",
24466=>"001001000",
24467=>"001001001",
24468=>"001011111",
24469=>"000110110",
24470=>"000011010",
24471=>"111011011",
24472=>"100100111",
24473=>"111110011",
24474=>"011110011",
24475=>"100000000",
24476=>"000100100",
24477=>"111110101",
24478=>"010000110",
24479=>"001100101",
24480=>"110100000",
24481=>"111110100",
24482=>"111001000",
24483=>"111010100",
24484=>"110000111",
24485=>"011001001",
24486=>"110101001",
24487=>"001111111",
24488=>"100010110",
24489=>"001001111",
24490=>"111000000",
24491=>"110000001",
24492=>"000010101",
24493=>"011000001",
24494=>"011100100",
24495=>"111110000",
24496=>"010110000",
24497=>"100111111",
24498=>"110000011",
24499=>"000000000",
24500=>"111111001",
24501=>"001100100",
24502=>"011011111",
24503=>"000000001",
24504=>"100100110",
24505=>"010000000",
24506=>"111110100",
24507=>"000011011",
24508=>"000000111",
24509=>"111111111",
24510=>"111001000",
24511=>"011011110",
24512=>"110110000",
24513=>"010000000",
24514=>"000001011",
24515=>"000011100",
24516=>"000000000",
24517=>"010000101",
24518=>"100011001",
24519=>"111100100",
24520=>"001000011",
24521=>"000000010",
24522=>"001010000",
24523=>"011010111",
24524=>"000111000",
24525=>"001001001",
24526=>"000001100",
24527=>"111111111",
24528=>"011111110",
24529=>"000001011",
24530=>"011100000",
24531=>"111101000",
24532=>"010010001",
24533=>"000000000",
24534=>"110111111",
24535=>"010011111",
24536=>"111111001",
24537=>"010010000",
24538=>"001001001",
24539=>"111100100",
24540=>"001011011",
24541=>"101101101",
24542=>"000010000",
24543=>"001011110",
24544=>"110111011",
24545=>"000010011",
24546=>"111100110",
24547=>"111110110",
24548=>"000110100",
24549=>"010100111",
24550=>"001111000",
24551=>"100100110",
24552=>"110111111",
24553=>"101110000",
24554=>"110111010",
24555=>"111111110",
24556=>"001100000",
24557=>"001011111",
24558=>"000111100",
24559=>"110000110",
24560=>"111001001",
24561=>"100101111",
24562=>"110000010",
24563=>"101011000",
24564=>"001101001",
24565=>"110000000",
24566=>"000100110",
24567=>"000000111",
24568=>"011111110",
24569=>"110111100",
24570=>"110111101",
24571=>"100001001",
24572=>"000001001",
24573=>"100010110",
24574=>"110000001",
24575=>"001001011",
24576=>"100100111",
24577=>"010010010",
24578=>"101111111",
24579=>"000000000",
24580=>"000100100",
24581=>"000111111",
24582=>"100100100",
24583=>"011111111",
24584=>"101101101",
24585=>"000000000",
24586=>"111100100",
24587=>"110000000",
24588=>"000100111",
24589=>"000000111",
24590=>"011000000",
24591=>"111111111",
24592=>"000000000",
24593=>"000000101",
24594=>"001000000",
24595=>"011011000",
24596=>"111011111",
24597=>"110000000",
24598=>"111111011",
24599=>"011000000",
24600=>"100000000",
24601=>"111111111",
24602=>"000000000",
24603=>"000000100",
24604=>"111101111",
24605=>"000000000",
24606=>"000000111",
24607=>"010010000",
24608=>"010110010",
24609=>"000010000",
24610=>"000000000",
24611=>"100110011",
24612=>"110011001",
24613=>"111001011",
24614=>"111000000",
24615=>"111110101",
24616=>"010111011",
24617=>"011101100",
24618=>"111111000",
24619=>"000001000",
24620=>"111001000",
24621=>"110011010",
24622=>"100000000",
24623=>"010111111",
24624=>"110111010",
24625=>"001000000",
24626=>"011100001",
24627=>"110000000",
24628=>"111100110",
24629=>"110000000",
24630=>"011000000",
24631=>"011000010",
24632=>"000110111",
24633=>"011101100",
24634=>"110011100",
24635=>"100110110",
24636=>"010011011",
24637=>"011000111",
24638=>"000011111",
24639=>"000000100",
24640=>"011111101",
24641=>"110101111",
24642=>"100000001",
24643=>"101101111",
24644=>"111111111",
24645=>"000000000",
24646=>"111101111",
24647=>"011110011",
24648=>"110011111",
24649=>"000010010",
24650=>"000010000",
24651=>"101100101",
24652=>"100110111",
24653=>"011111111",
24654=>"100110010",
24655=>"111000000",
24656=>"110000000",
24657=>"111111010",
24658=>"111110111",
24659=>"110110100",
24660=>"010100100",
24661=>"110101001",
24662=>"111111000",
24663=>"111001111",
24664=>"101111101",
24665=>"111001010",
24666=>"000001000",
24667=>"110000100",
24668=>"100000000",
24669=>"011011011",
24670=>"101100101",
24671=>"001001111",
24672=>"000100100",
24673=>"010010010",
24674=>"000000000",
24675=>"100100000",
24676=>"111111111",
24677=>"101111011",
24678=>"010010110",
24679=>"011110000",
24680=>"000000000",
24681=>"011011111",
24682=>"010111101",
24683=>"111101101",
24684=>"001100000",
24685=>"010111001",
24686=>"000111110",
24687=>"111111101",
24688=>"110110110",
24689=>"000000000",
24690=>"001000000",
24691=>"101000000",
24692=>"000110000",
24693=>"000011010",
24694=>"000000000",
24695=>"100111111",
24696=>"000000000",
24697=>"011000000",
24698=>"111111010",
24699=>"000100011",
24700=>"111011001",
24701=>"011011011",
24702=>"000101000",
24703=>"101000011",
24704=>"000010110",
24705=>"011111000",
24706=>"000000000",
24707=>"011011101",
24708=>"000000000",
24709=>"111101000",
24710=>"110100110",
24711=>"111110110",
24712=>"011011011",
24713=>"111101111",
24714=>"000000000",
24715=>"101101000",
24716=>"111111111",
24717=>"011010010",
24718=>"000000000",
24719=>"101000100",
24720=>"110110110",
24721=>"001000000",
24722=>"100101000",
24723=>"011101110",
24724=>"000100000",
24725=>"010111111",
24726=>"111100000",
24727=>"001110010",
24728=>"111101100",
24729=>"010111101",
24730=>"000000000",
24731=>"000011000",
24732=>"010100100",
24733=>"000000000",
24734=>"010111111",
24735=>"110000000",
24736=>"111110111",
24737=>"000011000",
24738=>"111111000",
24739=>"011011000",
24740=>"000001110",
24741=>"011011011",
24742=>"000010010",
24743=>"000000000",
24744=>"100110000",
24745=>"111101000",
24746=>"000010111",
24747=>"110111111",
24748=>"110010010",
24749=>"010111111",
24750=>"011001001",
24751=>"001000111",
24752=>"100001111",
24753=>"110110111",
24754=>"000000000",
24755=>"010011000",
24756=>"111110000",
24757=>"001000001",
24758=>"001111000",
24759=>"111001110",
24760=>"110110010",
24761=>"011001001",
24762=>"110000000",
24763=>"000110111",
24764=>"000100100",
24765=>"111111111",
24766=>"110100000",
24767=>"000000110",
24768=>"111011011",
24769=>"000010000",
24770=>"000101110",
24771=>"110011011",
24772=>"101000000",
24773=>"011111110",
24774=>"000010000",
24775=>"100000100",
24776=>"111111111",
24777=>"101101111",
24778=>"000011000",
24779=>"110100101",
24780=>"110000000",
24781=>"110110000",
24782=>"111111100",
24783=>"000000000",
24784=>"010100000",
24785=>"110110110",
24786=>"010000000",
24787=>"010100000",
24788=>"000011111",
24789=>"111111110",
24790=>"101101000",
24791=>"001010000",
24792=>"000000000",
24793=>"000000000",
24794=>"111111101",
24795=>"110110000",
24796=>"101011110",
24797=>"010000000",
24798=>"100100000",
24799=>"000000101",
24800=>"000000000",
24801=>"000011010",
24802=>"000000000",
24803=>"111010011",
24804=>"111000000",
24805=>"111100100",
24806=>"110000100",
24807=>"110010000",
24808=>"110111111",
24809=>"110100000",
24810=>"111000000",
24811=>"111101101",
24812=>"000000010",
24813=>"110000000",
24814=>"000111010",
24815=>"000111010",
24816=>"010000000",
24817=>"110101111",
24818=>"000101111",
24819=>"110000000",
24820=>"100000011",
24821=>"100100000",
24822=>"111111111",
24823=>"100100000",
24824=>"000111101",
24825=>"111111100",
24826=>"111111110",
24827=>"010110000",
24828=>"101101101",
24829=>"010010111",
24830=>"111111111",
24831=>"000000000",
24832=>"010100100",
24833=>"011111111",
24834=>"000010111",
24835=>"111111101",
24836=>"010010111",
24837=>"010011011",
24838=>"000000000",
24839=>"000111000",
24840=>"010100000",
24841=>"000000101",
24842=>"001100100",
24843=>"010101101",
24844=>"000000000",
24845=>"110100000",
24846=>"110000000",
24847=>"100000000",
24848=>"110111101",
24849=>"000111101",
24850=>"110111110",
24851=>"000100111",
24852=>"101000010",
24853=>"010011001",
24854=>"010110111",
24855=>"111111000",
24856=>"000000000",
24857=>"000000001",
24858=>"000000111",
24859=>"000111111",
24860=>"011111001",
24861=>"111110101",
24862=>"010111111",
24863=>"000000111",
24864=>"111000101",
24865=>"000001110",
24866=>"000001100",
24867=>"000111111",
24868=>"110110110",
24869=>"110000000",
24870=>"000010100",
24871=>"011011101",
24872=>"111110010",
24873=>"010000000",
24874=>"110000000",
24875=>"111000100",
24876=>"110111000",
24877=>"111101101",
24878=>"110111101",
24879=>"110001000",
24880=>"100000100",
24881=>"011111110",
24882=>"000000000",
24883=>"011101001",
24884=>"110110000",
24885=>"111111101",
24886=>"111100000",
24887=>"111101111",
24888=>"001000011",
24889=>"000000111",
24890=>"111101000",
24891=>"000000010",
24892=>"011001001",
24893=>"111111111",
24894=>"101000100",
24895=>"111011111",
24896=>"111100000",
24897=>"010000010",
24898=>"011001000",
24899=>"110110110",
24900=>"110001110",
24901=>"000101101",
24902=>"000100000",
24903=>"101101101",
24904=>"111010000",
24905=>"000000101",
24906=>"000000000",
24907=>"000000000",
24908=>"111000100",
24909=>"111010011",
24910=>"110110011",
24911=>"011111010",
24912=>"101001000",
24913=>"111111110",
24914=>"111111101",
24915=>"111011000",
24916=>"010111010",
24917=>"011110111",
24918=>"000110011",
24919=>"000010010",
24920=>"011111111",
24921=>"001001101",
24922=>"110101100",
24923=>"110010000",
24924=>"000000101",
24925=>"001001100",
24926=>"111111010",
24927=>"110111110",
24928=>"000001111",
24929=>"000111011",
24930=>"101000000",
24931=>"110110001",
24932=>"010000001",
24933=>"000100000",
24934=>"010111000",
24935=>"111010000",
24936=>"000111111",
24937=>"100000111",
24938=>"000011111",
24939=>"111011000",
24940=>"111110100",
24941=>"101111100",
24942=>"100000000",
24943=>"101101000",
24944=>"000000110",
24945=>"000000010",
24946=>"001000000",
24947=>"100000000",
24948=>"010111111",
24949=>"000101111",
24950=>"000000010",
24951=>"100100000",
24952=>"000111111",
24953=>"000111110",
24954=>"101000101",
24955=>"110000101",
24956=>"111111000",
24957=>"110001011",
24958=>"111000001",
24959=>"000111101",
24960=>"010011011",
24961=>"111101100",
24962=>"111000001",
24963=>"101111110",
24964=>"010111111",
24965=>"011001001",
24966=>"010001110",
24967=>"010000100",
24968=>"010000001",
24969=>"110000101",
24970=>"000011011",
24971=>"000100111",
24972=>"101000101",
24973=>"101000101",
24974=>"100101000",
24975=>"000000000",
24976=>"111011001",
24977=>"011001111",
24978=>"101001100",
24979=>"000111000",
24980=>"110011100",
24981=>"000000111",
24982=>"110000111",
24983=>"100100100",
24984=>"100101001",
24985=>"011111111",
24986=>"111000000",
24987=>"000110000",
24988=>"010101000",
24989=>"110100000",
24990=>"000010111",
24991=>"100000001",
24992=>"111010010",
24993=>"000110110",
24994=>"000001000",
24995=>"000000000",
24996=>"110001101",
24997=>"101110111",
24998=>"001000110",
24999=>"111111101",
25000=>"101011011",
25001=>"100101101",
25002=>"000000101",
25003=>"111000000",
25004=>"100101101",
25005=>"001000100",
25006=>"011000100",
25007=>"010000010",
25008=>"110111010",
25009=>"110100101",
25010=>"000001011",
25011=>"000000000",
25012=>"000011011",
25013=>"000000000",
25014=>"110010110",
25015=>"010000001",
25016=>"110110000",
25017=>"000010011",
25018=>"000000000",
25019=>"001000101",
25020=>"011000010",
25021=>"101000101",
25022=>"100100100",
25023=>"000000000",
25024=>"000010110",
25025=>"000000001",
25026=>"011000000",
25027=>"011000101",
25028=>"110000000",
25029=>"111100000",
25030=>"000011100",
25031=>"010011010",
25032=>"110111000",
25033=>"001111111",
25034=>"110001111",
25035=>"111110110",
25036=>"000011010",
25037=>"011110000",
25038=>"101001100",
25039=>"100000010",
25040=>"111111111",
25041=>"010011110",
25042=>"010111011",
25043=>"101100110",
25044=>"011011000",
25045=>"000001001",
25046=>"010011111",
25047=>"100001111",
25048=>"010011010",
25049=>"100000000",
25050=>"011010000",
25051=>"101000000",
25052=>"111111111",
25053=>"010111100",
25054=>"000000000",
25055=>"100101111",
25056=>"010011010",
25057=>"100000110",
25058=>"000111111",
25059=>"011010000",
25060=>"000010010",
25061=>"011111000",
25062=>"111001000",
25063=>"100111011",
25064=>"111111111",
25065=>"000000000",
25066=>"010000000",
25067=>"111101111",
25068=>"000000000",
25069=>"000000010",
25070=>"000000100",
25071=>"010111111",
25072=>"010100101",
25073=>"111000000",
25074=>"010000000",
25075=>"010110100",
25076=>"001001001",
25077=>"101110101",
25078=>"111001001",
25079=>"111111100",
25080=>"111000000",
25081=>"001000000",
25082=>"011111111",
25083=>"000000101",
25084=>"010010111",
25085=>"111111111",
25086=>"010010100",
25087=>"000101000",
25088=>"010010000",
25089=>"100110010",
25090=>"100111000",
25091=>"000101110",
25092=>"100011011",
25093=>"110000000",
25094=>"111111111",
25095=>"010000010",
25096=>"000000000",
25097=>"111111000",
25098=>"110110100",
25099=>"101101111",
25100=>"100111111",
25101=>"110011111",
25102=>"100010011",
25103=>"110100000",
25104=>"110001101",
25105=>"000000001",
25106=>"000000000",
25107=>"111001000",
25108=>"000000000",
25109=>"011010000",
25110=>"011000000",
25111=>"010111011",
25112=>"100000011",
25113=>"111111111",
25114=>"010000111",
25115=>"000000000",
25116=>"100110111",
25117=>"000000101",
25118=>"111000000",
25119=>"001111111",
25120=>"111101101",
25121=>"100111111",
25122=>"000110111",
25123=>"010000000",
25124=>"000001101",
25125=>"001010101",
25126=>"010010010",
25127=>"000001001",
25128=>"111000000",
25129=>"111101111",
25130=>"010010000",
25131=>"101111111",
25132=>"011000011",
25133=>"001000000",
25134=>"111111011",
25135=>"000000000",
25136=>"000101111",
25137=>"111111011",
25138=>"000001001",
25139=>"000000000",
25140=>"000000000",
25141=>"101110000",
25142=>"010001011",
25143=>"000000000",
25144=>"000000010",
25145=>"000000000",
25146=>"010000000",
25147=>"001101101",
25148=>"000000000",
25149=>"011111111",
25150=>"100100101",
25151=>"110110110",
25152=>"111111011",
25153=>"001001010",
25154=>"110110000",
25155=>"011000000",
25156=>"000111111",
25157=>"000001111",
25158=>"111111000",
25159=>"010001000",
25160=>"100000101",
25161=>"011001111",
25162=>"000001000",
25163=>"000001001",
25164=>"000001001",
25165=>"000001110",
25166=>"110110100",
25167=>"111011111",
25168=>"000111000",
25169=>"111111111",
25170=>"101110000",
25171=>"111011100",
25172=>"111010000",
25173=>"001000101",
25174=>"001001000",
25175=>"000000000",
25176=>"011110110",
25177=>"111001001",
25178=>"011011010",
25179=>"101000100",
25180=>"000001111",
25181=>"010001001",
25182=>"000101111",
25183=>"000000001",
25184=>"111111011",
25185=>"001001010",
25186=>"001011010",
25187=>"100000000",
25188=>"111100000",
25189=>"111111000",
25190=>"000100010",
25191=>"110010000",
25192=>"111111111",
25193=>"000000011",
25194=>"010000111",
25195=>"100111001",
25196=>"000100111",
25197=>"010111101",
25198=>"010110000",
25199=>"010000001",
25200=>"111011111",
25201=>"000000010",
25202=>"110100110",
25203=>"111111010",
25204=>"110110111",
25205=>"000000000",
25206=>"000000110",
25207=>"000000000",
25208=>"100000000",
25209=>"111101111",
25210=>"111011001",
25211=>"010000000",
25212=>"001100000",
25213=>"000000000",
25214=>"110011111",
25215=>"000000000",
25216=>"110111101",
25217=>"110100000",
25218=>"000000111",
25219=>"000000000",
25220=>"111100000",
25221=>"011000101",
25222=>"100100100",
25223=>"100101011",
25224=>"111101001",
25225=>"000001000",
25226=>"010101010",
25227=>"101000001",
25228=>"000001001",
25229=>"000101111",
25230=>"000000111",
25231=>"101000000",
25232=>"000101100",
25233=>"110110111",
25234=>"000000111",
25235=>"111000001",
25236=>"100111111",
25237=>"001000000",
25238=>"000000111",
25239=>"011001011",
25240=>"101101111",
25241=>"000000001",
25242=>"100110111",
25243=>"111000000",
25244=>"001000001",
25245=>"100001101",
25246=>"111111101",
25247=>"001001000",
25248=>"111101101",
25249=>"010000101",
25250=>"000101101",
25251=>"111100000",
25252=>"110000111",
25253=>"111110000",
25254=>"001001000",
25255=>"010000001",
25256=>"111100000",
25257=>"000010000",
25258=>"010010000",
25259=>"000000010",
25260=>"000000000",
25261=>"001000000",
25262=>"110001000",
25263=>"111111010",
25264=>"001100111",
25265=>"110111111",
25266=>"000000101",
25267=>"000110100",
25268=>"111111111",
25269=>"000000000",
25270=>"101111011",
25271=>"101111101",
25272=>"000000000",
25273=>"000110110",
25274=>"110000010",
25275=>"110110100",
25276=>"101101101",
25277=>"010001111",
25278=>"001001110",
25279=>"111111111",
25280=>"000111001",
25281=>"000111111",
25282=>"111010001",
25283=>"001000000",
25284=>"000000000",
25285=>"100100001",
25286=>"110010011",
25287=>"010010010",
25288=>"001000111",
25289=>"001111000",
25290=>"111110111",
25291=>"000001111",
25292=>"111000001",
25293=>"100111110",
25294=>"111010001",
25295=>"111101111",
25296=>"000001111",
25297=>"110010010",
25298=>"111001011",
25299=>"001110111",
25300=>"110101001",
25301=>"111110001",
25302=>"011000000",
25303=>"110010101",
25304=>"000000000",
25305=>"101001010",
25306=>"111111101",
25307=>"000111010",
25308=>"100001000",
25309=>"011111000",
25310=>"111111110",
25311=>"011111000",
25312=>"000010110",
25313=>"000000101",
25314=>"000110111",
25315=>"110100000",
25316=>"010000000",
25317=>"101111110",
25318=>"011010111",
25319=>"000100100",
25320=>"100111111",
25321=>"000101111",
25322=>"001000011",
25323=>"010111010",
25324=>"111110000",
25325=>"011111111",
25326=>"000110000",
25327=>"000000110",
25328=>"110010000",
25329=>"001001001",
25330=>"110110000",
25331=>"110100110",
25332=>"001000110",
25333=>"111111000",
25334=>"000010001",
25335=>"100110000",
25336=>"000100101",
25337=>"000001000",
25338=>"111010111",
25339=>"000101000",
25340=>"000000111",
25341=>"011111111",
25342=>"111000000",
25343=>"000000000",
25344=>"000110110",
25345=>"110100000",
25346=>"001000100",
25347=>"101100000",
25348=>"111111111",
25349=>"111111000",
25350=>"000011011",
25351=>"000000000",
25352=>"100000001",
25353=>"101000100",
25354=>"111111111",
25355=>"010101100",
25356=>"111110100",
25357=>"111110000",
25358=>"110110100",
25359=>"000000000",
25360=>"100111111",
25361=>"111111111",
25362=>"000011111",
25363=>"110010000",
25364=>"100010010",
25365=>"111111111",
25366=>"000000001",
25367=>"111111111",
25368=>"101010011",
25369=>"000000110",
25370=>"111110000",
25371=>"010100010",
25372=>"000000001",
25373=>"001000000",
25374=>"000001111",
25375=>"000010000",
25376=>"001000000",
25377=>"000010000",
25378=>"000011100",
25379=>"010000010",
25380=>"001010111",
25381=>"011011011",
25382=>"000110010",
25383=>"000000101",
25384=>"000000100",
25385=>"010100111",
25386=>"010011011",
25387=>"000010000",
25388=>"011111110",
25389=>"111010000",
25390=>"111110011",
25391=>"000000000",
25392=>"000000000",
25393=>"000110110",
25394=>"011000000",
25395=>"010111101",
25396=>"111101111",
25397=>"111101010",
25398=>"001001000",
25399=>"010011101",
25400=>"111110110",
25401=>"111010000",
25402=>"001000000",
25403=>"000000000",
25404=>"001100001",
25405=>"111011111",
25406=>"000100000",
25407=>"011011011",
25408=>"110000111",
25409=>"101000111",
25410=>"111000000",
25411=>"010001001",
25412=>"111111110",
25413=>"000000000",
25414=>"000000001",
25415=>"101101001",
25416=>"110000010",
25417=>"000111111",
25418=>"100100101",
25419=>"011101111",
25420=>"001101111",
25421=>"100010110",
25422=>"001111111",
25423=>"011111111",
25424=>"111100000",
25425=>"100101111",
25426=>"000010000",
25427=>"000110000",
25428=>"011000100",
25429=>"010011001",
25430=>"000110011",
25431=>"000000101",
25432=>"111111101",
25433=>"011011011",
25434=>"011010000",
25435=>"100111111",
25436=>"000101101",
25437=>"001100100",
25438=>"000011010",
25439=>"110101001",
25440=>"111101000",
25441=>"010000100",
25442=>"000000110",
25443=>"001011010",
25444=>"011011011",
25445=>"010100001",
25446=>"000000111",
25447=>"011111111",
25448=>"000000000",
25449=>"111011111",
25450=>"110010001",
25451=>"000111100",
25452=>"010011111",
25453=>"101111010",
25454=>"000000000",
25455=>"111111111",
25456=>"111011110",
25457=>"111111111",
25458=>"001000000",
25459=>"000110100",
25460=>"010111101",
25461=>"000000000",
25462=>"111111101",
25463=>"001000000",
25464=>"101000000",
25465=>"111111111",
25466=>"000101111",
25467=>"111111101",
25468=>"000000000",
25469=>"001001001",
25470=>"001000100",
25471=>"101100110",
25472=>"000010010",
25473=>"000010000",
25474=>"101100100",
25475=>"000111111",
25476=>"000010000",
25477=>"101000101",
25478=>"101100001",
25479=>"100000110",
25480=>"100110111",
25481=>"101101011",
25482=>"111111110",
25483=>"000101111",
25484=>"111111100",
25485=>"000101111",
25486=>"100111111",
25487=>"000000001",
25488=>"001011011",
25489=>"111111100",
25490=>"101101111",
25491=>"100100100",
25492=>"000100110",
25493=>"101101111",
25494=>"111111111",
25495=>"110110110",
25496=>"010011111",
25497=>"100000000",
25498=>"101100101",
25499=>"000000000",
25500=>"110110111",
25501=>"000000000",
25502=>"100111111",
25503=>"111111111",
25504=>"011000111",
25505=>"001111111",
25506=>"111101111",
25507=>"111010111",
25508=>"000010000",
25509=>"011011011",
25510=>"000000001",
25511=>"011111111",
25512=>"100001000",
25513=>"101000000",
25514=>"001000000",
25515=>"000110000",
25516=>"100010000",
25517=>"000111111",
25518=>"000101111",
25519=>"111000001",
25520=>"100000100",
25521=>"100110110",
25522=>"000000000",
25523=>"011011001",
25524=>"010111111",
25525=>"001100000",
25526=>"011110000",
25527=>"100111101",
25528=>"100101000",
25529=>"001001001",
25530=>"001100101",
25531=>"010000111",
25532=>"101111111",
25533=>"101001001",
25534=>"100100100",
25535=>"111110010",
25536=>"000000010",
25537=>"101000000",
25538=>"110011001",
25539=>"000000100",
25540=>"111101111",
25541=>"011001011",
25542=>"001000100",
25543=>"101001101",
25544=>"000010000",
25545=>"111111000",
25546=>"110011011",
25547=>"101000000",
25548=>"100110111",
25549=>"000000100",
25550=>"010111101",
25551=>"100111011",
25552=>"010111010",
25553=>"111110110",
25554=>"111000101",
25555=>"111110111",
25556=>"001111111",
25557=>"010001011",
25558=>"111011010",
25559=>"100011010",
25560=>"100010111",
25561=>"000011111",
25562=>"000110100",
25563=>"000000000",
25564=>"000110010",
25565=>"010000000",
25566=>"010000001",
25567=>"000001001",
25568=>"011100011",
25569=>"010101101",
25570=>"000111111",
25571=>"000111011",
25572=>"001000000",
25573=>"010111010",
25574=>"110000101",
25575=>"000110110",
25576=>"000101111",
25577=>"000100000",
25578=>"011111100",
25579=>"011001100",
25580=>"111100000",
25581=>"110100111",
25582=>"010000011",
25583=>"000000100",
25584=>"101111111",
25585=>"110100111",
25586=>"000000010",
25587=>"000010010",
25588=>"000001011",
25589=>"011111000",
25590=>"000001000",
25591=>"001100000",
25592=>"000000000",
25593=>"000111010",
25594=>"110000000",
25595=>"000111111",
25596=>"000000000",
25597=>"000101101",
25598=>"000110110",
25599=>"000111011",
25600=>"000100101",
25601=>"101111111",
25602=>"111100100",
25603=>"000010011",
25604=>"111101101",
25605=>"000111100",
25606=>"011111101",
25607=>"100110100",
25608=>"000000001",
25609=>"111101100",
25610=>"101101100",
25611=>"101100100",
25612=>"000000111",
25613=>"000000111",
25614=>"111100100",
25615=>"111010000",
25616=>"000000100",
25617=>"111000000",
25618=>"011111000",
25619=>"111011000",
25620=>"111011111",
25621=>"111100100",
25622=>"101000111",
25623=>"001001000",
25624=>"000100000",
25625=>"000000000",
25626=>"000000111",
25627=>"111000100",
25628=>"000100000",
25629=>"011100101",
25630=>"000011111",
25631=>"101100100",
25632=>"000000000",
25633=>"111011011",
25634=>"011000100",
25635=>"000011011",
25636=>"000001110",
25637=>"000000100",
25638=>"100011011",
25639=>"010010000",
25640=>"001011011",
25641=>"001001100",
25642=>"111110101",
25643=>"000011010",
25644=>"100001011",
25645=>"000010011",
25646=>"000000111",
25647=>"111010110",
25648=>"001000101",
25649=>"111001001",
25650=>"000010011",
25651=>"001110100",
25652=>"010000001",
25653=>"101111111",
25654=>"000010110",
25655=>"111101101",
25656=>"011011101",
25657=>"111101100",
25658=>"111001100",
25659=>"111000100",
25660=>"011000000",
25661=>"010111111",
25662=>"111100000",
25663=>"000001111",
25664=>"000010000",
25665=>"000000101",
25666=>"111111110",
25667=>"000100111",
25668=>"111101111",
25669=>"111100100",
25670=>"000111111",
25671=>"000011010",
25672=>"000011111",
25673=>"110100111",
25674=>"110100101",
25675=>"111100101",
25676=>"111100000",
25677=>"010110011",
25678=>"111000010",
25679=>"111011100",
25680=>"111101000",
25681=>"000010010",
25682=>"111000111",
25683=>"000011001",
25684=>"111100100",
25685=>"011011011",
25686=>"011011011",
25687=>"100100101",
25688=>"100000100",
25689=>"000000000",
25690=>"111110000",
25691=>"001011111",
25692=>"001000111",
25693=>"111100101",
25694=>"100000011",
25695=>"001000111",
25696=>"000000011",
25697=>"111111100",
25698=>"011100100",
25699=>"111101101",
25700=>"111000011",
25701=>"111111100",
25702=>"000011011",
25703=>"100001000",
25704=>"010110111",
25705=>"011111000",
25706=>"100001000",
25707=>"000101011",
25708=>"000010111",
25709=>"111000001",
25710=>"000000101",
25711=>"111000000",
25712=>"110110111",
25713=>"001011111",
25714=>"110000000",
25715=>"000000000",
25716=>"100000011",
25717=>"010101100",
25718=>"011111100",
25719=>"000000011",
25720=>"000110011",
25721=>"110011111",
25722=>"101111111",
25723=>"110011101",
25724=>"110110010",
25725=>"000010010",
25726=>"110010010",
25727=>"111100100",
25728=>"000010101",
25729=>"010111100",
25730=>"000001001",
25731=>"000000111",
25732=>"010010100",
25733=>"001011011",
25734=>"000101001",
25735=>"001000000",
25736=>"010000101",
25737=>"111111000",
25738=>"001100100",
25739=>"001011010",
25740=>"100100011",
25741=>"100101100",
25742=>"111110100",
25743=>"111000000",
25744=>"011101011",
25745=>"000000111",
25746=>"011000000",
25747=>"001011111",
25748=>"001000000",
25749=>"101100100",
25750=>"111100100",
25751=>"000010011",
25752=>"001011001",
25753=>"100100111",
25754=>"000000011",
25755=>"000000000",
25756=>"111110111",
25757=>"101111111",
25758=>"001100110",
25759=>"111101000",
25760=>"000101001",
25761=>"000000100",
25762=>"000010101",
25763=>"000000101",
25764=>"111000110",
25765=>"110100010",
25766=>"000011111",
25767=>"000011011",
25768=>"110111000",
25769=>"010110000",
25770=>"000000100",
25771=>"111101100",
25772=>"000011011",
25773=>"100000000",
25774=>"101000000",
25775=>"100010010",
25776=>"110000000",
25777=>"111001011",
25778=>"111100110",
25779=>"000010010",
25780=>"010011011",
25781=>"010011111",
25782=>"000001011",
25783=>"000010010",
25784=>"110011000",
25785=>"010000001",
25786=>"000100100",
25787=>"000010011",
25788=>"111111111",
25789=>"010000011",
25790=>"000010001",
25791=>"000101101",
25792=>"001000100",
25793=>"000000000",
25794=>"100100111",
25795=>"111101000",
25796=>"111101101",
25797=>"000110010",
25798=>"100000000",
25799=>"000010010",
25800=>"010100000",
25801=>"111100100",
25802=>"000000000",
25803=>"111101101",
25804=>"111110100",
25805=>"011010011",
25806=>"011101100",
25807=>"111000011",
25808=>"111101000",
25809=>"001000111",
25810=>"000000010",
25811=>"010100111",
25812=>"111111110",
25813=>"001001010",
25814=>"011100100",
25815=>"000000100",
25816=>"001011011",
25817=>"111100000",
25818=>"001000100",
25819=>"011000000",
25820=>"000110101",
25821=>"100100011",
25822=>"111011111",
25823=>"000000010",
25824=>"111100100",
25825=>"101100100",
25826=>"111100000",
25827=>"000000001",
25828=>"000000000",
25829=>"110000111",
25830=>"111111000",
25831=>"100000000",
25832=>"011011011",
25833=>"000000000",
25834=>"101100001",
25835=>"000011111",
25836=>"000100111",
25837=>"001000011",
25838=>"000000000",
25839=>"000000000",
25840=>"001000000",
25841=>"110001000",
25842=>"000001101",
25843=>"111010111",
25844=>"000000110",
25845=>"111111100",
25846=>"011100000",
25847=>"000011011",
25848=>"011000001",
25849=>"010111111",
25850=>"000000001",
25851=>"000000111",
25852=>"111100100",
25853=>"000000000",
25854=>"000000001",
25855=>"111111000",
25856=>"011011101",
25857=>"000000100",
25858=>"101101101",
25859=>"010111000",
25860=>"011111010",
25861=>"100000101",
25862=>"010000011",
25863=>"000001000",
25864=>"000001110",
25865=>"000010001",
25866=>"000110111",
25867=>"001001100",
25868=>"000001111",
25869=>"000001111",
25870=>"111111001",
25871=>"111110010",
25872=>"000010111",
25873=>"010010111",
25874=>"100000110",
25875=>"011010100",
25876=>"000000000",
25877=>"110010000",
25878=>"000001100",
25879=>"000000000",
25880=>"000000010",
25881=>"111000111",
25882=>"000001011",
25883=>"010011000",
25884=>"000000000",
25885=>"110010000",
25886=>"101000111",
25887=>"000000111",
25888=>"111001101",
25889=>"000000101",
25890=>"100000010",
25891=>"110000010",
25892=>"001001011",
25893=>"100010100",
25894=>"000000011",
25895=>"000001111",
25896=>"010010000",
25897=>"101001000",
25898=>"101000110",
25899=>"001000010",
25900=>"111111111",
25901=>"111101100",
25902=>"011001000",
25903=>"011001001",
25904=>"000000000",
25905=>"001101111",
25906=>"010000100",
25907=>"110111111",
25908=>"101001111",
25909=>"111111100",
25910=>"000000100",
25911=>"000100000",
25912=>"000101001",
25913=>"111111000",
25914=>"000000110",
25915=>"011110001",
25916=>"001001001",
25917=>"111111011",
25918=>"001010000",
25919=>"011011001",
25920=>"000010111",
25921=>"010000000",
25922=>"100000111",
25923=>"000000110",
25924=>"000000000",
25925=>"000000110",
25926=>"100011010",
25927=>"010010111",
25928=>"111100101",
25929=>"010010000",
25930=>"010000000",
25931=>"000100100",
25932=>"000100000",
25933=>"111111110",
25934=>"101010000",
25935=>"101100001",
25936=>"101000111",
25937=>"111010010",
25938=>"001000100",
25939=>"001001001",
25940=>"001101001",
25941=>"100001101",
25942=>"111111100",
25943=>"101101110",
25944=>"101001101",
25945=>"110110110",
25946=>"000000101",
25947=>"000010111",
25948=>"000000000",
25949=>"001000001",
25950=>"000111111",
25951=>"000100001",
25952=>"000001111",
25953=>"110000101",
25954=>"101111111",
25955=>"000000100",
25956=>"111111110",
25957=>"011000001",
25958=>"111011001",
25959=>"000000010",
25960=>"110111000",
25961=>"111111100",
25962=>"000001111",
25963=>"000000110",
25964=>"111111111",
25965=>"110111010",
25966=>"000100000",
25967=>"111111101",
25968=>"101111101",
25969=>"001000100",
25970=>"000000001",
25971=>"001000000",
25972=>"010000000",
25973=>"101100100",
25974=>"000010110",
25975=>"100111111",
25976=>"000000011",
25977=>"110010000",
25978=>"001101111",
25979=>"111111100",
25980=>"111111001",
25981=>"100100000",
25982=>"010010111",
25983=>"001000000",
25984=>"010100101",
25985=>"101000010",
25986=>"010010010",
25987=>"110000111",
25988=>"111010010",
25989=>"010111111",
25990=>"001001001",
25991=>"001011000",
25992=>"111111101",
25993=>"110010101",
25994=>"010000000",
25995=>"010010011",
25996=>"000010001",
25997=>"001011001",
25998=>"110010110",
25999=>"000000001",
26000=>"111111101",
26001=>"111101000",
26002=>"011000001",
26003=>"001000100",
26004=>"011111111",
26005=>"000000001",
26006=>"011101111",
26007=>"000000000",
26008=>"010111111",
26009=>"110111111",
26010=>"010111000",
26011=>"000000010",
26012=>"000000000",
26013=>"011111111",
26014=>"000000000",
26015=>"111011000",
26016=>"101101101",
26017=>"000110111",
26018=>"111101101",
26019=>"000000001",
26020=>"000000101",
26021=>"110000000",
26022=>"101001111",
26023=>"011111001",
26024=>"111010110",
26025=>"001010011",
26026=>"100000000",
26027=>"000010111",
26028=>"110111111",
26029=>"001001000",
26030=>"000100101",
26031=>"000010010",
26032=>"011000011",
26033=>"011001001",
26034=>"010010010",
26035=>"001001001",
26036=>"011101001",
26037=>"010010011",
26038=>"011010000",
26039=>"010000001",
26040=>"100100110",
26041=>"110110100",
26042=>"000111110",
26043=>"000100010",
26044=>"111111000",
26045=>"110111010",
26046=>"101100101",
26047=>"010010000",
26048=>"001001101",
26049=>"010010000",
26050=>"010000101",
26051=>"111111110",
26052=>"010011000",
26053=>"110110111",
26054=>"111100000",
26055=>"110010110",
26056=>"101000011",
26057=>"000101111",
26058=>"110110011",
26059=>"111111111",
26060=>"000000000",
26061=>"111100100",
26062=>"000111111",
26063=>"000011010",
26064=>"011000000",
26065=>"110101111",
26066=>"000000100",
26067=>"010111110",
26068=>"001000111",
26069=>"100100100",
26070=>"111101000",
26071=>"110101000",
26072=>"111101101",
26073=>"100000111",
26074=>"101101001",
26075=>"000010010",
26076=>"000001001",
26077=>"000000010",
26078=>"101001101",
26079=>"000000100",
26080=>"000000111",
26081=>"000100000",
26082=>"000010110",
26083=>"101111110",
26084=>"001000101",
26085=>"010110111",
26086=>"010010010",
26087=>"010011010",
26088=>"000000000",
26089=>"000000000",
26090=>"000001111",
26091=>"101110111",
26092=>"101000101",
26093=>"000000000",
26094=>"001110000",
26095=>"001111010",
26096=>"111111000",
26097=>"011101111",
26098=>"100001100",
26099=>"001001101",
26100=>"110110110",
26101=>"000000101",
26102=>"000000000",
26103=>"000000001",
26104=>"000011011",
26105=>"010000100",
26106=>"111010010",
26107=>"000101000",
26108=>"110110110",
26109=>"000000001",
26110=>"111101110",
26111=>"011111111",
26112=>"111000000",
26113=>"000010111",
26114=>"000000110",
26115=>"111000101",
26116=>"110111111",
26117=>"110100101",
26118=>"000001101",
26119=>"000000100",
26120=>"011000000",
26121=>"000100000",
26122=>"000011001",
26123=>"000000000",
26124=>"110000000",
26125=>"101011011",
26126=>"100001000",
26127=>"111010110",
26128=>"000101011",
26129=>"010111111",
26130=>"111000000",
26131=>"000011111",
26132=>"010100110",
26133=>"111111101",
26134=>"000111011",
26135=>"101011110",
26136=>"111000000",
26137=>"111111111",
26138=>"111001000",
26139=>"000000111",
26140=>"000000111",
26141=>"101011000",
26142=>"100000001",
26143=>"111010010",
26144=>"000111111",
26145=>"111100000",
26146=>"000000010",
26147=>"011001111",
26148=>"011101101",
26149=>"000000000",
26150=>"111101101",
26151=>"101001110",
26152=>"111101001",
26153=>"000010111",
26154=>"000101101",
26155=>"000010000",
26156=>"000000111",
26157=>"001100000",
26158=>"001000100",
26159=>"101100110",
26160=>"011111110",
26161=>"111111001",
26162=>"000111111",
26163=>"111011001",
26164=>"000111110",
26165=>"000000001",
26166=>"000011010",
26167=>"111100100",
26168=>"000010101",
26169=>"001001001",
26170=>"111001000",
26171=>"000011111",
26172=>"001100101",
26173=>"101111010",
26174=>"010000000",
26175=>"010110011",
26176=>"001110010",
26177=>"011000000",
26178=>"110111000",
26179=>"111000100",
26180=>"111111101",
26181=>"100010111",
26182=>"000001101",
26183=>"101111111",
26184=>"110001001",
26185=>"011000111",
26186=>"111000100",
26187=>"111101011",
26188=>"000000010",
26189=>"110001100",
26190=>"011111111",
26191=>"000010110",
26192=>"010110110",
26193=>"100111110",
26194=>"001000101",
26195=>"010011000",
26196=>"000000100",
26197=>"000100101",
26198=>"001001100",
26199=>"000000101",
26200=>"000010101",
26201=>"000000011",
26202=>"010011001",
26203=>"111011001",
26204=>"100000000",
26205=>"111101001",
26206=>"011111111",
26207=>"111001001",
26208=>"000000000",
26209=>"111101000",
26210=>"111101000",
26211=>"100101011",
26212=>"111110100",
26213=>"000011111",
26214=>"110001011",
26215=>"011000000",
26216=>"111001000",
26217=>"000110001",
26218=>"000011111",
26219=>"111011000",
26220=>"111110000",
26221=>"111000000",
26222=>"111001100",
26223=>"000101111",
26224=>"010011101",
26225=>"000000000",
26226=>"000110011",
26227=>"110110100",
26228=>"110111111",
26229=>"111000101",
26230=>"111000000",
26231=>"000001010",
26232=>"000000111",
26233=>"000000111",
26234=>"001000000",
26235=>"111111101",
26236=>"100100111",
26237=>"111111100",
26238=>"000111010",
26239=>"111001000",
26240=>"010111000",
26241=>"000111000",
26242=>"000000000",
26243=>"101111010",
26244=>"011101000",
26245=>"101000000",
26246=>"100000000",
26247=>"111000000",
26248=>"110100101",
26249=>"101010110",
26250=>"011000101",
26251=>"101111111",
26252=>"001000100",
26253=>"100111101",
26254=>"010000000",
26255=>"000000110",
26256=>"011011011",
26257=>"111001000",
26258=>"101011011",
26259=>"111011011",
26260=>"101110010",
26261=>"011000000",
26262=>"011000000",
26263=>"000100000",
26264=>"010000111",
26265=>"000000111",
26266=>"111111111",
26267=>"000000010",
26268=>"111101101",
26269=>"011100001",
26270=>"110011000",
26271=>"000000010",
26272=>"001100000",
26273=>"000011010",
26274=>"111111001",
26275=>"000000110",
26276=>"100000000",
26277=>"110101001",
26278=>"000010001",
26279=>"010000000",
26280=>"000000010",
26281=>"000101100",
26282=>"111000000",
26283=>"000111110",
26284=>"001101010",
26285=>"000000000",
26286=>"001011011",
26287=>"011101000",
26288=>"000001100",
26289=>"111011001",
26290=>"011111100",
26291=>"010100110",
26292=>"010111111",
26293=>"000111111",
26294=>"000100111",
26295=>"001011111",
26296=>"000100100",
26297=>"011011000",
26298=>"000100000",
26299=>"110000000",
26300=>"110000000",
26301=>"111111000",
26302=>"010001001",
26303=>"000110111",
26304=>"101101000",
26305=>"001000000",
26306=>"111101111",
26307=>"011011000",
26308=>"111000000",
26309=>"101100111",
26310=>"000000100",
26311=>"011001011",
26312=>"111101100",
26313=>"000100110",
26314=>"101111110",
26315=>"010110100",
26316=>"000001111",
26317=>"001001110",
26318=>"000111010",
26319=>"111100000",
26320=>"000000110",
26321=>"011011001",
26322=>"011100100",
26323=>"111111010",
26324=>"111011111",
26325=>"100000100",
26326=>"111111101",
26327=>"111111001",
26328=>"000111111",
26329=>"111111000",
26330=>"100001101",
26331=>"111100000",
26332=>"000111111",
26333=>"100000000",
26334=>"000000111",
26335=>"111101000",
26336=>"111100101",
26337=>"111111001",
26338=>"000100100",
26339=>"011001101",
26340=>"000000101",
26341=>"000101111",
26342=>"000001111",
26343=>"100100100",
26344=>"111111101",
26345=>"100111111",
26346=>"100010110",
26347=>"100000011",
26348=>"101100100",
26349=>"000000100",
26350=>"110100000",
26351=>"000111010",
26352=>"000110011",
26353=>"001011101",
26354=>"000000101",
26355=>"010111111",
26356=>"000000100",
26357=>"101000000",
26358=>"111100000",
26359=>"000101111",
26360=>"111110111",
26361=>"111011101",
26362=>"001111001",
26363=>"000101101",
26364=>"011110000",
26365=>"100111010",
26366=>"000001111",
26367=>"010000100",
26368=>"110000000",
26369=>"110000000",
26370=>"110111010",
26371=>"111101111",
26372=>"001001001",
26373=>"100000000",
26374=>"110110010",
26375=>"000000001",
26376=>"000110111",
26377=>"111011001",
26378=>"111000110",
26379=>"101000001",
26380=>"000000000",
26381=>"000010000",
26382=>"110010001",
26383=>"011111111",
26384=>"000000110",
26385=>"110111110",
26386=>"000000000",
26387=>"000111111",
26388=>"010111110",
26389=>"111001000",
26390=>"100001001",
26391=>"010110011",
26392=>"000000000",
26393=>"111100010",
26394=>"100101110",
26395=>"100000100",
26396=>"000000000",
26397=>"100000000",
26398=>"010000000",
26399=>"101101101",
26400=>"100000111",
26401=>"000000000",
26402=>"000111001",
26403=>"111000101",
26404=>"111110000",
26405=>"000000000",
26406=>"011111010",
26407=>"111110111",
26408=>"111111001",
26409=>"111111001",
26410=>"110111110",
26411=>"001001001",
26412=>"111001001",
26413=>"100100000",
26414=>"000000000",
26415=>"000000000",
26416=>"000000001",
26417=>"100001001",
26418=>"000000000",
26419=>"111101111",
26420=>"010000000",
26421=>"111111110",
26422=>"111011011",
26423=>"000000000",
26424=>"000000000",
26425=>"101000000",
26426=>"010000100",
26427=>"111111001",
26428=>"001101100",
26429=>"000101000",
26430=>"101100001",
26431=>"011011011",
26432=>"111111111",
26433=>"000000010",
26434=>"100100000",
26435=>"000100100",
26436=>"110111111",
26437=>"101000101",
26438=>"000111111",
26439=>"011111111",
26440=>"000101001",
26441=>"110000010",
26442=>"111101001",
26443=>"110110010",
26444=>"101101001",
26445=>"011011000",
26446=>"110000000",
26447=>"101110000",
26448=>"001011001",
26449=>"010000000",
26450=>"001000111",
26451=>"001000101",
26452=>"000000000",
26453=>"100100100",
26454=>"100100100",
26455=>"000001111",
26456=>"001111111",
26457=>"011011001",
26458=>"100110110",
26459=>"111111111",
26460=>"001101101",
26461=>"110000000",
26462=>"010110110",
26463=>"000001011",
26464=>"001111111",
26465=>"001101000",
26466=>"000001101",
26467=>"100111101",
26468=>"101111100",
26469=>"001100000",
26470=>"011001100",
26471=>"110000001",
26472=>"110000111",
26473=>"000000011",
26474=>"001000101",
26475=>"001000000",
26476=>"011000110",
26477=>"111111110",
26478=>"000000000",
26479=>"111000000",
26480=>"100110111",
26481=>"001111000",
26482=>"111110110",
26483=>"000000000",
26484=>"000000001",
26485=>"011000000",
26486=>"111111100",
26487=>"110111010",
26488=>"111101101",
26489=>"111001001",
26490=>"111000111",
26491=>"000001111",
26492=>"001000110",
26493=>"000000001",
26494=>"010000000",
26495=>"000000101",
26496=>"010010000",
26497=>"000000000",
26498=>"111000010",
26499=>"111111100",
26500=>"101000000",
26501=>"111111011",
26502=>"000000010",
26503=>"001110011",
26504=>"011011011",
26505=>"110010000",
26506=>"011101000",
26507=>"011111111",
26508=>"111110111",
26509=>"000001111",
26510=>"000000111",
26511=>"100000111",
26512=>"001011011",
26513=>"000100111",
26514=>"100000000",
26515=>"001111111",
26516=>"000000111",
26517=>"001000110",
26518=>"100100000",
26519=>"100100000",
26520=>"000000000",
26521=>"001101000",
26522=>"110100111",
26523=>"000000100",
26524=>"100100000",
26525=>"111111011",
26526=>"010000001",
26527=>"111000011",
26528=>"111111111",
26529=>"111111000",
26530=>"011111111",
26531=>"111111111",
26532=>"011000000",
26533=>"110110110",
26534=>"001001001",
26535=>"111111010",
26536=>"111111111",
26537=>"001000111",
26538=>"000001111",
26539=>"111000000",
26540=>"001111101",
26541=>"101101100",
26542=>"101001000",
26543=>"000000101",
26544=>"000101101",
26545=>"111100110",
26546=>"000000000",
26547=>"001000000",
26548=>"111000000",
26549=>"111111011",
26550=>"111111110",
26551=>"111111101",
26552=>"100000000",
26553=>"000000100",
26554=>"101001000",
26555=>"000100111",
26556=>"010000000",
26557=>"101101111",
26558=>"001111110",
26559=>"010010010",
26560=>"000111111",
26561=>"011111010",
26562=>"010000010",
26563=>"101100100",
26564=>"010000000",
26565=>"100100000",
26566=>"000000000",
26567=>"100000000",
26568=>"111111101",
26569=>"111111111",
26570=>"111111011",
26571=>"111011111",
26572=>"111111101",
26573=>"100111011",
26574=>"000010010",
26575=>"000000000",
26576=>"101111000",
26577=>"011000000",
26578=>"100000000",
26579=>"100000100",
26580=>"001000101",
26581=>"001000000",
26582=>"001001101",
26583=>"010000011",
26584=>"000000000",
26585=>"111001111",
26586=>"110110110",
26587=>"000000011",
26588=>"101100001",
26589=>"101000111",
26590=>"111111110",
26591=>"000000000",
26592=>"111101000",
26593=>"000000000",
26594=>"000001101",
26595=>"110110100",
26596=>"000000100",
26597=>"010010111",
26598=>"111001111",
26599=>"111111000",
26600=>"011010000",
26601=>"101100001",
26602=>"100000101",
26603=>"000111111",
26604=>"000110000",
26605=>"001001001",
26606=>"000000000",
26607=>"000000111",
26608=>"000000000",
26609=>"001001011",
26610=>"000000111",
26611=>"011101001",
26612=>"011011001",
26613=>"110111111",
26614=>"000000000",
26615=>"000000111",
26616=>"010010111",
26617=>"010000000",
26618=>"111000000",
26619=>"000000000",
26620=>"011111100",
26621=>"100000111",
26622=>"111110110",
26623=>"000000000",
26624=>"111100110",
26625=>"001011000",
26626=>"111000000",
26627=>"111010101",
26628=>"110100110",
26629=>"111111111",
26630=>"111100100",
26631=>"000001000",
26632=>"000001001",
26633=>"111001011",
26634=>"000001000",
26635=>"100000000",
26636=>"110111111",
26637=>"001101000",
26638=>"110100000",
26639=>"111111010",
26640=>"110100010",
26641=>"000000001",
26642=>"100000000",
26643=>"011111000",
26644=>"000010000",
26645=>"000000001",
26646=>"111011000",
26647=>"011111000",
26648=>"101000101",
26649=>"101000000",
26650=>"011001111",
26651=>"111000110",
26652=>"001101101",
26653=>"101000000",
26654=>"111111111",
26655=>"110000000",
26656=>"111111110",
26657=>"111111101",
26658=>"001100000",
26659=>"010111010",
26660=>"100110010",
26661=>"011001101",
26662=>"000111111",
26663=>"000001000",
26664=>"000111010",
26665=>"111001111",
26666=>"111000000",
26667=>"101000001",
26668=>"110100010",
26669=>"001000000",
26670=>"011111111",
26671=>"111001001",
26672=>"011011000",
26673=>"010111111",
26674=>"101101010",
26675=>"111101001",
26676=>"101000000",
26677=>"111001111",
26678=>"111111111",
26679=>"000000000",
26680=>"010111001",
26681=>"000000100",
26682=>"000011000",
26683=>"111000010",
26684=>"001000000",
26685=>"100111111",
26686=>"111000010",
26687=>"000000100",
26688=>"101111000",
26689=>"000001110",
26690=>"111111000",
26691=>"001000111",
26692=>"000111011",
26693=>"000101111",
26694=>"011111010",
26695=>"100101000",
26696=>"101111010",
26697=>"100000000",
26698=>"011101111",
26699=>"000000000",
26700=>"000000111",
26701=>"011110111",
26702=>"001111111",
26703=>"000000111",
26704=>"000101001",
26705=>"111111111",
26706=>"000001010",
26707=>"000110000",
26708=>"000000000",
26709=>"111011010",
26710=>"011011001",
26711=>"000000000",
26712=>"011111000",
26713=>"001111010",
26714=>"011001000",
26715=>"010001011",
26716=>"111111011",
26717=>"000110000",
26718=>"101111101",
26719=>"100100111",
26720=>"100000101",
26721=>"010101011",
26722=>"000100101",
26723=>"010000000",
26724=>"111011001",
26725=>"010000001",
26726=>"111101101",
26727=>"111000111",
26728=>"111111100",
26729=>"011111111",
26730=>"000000111",
26731=>"110101111",
26732=>"111111111",
26733=>"011011001",
26734=>"101100101",
26735=>"000000111",
26736=>"000110111",
26737=>"000011111",
26738=>"011111111",
26739=>"111101000",
26740=>"000111111",
26741=>"111100111",
26742=>"011101000",
26743=>"111101111",
26744=>"001000000",
26745=>"010110100",
26746=>"000000000",
26747=>"010110011",
26748=>"000011000",
26749=>"100001000",
26750=>"001111110",
26751=>"000000000",
26752=>"010111101",
26753=>"001000000",
26754=>"001010111",
26755=>"010111111",
26756=>"000111011",
26757=>"100000001",
26758=>"000100001",
26759=>"000000110",
26760=>"000001111",
26761=>"000000000",
26762=>"110000000",
26763=>"101011010",
26764=>"000000000",
26765=>"000000000",
26766=>"000010010",
26767=>"001000000",
26768=>"111100011",
26769=>"110000000",
26770=>"000000110",
26771=>"101000110",
26772=>"100110000",
26773=>"000111101",
26774=>"111011000",
26775=>"000100000",
26776=>"101000000",
26777=>"101111000",
26778=>"010011011",
26779=>"111000000",
26780=>"010111000",
26781=>"111011001",
26782=>"111011000",
26783=>"000000000",
26784=>"011011110",
26785=>"100010000",
26786=>"000010011",
26787=>"111111001",
26788=>"101111100",
26789=>"000000000",
26790=>"001111000",
26791=>"001000100",
26792=>"000000111",
26793=>"111011000",
26794=>"111111000",
26795=>"010010000",
26796=>"101010000",
26797=>"101101111",
26798=>"000001001",
26799=>"000000001",
26800=>"000010000",
26801=>"000110110",
26802=>"101010011",
26803=>"011010010",
26804=>"111001000",
26805=>"001000000",
26806=>"110000101",
26807=>"001100101",
26808=>"110010000",
26809=>"011001001",
26810=>"010000100",
26811=>"111111111",
26812=>"000100001",
26813=>"010000000",
26814=>"100000000",
26815=>"000100111",
26816=>"000101100",
26817=>"101000000",
26818=>"010111000",
26819=>"010110110",
26820=>"000111011",
26821=>"110011111",
26822=>"010111001",
26823=>"101000111",
26824=>"010000010",
26825=>"000000000",
26826=>"011100110",
26827=>"011111010",
26828=>"100000000",
26829=>"000110000",
26830=>"110111000",
26831=>"111111001",
26832=>"000101101",
26833=>"010110011",
26834=>"011000000",
26835=>"111010110",
26836=>"101000000",
26837=>"000011000",
26838=>"110000000",
26839=>"100001111",
26840=>"000000000",
26841=>"000000000",
26842=>"110100011",
26843=>"111111000",
26844=>"111111000",
26845=>"110000000",
26846=>"100100000",
26847=>"101111111",
26848=>"000100000",
26849=>"011111111",
26850=>"110101111",
26851=>"011001001",
26852=>"000000000",
26853=>"111111111",
26854=>"000000000",
26855=>"000110010",
26856=>"000000100",
26857=>"000000000",
26858=>"000000000",
26859=>"100000011",
26860=>"011000000",
26861=>"001101011",
26862=>"000001000",
26863=>"000000000",
26864=>"000000110",
26865=>"010100110",
26866=>"101000111",
26867=>"001111000",
26868=>"011001011",
26869=>"111110000",
26870=>"000100111",
26871=>"111111000",
26872=>"000111010",
26873=>"000111101",
26874=>"000000000",
26875=>"000000000",
26876=>"111111011",
26877=>"111111111",
26878=>"000000000",
26879=>"000000000",
26880=>"100100110",
26881=>"111101000",
26882=>"100000111",
26883=>"111101010",
26884=>"000000000",
26885=>"000000000",
26886=>"011000100",
26887=>"111111000",
26888=>"000101110",
26889=>"011011000",
26890=>"110011001",
26891=>"111000000",
26892=>"010111000",
26893=>"000000000",
26894=>"110100010",
26895=>"111111111",
26896=>"010011000",
26897=>"010010010",
26898=>"010000000",
26899=>"000100000",
26900=>"010011000",
26901=>"000000100",
26902=>"000011111",
26903=>"110111111",
26904=>"111000000",
26905=>"011011111",
26906=>"101100000",
26907=>"111111111",
26908=>"000001111",
26909=>"000000000",
26910=>"001111110",
26911=>"100000011",
26912=>"111111100",
26913=>"000000000",
26914=>"100000000",
26915=>"000000011",
26916=>"000000001",
26917=>"000001111",
26918=>"000000010",
26919=>"000011100",
26920=>"000111111",
26921=>"000101000",
26922=>"010000100",
26923=>"110010000",
26924=>"111111001",
26925=>"011001111",
26926=>"100111010",
26927=>"000000000",
26928=>"111110001",
26929=>"001000011",
26930=>"101000111",
26931=>"111010000",
26932=>"000101000",
26933=>"011111010",
26934=>"100100000",
26935=>"000000001",
26936=>"111111010",
26937=>"110100111",
26938=>"110000000",
26939=>"111101111",
26940=>"001111101",
26941=>"111000111",
26942=>"100000000",
26943=>"111100100",
26944=>"111100010",
26945=>"000110011",
26946=>"000000111",
26947=>"111000111",
26948=>"000000000",
26949=>"100011001",
26950=>"111000111",
26951=>"001000000",
26952=>"010101110",
26953=>"011111111",
26954=>"100100100",
26955=>"111111110",
26956=>"000000000",
26957=>"100110100",
26958=>"001010100",
26959=>"101100100",
26960=>"000000000",
26961=>"010111111",
26962=>"111110101",
26963=>"101000100",
26964=>"000100111",
26965=>"001000100",
26966=>"101010000",
26967=>"111011011",
26968=>"000000010",
26969=>"000000100",
26970=>"001000000",
26971=>"111011111",
26972=>"000000110",
26973=>"110010000",
26974=>"000111100",
26975=>"111011011",
26976=>"111111111",
26977=>"000000100",
26978=>"000010010",
26979=>"100000000",
26980=>"100101111",
26981=>"011011010",
26982=>"000000000",
26983=>"101000111",
26984=>"101011111",
26985=>"000000000",
26986=>"010000000",
26987=>"010111111",
26988=>"111111101",
26989=>"011111011",
26990=>"000000000",
26991=>"111000000",
26992=>"000111001",
26993=>"110000000",
26994=>"000000000",
26995=>"010011011",
26996=>"010010000",
26997=>"111001011",
26998=>"100000001",
26999=>"010111000",
27000=>"100000001",
27001=>"000011111",
27002=>"101000101",
27003=>"000011011",
27004=>"001001101",
27005=>"101001000",
27006=>"111010010",
27007=>"111100111",
27008=>"101101100",
27009=>"111111011",
27010=>"000000011",
27011=>"000101000",
27012=>"011000000",
27013=>"100000000",
27014=>"100100101",
27015=>"110000000",
27016=>"010110100",
27017=>"000100111",
27018=>"011111001",
27019=>"000001111",
27020=>"000000011",
27021=>"111010000",
27022=>"000000111",
27023=>"000000100",
27024=>"110010010",
27025=>"000000000",
27026=>"001000000",
27027=>"111100000",
27028=>"000000100",
27029=>"110110000",
27030=>"111111000",
27031=>"110100110",
27032=>"010010001",
27033=>"010000011",
27034=>"010010000",
27035=>"111000000",
27036=>"111111111",
27037=>"111111000",
27038=>"100000000",
27039=>"111111111",
27040=>"000000010",
27041=>"111110111",
27042=>"111111111",
27043=>"110011000",
27044=>"101000000",
27045=>"100000000",
27046=>"010000110",
27047=>"111101100",
27048=>"000000000",
27049=>"001101000",
27050=>"000001000",
27051=>"000000000",
27052=>"011001010",
27053=>"100100100",
27054=>"110100101",
27055=>"011010000",
27056=>"111000001",
27057=>"101101010",
27058=>"000010111",
27059=>"100000000",
27060=>"111011000",
27061=>"001000000",
27062=>"000000000",
27063=>"000001001",
27064=>"010000011",
27065=>"010011101",
27066=>"000010011",
27067=>"111111111",
27068=>"001111111",
27069=>"011111111",
27070=>"111111001",
27071=>"111010000",
27072=>"011000100",
27073=>"000000000",
27074=>"111111111",
27075=>"000000000",
27076=>"000111111",
27077=>"010111100",
27078=>"011111011",
27079=>"111000000",
27080=>"011111010",
27081=>"100000000",
27082=>"000000100",
27083=>"000000000",
27084=>"111100101",
27085=>"110110001",
27086=>"100100100",
27087=>"111111111",
27088=>"111111111",
27089=>"100011011",
27090=>"100100101",
27091=>"101111011",
27092=>"101000100",
27093=>"111111111",
27094=>"100000000",
27095=>"011010000",
27096=>"000101101",
27097=>"000110101",
27098=>"000100101",
27099=>"011010000",
27100=>"100110101",
27101=>"011111001",
27102=>"101001000",
27103=>"111111011",
27104=>"000000000",
27105=>"101011011",
27106=>"111111111",
27107=>"111011000",
27108=>"000001100",
27109=>"011011010",
27110=>"000000000",
27111=>"000100100",
27112=>"000000011",
27113=>"111111000",
27114=>"110110110",
27115=>"011011000",
27116=>"001111011",
27117=>"000000100",
27118=>"100010111",
27119=>"000000000",
27120=>"101111111",
27121=>"000000100",
27122=>"000100111",
27123=>"100100000",
27124=>"001001111",
27125=>"000000000",
27126=>"011011010",
27127=>"100010111",
27128=>"000010000",
27129=>"111111101",
27130=>"000000000",
27131=>"000110111",
27132=>"000000111",
27133=>"000011111",
27134=>"001000001",
27135=>"111111000",
27136=>"000000100",
27137=>"000000011",
27138=>"111000000",
27139=>"110000111",
27140=>"000001001",
27141=>"010011001",
27142=>"001000001",
27143=>"000001110",
27144=>"000011001",
27145=>"100000000",
27146=>"000100011",
27147=>"101101111",
27148=>"000100101",
27149=>"100110110",
27150=>"000001000",
27151=>"011011001",
27152=>"100101000",
27153=>"110111001",
27154=>"111101000",
27155=>"011111111",
27156=>"011011101",
27157=>"111111011",
27158=>"111111001",
27159=>"111111101",
27160=>"001010000",
27161=>"101000000",
27162=>"100011011",
27163=>"000000000",
27164=>"011011010",
27165=>"011010010",
27166=>"110001000",
27167=>"000000111",
27168=>"000010110",
27169=>"111010011",
27170=>"001000111",
27171=>"001111111",
27172=>"000000000",
27173=>"011011111",
27174=>"100010010",
27175=>"001000001",
27176=>"001000010",
27177=>"000000111",
27178=>"101111101",
27179=>"000001111",
27180=>"000000111",
27181=>"011111111",
27182=>"010010111",
27183=>"000000001",
27184=>"111111110",
27185=>"101101000",
27186=>"000000101",
27187=>"111001000",
27188=>"000000010",
27189=>"000111110",
27190=>"011011110",
27191=>"110111100",
27192=>"111101000",
27193=>"000001000",
27194=>"000000101",
27195=>"111111011",
27196=>"000111011",
27197=>"111010110",
27198=>"000001000",
27199=>"111011011",
27200=>"111001000",
27201=>"010111010",
27202=>"111000100",
27203=>"111011100",
27204=>"111100111",
27205=>"000000111",
27206=>"000000000",
27207=>"001000000",
27208=>"000111110",
27209=>"000001111",
27210=>"000000000",
27211=>"100111010",
27212=>"011000000",
27213=>"000111011",
27214=>"001001000",
27215=>"110111111",
27216=>"011010111",
27217=>"111010000",
27218=>"011111111",
27219=>"011011101",
27220=>"001000110",
27221=>"111111000",
27222=>"000010010",
27223=>"111000000",
27224=>"000000000",
27225=>"000000011",
27226=>"000000111",
27227=>"110000110",
27228=>"100111000",
27229=>"000001001",
27230=>"111010111",
27231=>"111101001",
27232=>"110000000",
27233=>"000010011",
27234=>"110000000",
27235=>"000001110",
27236=>"000100111",
27237=>"101000111",
27238=>"000111111",
27239=>"001110111",
27240=>"001001111",
27241=>"000000000",
27242=>"110100101",
27243=>"010000000",
27244=>"010011010",
27245=>"000000111",
27246=>"000100101",
27247=>"000000001",
27248=>"011101111",
27249=>"000000000",
27250=>"110110011",
27251=>"101110010",
27252=>"111001010",
27253=>"011000000",
27254=>"000000000",
27255=>"111110010",
27256=>"000000100",
27257=>"000101101",
27258=>"000001000",
27259=>"101100111",
27260=>"011001100",
27261=>"010100100",
27262=>"111110110",
27263=>"111001100",
27264=>"111010000",
27265=>"111111101",
27266=>"010010000",
27267=>"000011110",
27268=>"011111101",
27269=>"111111111",
27270=>"110110110",
27271=>"000100000",
27272=>"100111011",
27273=>"101110110",
27274=>"000011110",
27275=>"001000110",
27276=>"111000000",
27277=>"011110110",
27278=>"111111000",
27279=>"111101000",
27280=>"001011101",
27281=>"000100000",
27282=>"001000000",
27283=>"000001000",
27284=>"000111000",
27285=>"111100000",
27286=>"111010111",
27287=>"000011111",
27288=>"000000111",
27289=>"100000100",
27290=>"111101001",
27291=>"111100100",
27292=>"111000010",
27293=>"111110100",
27294=>"111101011",
27295=>"000001000",
27296=>"000000001",
27297=>"011000110",
27298=>"000111101",
27299=>"100100101",
27300=>"100001100",
27301=>"011010111",
27302=>"111111111",
27303=>"001010001",
27304=>"111010111",
27305=>"111101111",
27306=>"111111101",
27307=>"111101110",
27308=>"000000110",
27309=>"111001000",
27310=>"000000011",
27311=>"100100101",
27312=>"011111100",
27313=>"000001001",
27314=>"000000000",
27315=>"001101100",
27316=>"000111111",
27317=>"000110111",
27318=>"000011000",
27319=>"000001100",
27320=>"000111111",
27321=>"000001001",
27322=>"011110110",
27323=>"001101000",
27324=>"000001010",
27325=>"111111100",
27326=>"100000001",
27327=>"000111111",
27328=>"000000000",
27329=>"000111110",
27330=>"011111111",
27331=>"000000110",
27332=>"001000000",
27333=>"001010101",
27334=>"000000000",
27335=>"111000100",
27336=>"000001101",
27337=>"110010000",
27338=>"011010000",
27339=>"111100010",
27340=>"000000000",
27341=>"100100101",
27342=>"000000101",
27343=>"111000000",
27344=>"000010111",
27345=>"110110111",
27346=>"000001011",
27347=>"000000000",
27348=>"111101000",
27349=>"000100111",
27350=>"110110111",
27351=>"001101111",
27352=>"000000111",
27353=>"000111111",
27354=>"011000000",
27355=>"111101000",
27356=>"111110000",
27357=>"111001111",
27358=>"101111001",
27359=>"000100000",
27360=>"111111000",
27361=>"110000111",
27362=>"001000100",
27363=>"101111111",
27364=>"000100111",
27365=>"000110111",
27366=>"010011100",
27367=>"000000111",
27368=>"001010110",
27369=>"000010111",
27370=>"001001111",
27371=>"001101101",
27372=>"000000000",
27373=>"000010000",
27374=>"111000000",
27375=>"000101101",
27376=>"011011110",
27377=>"111011111",
27378=>"100000000",
27379=>"010011101",
27380=>"000011001",
27381=>"100000111",
27382=>"001000000",
27383=>"101010110",
27384=>"100000000",
27385=>"001000011",
27386=>"010110111",
27387=>"000010110",
27388=>"110110100",
27389=>"111111111",
27390=>"100111001",
27391=>"001100000",
27392=>"011000101",
27393=>"100000000",
27394=>"111111111",
27395=>"110010000",
27396=>"010111111",
27397=>"010100111",
27398=>"101100100",
27399=>"000000000",
27400=>"110111100",
27401=>"000100000",
27402=>"000001000",
27403=>"000000000",
27404=>"111100000",
27405=>"000000000",
27406=>"100100100",
27407=>"010111111",
27408=>"111111000",
27409=>"101111001",
27410=>"111111110",
27411=>"101011111",
27412=>"000000100",
27413=>"110110010",
27414=>"000011111",
27415=>"111000010",
27416=>"100000000",
27417=>"000000000",
27418=>"100000000",
27419=>"000011111",
27420=>"001111111",
27421=>"011101011",
27422=>"000000100",
27423=>"101101101",
27424=>"010111111",
27425=>"000000000",
27426=>"111101000",
27427=>"110101010",
27428=>"010110000",
27429=>"000011011",
27430=>"111000000",
27431=>"000111010",
27432=>"000000000",
27433=>"111111110",
27434=>"111011111",
27435=>"000111100",
27436=>"000100100",
27437=>"111001000",
27438=>"000111111",
27439=>"001011010",
27440=>"111001000",
27441=>"100100101",
27442=>"000000000",
27443=>"000000000",
27444=>"000111110",
27445=>"111011011",
27446=>"100100001",
27447=>"000011011",
27448=>"000011000",
27449=>"000000000",
27450=>"000100000",
27451=>"111111111",
27452=>"110011011",
27453=>"111111011",
27454=>"000100111",
27455=>"111010011",
27456=>"111111000",
27457=>"011000111",
27458=>"000001000",
27459=>"010011011",
27460=>"010011010",
27461=>"100111111",
27462=>"000000110",
27463=>"000000101",
27464=>"000001000",
27465=>"000000101",
27466=>"110100001",
27467=>"101000000",
27468=>"111111111",
27469=>"011011011",
27470=>"011011101",
27471=>"101001111",
27472=>"101101111",
27473=>"001111010",
27474=>"000100101",
27475=>"010110110",
27476=>"100000001",
27477=>"000110110",
27478=>"001001001",
27479=>"111000001",
27480=>"110000000",
27481=>"110111100",
27482=>"001011011",
27483=>"110111011",
27484=>"000000100",
27485=>"100110000",
27486=>"000111110",
27487=>"110110111",
27488=>"000000000",
27489=>"111101101",
27490=>"101000000",
27491=>"000110110",
27492=>"011111111",
27493=>"000111110",
27494=>"000000000",
27495=>"000010010",
27496=>"101010100",
27497=>"111010000",
27498=>"000000010",
27499=>"000001111",
27500=>"111010010",
27501=>"000000111",
27502=>"000110111",
27503=>"010000010",
27504=>"000111100",
27505=>"111001000",
27506=>"001010110",
27507=>"001000000",
27508=>"101011000",
27509=>"000000011",
27510=>"101001000",
27511=>"011011111",
27512=>"000010100",
27513=>"111011111",
27514=>"111101001",
27515=>"000001100",
27516=>"011101111",
27517=>"000000010",
27518=>"111111111",
27519=>"101000001",
27520=>"111101111",
27521=>"010100000",
27522=>"111111010",
27523=>"011111111",
27524=>"000000000",
27525=>"000111110",
27526=>"000111111",
27527=>"110100000",
27528=>"000111010",
27529=>"010111001",
27530=>"001011010",
27531=>"000101111",
27532=>"000000000",
27533=>"011111000",
27534=>"000111110",
27535=>"010001011",
27536=>"011011111",
27537=>"000000111",
27538=>"000010101",
27539=>"111101100",
27540=>"111111111",
27541=>"111111011",
27542=>"000111100",
27543=>"111100000",
27544=>"011101001",
27545=>"101000100",
27546=>"000000011",
27547=>"111111010",
27548=>"000000000",
27549=>"010011010",
27550=>"100101111",
27551=>"101000000",
27552=>"100101001",
27553=>"010110111",
27554=>"000100101",
27555=>"111101101",
27556=>"111000001",
27557=>"010111011",
27558=>"010001011",
27559=>"000000000",
27560=>"000000011",
27561=>"110101000",
27562=>"111001001",
27563=>"000000101",
27564=>"111111000",
27565=>"000011001",
27566=>"110111111",
27567=>"111111111",
27568=>"100100000",
27569=>"111001000",
27570=>"011011001",
27571=>"111000000",
27572=>"110010011",
27573=>"100101010",
27574=>"011101110",
27575=>"000000011",
27576=>"110111100",
27577=>"111111100",
27578=>"000001110",
27579=>"100010111",
27580=>"000100000",
27581=>"110111111",
27582=>"111110100",
27583=>"111100000",
27584=>"111111111",
27585=>"000011110",
27586=>"011000000",
27587=>"110000011",
27588=>"000000001",
27589=>"100011010",
27590=>"010010001",
27591=>"011111111",
27592=>"000010100",
27593=>"110000111",
27594=>"111111111",
27595=>"000101001",
27596=>"000111111",
27597=>"110111111",
27598=>"100111111",
27599=>"110011000",
27600=>"111111111",
27601=>"011110110",
27602=>"111100101",
27603=>"101110000",
27604=>"001101101",
27605=>"000000000",
27606=>"000000000",
27607=>"111100000",
27608=>"000000000",
27609=>"111000000",
27610=>"010110100",
27611=>"001000000",
27612=>"111110111",
27613=>"111101000",
27614=>"111101011",
27615=>"111111010",
27616=>"101000001",
27617=>"101101111",
27618=>"000001101",
27619=>"111111100",
27620=>"000000100",
27621=>"111001001",
27622=>"110111011",
27623=>"110110111",
27624=>"100101001",
27625=>"000000000",
27626=>"000100011",
27627=>"111101000",
27628=>"111100100",
27629=>"000011001",
27630=>"111010000",
27631=>"101000000",
27632=>"111011000",
27633=>"000101111",
27634=>"000000100",
27635=>"010111001",
27636=>"010000011",
27637=>"000000000",
27638=>"000111110",
27639=>"110100001",
27640=>"111111111",
27641=>"111011001",
27642=>"000100111",
27643=>"110110010",
27644=>"001000011",
27645=>"011000111",
27646=>"000110111",
27647=>"010111011",
27648=>"111000001",
27649=>"000010111",
27650=>"100100110",
27651=>"010000110",
27652=>"100001001",
27653=>"011110000",
27654=>"111101000",
27655=>"001000001",
27656=>"000111111",
27657=>"000101011",
27658=>"001011001",
27659=>"111111101",
27660=>"101001001",
27661=>"001111010",
27662=>"000101001",
27663=>"001011000",
27664=>"111110111",
27665=>"000111000",
27666=>"010110011",
27667=>"110101111",
27668=>"111100011",
27669=>"010100100",
27670=>"100100100",
27671=>"100011011",
27672=>"111110011",
27673=>"001011000",
27674=>"001100010",
27675=>"000101100",
27676=>"111111100",
27677=>"111111000",
27678=>"111100100",
27679=>"110001001",
27680=>"011000001",
27681=>"111111111",
27682=>"111110011",
27683=>"111101100",
27684=>"011001010",
27685=>"101011001",
27686=>"111110111",
27687=>"000011001",
27688=>"000110011",
27689=>"100110111",
27690=>"111110000",
27691=>"100010000",
27692=>"100111100",
27693=>"001010111",
27694=>"000110000",
27695=>"111100000",
27696=>"011010001",
27697=>"000100100",
27698=>"001000110",
27699=>"111100101",
27700=>"111011011",
27701=>"000000000",
27702=>"000000001",
27703=>"000001000",
27704=>"110110111",
27705=>"101000011",
27706=>"000001000",
27707=>"000001100",
27708=>"100100100",
27709=>"111111111",
27710=>"000000100",
27711=>"101111110",
27712=>"000110100",
27713=>"100001011",
27714=>"010110001",
27715=>"011001110",
27716=>"001111100",
27717=>"000000010",
27718=>"000001001",
27719=>"111110111",
27720=>"111110011",
27721=>"001001011",
27722=>"011000011",
27723=>"000011011",
27724=>"000100010",
27725=>"100100110",
27726=>"110111111",
27727=>"111111111",
27728=>"100100100",
27729=>"011111100",
27730=>"001001001",
27731=>"001001000",
27732=>"010111110",
27733=>"001010101",
27734=>"001011100",
27735=>"011100011",
27736=>"111111111",
27737=>"101000000",
27738=>"011101001",
27739=>"000001101",
27740=>"000011011",
27741=>"010000011",
27742=>"110111100",
27743=>"111010000",
27744=>"000110111",
27745=>"000100100",
27746=>"110110010",
27747=>"101011000",
27748=>"000000011",
27749=>"100001001",
27750=>"000001000",
27751=>"010100000",
27752=>"011111111",
27753=>"001000000",
27754=>"000010110",
27755=>"000011001",
27756=>"010100100",
27757=>"101100000",
27758=>"110000100",
27759=>"100101010",
27760=>"000110100",
27761=>"000000001",
27762=>"110101111",
27763=>"111101011",
27764=>"001001000",
27765=>"110000000",
27766=>"100011101",
27767=>"111100110",
27768=>"110100010",
27769=>"011111001",
27770=>"100000101",
27771=>"101101001",
27772=>"110110110",
27773=>"011011011",
27774=>"001000001",
27775=>"100010011",
27776=>"010001000",
27777=>"111110100",
27778=>"011011011",
27779=>"000101111",
27780=>"001101111",
27781=>"111011011",
27782=>"110001001",
27783=>"000000001",
27784=>"101101111",
27785=>"100100000",
27786=>"000001011",
27787=>"000001010",
27788=>"100110110",
27789=>"100000001",
27790=>"111011011",
27791=>"100000010",
27792=>"101110101",
27793=>"000001111",
27794=>"000001011",
27795=>"111101111",
27796=>"001011010",
27797=>"010100000",
27798=>"000000000",
27799=>"011010101",
27800=>"001000001",
27801=>"110100000",
27802=>"111110111",
27803=>"111110011",
27804=>"000000110",
27805=>"111110111",
27806=>"000000000",
27807=>"100101001",
27808=>"010001101",
27809=>"110000100",
27810=>"011110011",
27811=>"101110111",
27812=>"111100001",
27813=>"000011111",
27814=>"011000000",
27815=>"000001001",
27816=>"000100011",
27817=>"100111100",
27818=>"001111100",
27819=>"001110110",
27820=>"110100111",
27821=>"010010011",
27822=>"001110000",
27823=>"011000001",
27824=>"001011000",
27825=>"000000010",
27826=>"011011000",
27827=>"111100110",
27828=>"000001001",
27829=>"001010000",
27830=>"000000001",
27831=>"000000010",
27832=>"100000001",
27833=>"011101011",
27834=>"001101000",
27835=>"011000011",
27836=>"000011000",
27837=>"001111011",
27838=>"000000001",
27839=>"000001101",
27840=>"111100001",
27841=>"000100111",
27842=>"111111111",
27843=>"101101111",
27844=>"000001001",
27845=>"010010111",
27846=>"000001001",
27847=>"101110100",
27848=>"001001000",
27849=>"111000011",
27850=>"101110111",
27851=>"000011001",
27852=>"111101000",
27853=>"000110110",
27854=>"000001001",
27855=>"000000011",
27856=>"111101100",
27857=>"011000000",
27858=>"100001111",
27859=>"001001000",
27860=>"111010000",
27861=>"010111110",
27862=>"101010110",
27863=>"001001000",
27864=>"001010011",
27865=>"001001001",
27866=>"100111110",
27867=>"001000000",
27868=>"011110100",
27869=>"000111110",
27870=>"100010000",
27871=>"111101001",
27872=>"110110100",
27873=>"010100110",
27874=>"011011000",
27875=>"000110110",
27876=>"110100101",
27877=>"000111000",
27878=>"101111111",
27879=>"000101100",
27880=>"001000000",
27881=>"001011001",
27882=>"110001011",
27883=>"111110110",
27884=>"001001011",
27885=>"001011000",
27886=>"001001001",
27887=>"111010000",
27888=>"101000011",
27889=>"111100101",
27890=>"011111000",
27891=>"110111001",
27892=>"001110110",
27893=>"001101100",
27894=>"011010011",
27895=>"111000000",
27896=>"110100111",
27897=>"111011000",
27898=>"111110000",
27899=>"000011000",
27900=>"010011000",
27901=>"000001000",
27902=>"001001011",
27903=>"111110100",
27904=>"000000000",
27905=>"100100001",
27906=>"101000000",
27907=>"000000000",
27908=>"010111101",
27909=>"001011110",
27910=>"111111000",
27911=>"000000111",
27912=>"010010100",
27913=>"000000000",
27914=>"110001000",
27915=>"111101101",
27916=>"110111101",
27917=>"111111001",
27918=>"000100111",
27919=>"100001010",
27920=>"111111111",
27921=>"001111000",
27922=>"000111000",
27923=>"111111111",
27924=>"010110111",
27925=>"000001011",
27926=>"111110100",
27927=>"101110111",
27928=>"000000000",
27929=>"111111101",
27930=>"000000000",
27931=>"000000010",
27932=>"111111101",
27933=>"101101000",
27934=>"111000000",
27935=>"000101101",
27936=>"111111111",
27937=>"111111010",
27938=>"000000000",
27939=>"000000110",
27940=>"111111011",
27941=>"010100110",
27942=>"111101000",
27943=>"001000011",
27944=>"010111111",
27945=>"101110111",
27946=>"000110110",
27947=>"110111111",
27948=>"111111111",
27949=>"000110011",
27950=>"111111111",
27951=>"000000000",
27952=>"111001000",
27953=>"110110110",
27954=>"001000000",
27955=>"010010111",
27956=>"100000000",
27957=>"110101010",
27958=>"110111011",
27959=>"000000000",
27960=>"011001100",
27961=>"000000000",
27962=>"000000000",
27963=>"000000000",
27964=>"110000110",
27965=>"010111000",
27966=>"110000000",
27967=>"100100111",
27968=>"100110101",
27969=>"111101000",
27970=>"111110100",
27971=>"111100000",
27972=>"010111000",
27973=>"001101111",
27974=>"111111011",
27975=>"000111111",
27976=>"000000011",
27977=>"000010111",
27978=>"111010000",
27979=>"110110111",
27980=>"101000000",
27981=>"000110110",
27982=>"010110111",
27983=>"111110011",
27984=>"111000001",
27985=>"111110000",
27986=>"000010011",
27987=>"001000000",
27988=>"111000000",
27989=>"100100010",
27990=>"100110000",
27991=>"111101000",
27992=>"000000001",
27993=>"110110111",
27994=>"000100000",
27995=>"111111011",
27996=>"111101101",
27997=>"000000000",
27998=>"000000000",
27999=>"111111001",
28000=>"111111111",
28001=>"000111111",
28002=>"110111111",
28003=>"100000000",
28004=>"000000000",
28005=>"111010000",
28006=>"110111000",
28007=>"000000101",
28008=>"111111111",
28009=>"000000111",
28010=>"010110110",
28011=>"110010010",
28012=>"110111011",
28013=>"000000000",
28014=>"111111000",
28015=>"111010000",
28016=>"010110110",
28017=>"000000101",
28018=>"111101110",
28019=>"111111111",
28020=>"011000000",
28021=>"000000001",
28022=>"000111111",
28023=>"000101001",
28024=>"100111111",
28025=>"110110000",
28026=>"000110111",
28027=>"010010010",
28028=>"011000100",
28029=>"000000000",
28030=>"000010110",
28031=>"010000000",
28032=>"110011000",
28033=>"111100000",
28034=>"000111101",
28035=>"001010000",
28036=>"010000000",
28037=>"110111011",
28038=>"111100001",
28039=>"010011101",
28040=>"001011111",
28041=>"000001000",
28042=>"000000010",
28043=>"101111111",
28044=>"000000000",
28045=>"011001001",
28046=>"000000000",
28047=>"000000101",
28048=>"000010000",
28049=>"000000111",
28050=>"100000010",
28051=>"111110111",
28052=>"000110111",
28053=>"000000100",
28054=>"010000000",
28055=>"010110001",
28056=>"000000100",
28057=>"111111111",
28058=>"111111110",
28059=>"010110000",
28060=>"000010000",
28061=>"011111111",
28062=>"000110110",
28063=>"000000000",
28064=>"001011100",
28065=>"110110000",
28066=>"111100110",
28067=>"000000000",
28068=>"010011010",
28069=>"110110100",
28070=>"001000000",
28071=>"000111000",
28072=>"000000110",
28073=>"000001000",
28074=>"000110100",
28075=>"000110110",
28076=>"010111001",
28077=>"101000111",
28078=>"110011011",
28079=>"011111111",
28080=>"000010000",
28081=>"011100100",
28082=>"000000011",
28083=>"011111100",
28084=>"100100001",
28085=>"011111010",
28086=>"110110000",
28087=>"000101111",
28088=>"001000011",
28089=>"001110100",
28090=>"000000000",
28091=>"011111100",
28092=>"010011111",
28093=>"011111110",
28094=>"001011011",
28095=>"111000000",
28096=>"101000000",
28097=>"001000111",
28098=>"111111101",
28099=>"110001000",
28100=>"101000000",
28101=>"010100100",
28102=>"000111111",
28103=>"000001011",
28104=>"111111101",
28105=>"000111011",
28106=>"101111111",
28107=>"111111100",
28108=>"100010110",
28109=>"110001000",
28110=>"110110111",
28111=>"100111110",
28112=>"101111111",
28113=>"111110011",
28114=>"011111101",
28115=>"101000001",
28116=>"001000111",
28117=>"100001000",
28118=>"000000000",
28119=>"110000000",
28120=>"111000111",
28121=>"110000111",
28122=>"110111001",
28123=>"000010000",
28124=>"110011001",
28125=>"000111111",
28126=>"110010000",
28127=>"000010111",
28128=>"000010010",
28129=>"101000100",
28130=>"001000000",
28131=>"100110110",
28132=>"100000000",
28133=>"000001001",
28134=>"000110111",
28135=>"011001001",
28136=>"111111111",
28137=>"111101111",
28138=>"010010000",
28139=>"000010110",
28140=>"101111111",
28141=>"110100000",
28142=>"000110000",
28143=>"000011101",
28144=>"000101000",
28145=>"000011000",
28146=>"101101000",
28147=>"010011010",
28148=>"000100010",
28149=>"000010000",
28150=>"000101011",
28151=>"111000101",
28152=>"010000000",
28153=>"001111101",
28154=>"010010101",
28155=>"010000000",
28156=>"010010100",
28157=>"000000000",
28158=>"000110100",
28159=>"010010000",
28160=>"011001101",
28161=>"000000011",
28162=>"101101001",
28163=>"100000100",
28164=>"000000101",
28165=>"000000100",
28166=>"111111111",
28167=>"001010000",
28168=>"111000000",
28169=>"111000100",
28170=>"000110110",
28171=>"000000000",
28172=>"001000101",
28173=>"110000000",
28174=>"011000000",
28175=>"111111111",
28176=>"000011111",
28177=>"000000000",
28178=>"111000000",
28179=>"000100000",
28180=>"000000110",
28181=>"000000000",
28182=>"000111011",
28183=>"100000010",
28184=>"100000100",
28185=>"011111111",
28186=>"001000110",
28187=>"000011011",
28188=>"111111010",
28189=>"110010000",
28190=>"001111100",
28191=>"000000000",
28192=>"011010000",
28193=>"111101100",
28194=>"101111111",
28195=>"101000000",
28196=>"110110000",
28197=>"110101100",
28198=>"000000000",
28199=>"000000110",
28200=>"000011000",
28201=>"000000000",
28202=>"110100010",
28203=>"111111110",
28204=>"011010000",
28205=>"011001111",
28206=>"010000111",
28207=>"101100101",
28208=>"001000110",
28209=>"000111111",
28210=>"101000111",
28211=>"011111010",
28212=>"010111111",
28213=>"000000000",
28214=>"001011110",
28215=>"111111101",
28216=>"011000111",
28217=>"100000000",
28218=>"111111010",
28219=>"111111111",
28220=>"000111000",
28221=>"111111100",
28222=>"000000000",
28223=>"100011001",
28224=>"111111111",
28225=>"011010010",
28226=>"111111101",
28227=>"000000011",
28228=>"000000000",
28229=>"000000000",
28230=>"000100010",
28231=>"010000000",
28232=>"001001100",
28233=>"010111110",
28234=>"101000111",
28235=>"111111111",
28236=>"111100000",
28237=>"000000001",
28238=>"000001111",
28239=>"000000011",
28240=>"111111010",
28241=>"111111010",
28242=>"100000111",
28243=>"011001001",
28244=>"000010110",
28245=>"111111111",
28246=>"011111010",
28247=>"100101111",
28248=>"000000010",
28249=>"010100000",
28250=>"001011111",
28251=>"000100011",
28252=>"111111000",
28253=>"001011011",
28254=>"111111111",
28255=>"011011110",
28256=>"010000000",
28257=>"101011010",
28258=>"101000101",
28259=>"110111110",
28260=>"000001011",
28261=>"010111011",
28262=>"010010010",
28263=>"011000000",
28264=>"001111111",
28265=>"000001011",
28266=>"111111010",
28267=>"010000000",
28268=>"000000000",
28269=>"000100001",
28270=>"000000101",
28271=>"001001101",
28272=>"000100100",
28273=>"000000000",
28274=>"010110010",
28275=>"000101111",
28276=>"110001000",
28277=>"111000100",
28278=>"100101000",
28279=>"000001000",
28280=>"000011000",
28281=>"111111000",
28282=>"100111111",
28283=>"101000101",
28284=>"111111111",
28285=>"100100101",
28286=>"110111111",
28287=>"010000000",
28288=>"111001100",
28289=>"011111000",
28290=>"000000010",
28291=>"111111111",
28292=>"000101000",
28293=>"101001111",
28294=>"000110001",
28295=>"011011011",
28296=>"101001010",
28297=>"000000100",
28298=>"001011111",
28299=>"000000000",
28300=>"000100100",
28301=>"101000100",
28302=>"100000000",
28303=>"101001101",
28304=>"001000011",
28305=>"000010010",
28306=>"000000111",
28307=>"111010000",
28308=>"001111011",
28309=>"101100000",
28310=>"111111100",
28311=>"000000000",
28312=>"001000000",
28313=>"101100111",
28314=>"101101000",
28315=>"111011101",
28316=>"101000000",
28317=>"001101101",
28318=>"000000111",
28319=>"101000000",
28320=>"101001011",
28321=>"110111111",
28322=>"100000100",
28323=>"000000000",
28324=>"000000011",
28325=>"001001110",
28326=>"110000001",
28327=>"000000000",
28328=>"010011111",
28329=>"000000000",
28330=>"101101101",
28331=>"111001110",
28332=>"111110100",
28333=>"111000101",
28334=>"111111110",
28335=>"010001011",
28336=>"000000100",
28337=>"001101010",
28338=>"110111111",
28339=>"000100110",
28340=>"011101111",
28341=>"000000101",
28342=>"000110000",
28343=>"100000000",
28344=>"001011000",
28345=>"100110111",
28346=>"111011101",
28347=>"111110110",
28348=>"000101001",
28349=>"011111111",
28350=>"001100000",
28351=>"000000000",
28352=>"000000000",
28353=>"000000000",
28354=>"010000111",
28355=>"100000000",
28356=>"000000011",
28357=>"111110100",
28358=>"010111111",
28359=>"011111010",
28360=>"111100001",
28361=>"011011010",
28362=>"111000001",
28363=>"001000011",
28364=>"110110010",
28365=>"110111111",
28366=>"111111010",
28367=>"001010010",
28368=>"000000100",
28369=>"111111111",
28370=>"101000100",
28371=>"111111111",
28372=>"000100101",
28373=>"000010001",
28374=>"101000000",
28375=>"000010111",
28376=>"000000000",
28377=>"000000000",
28378=>"101001010",
28379=>"100100101",
28380=>"111111110",
28381=>"100000101",
28382=>"111111111",
28383=>"000000001",
28384=>"010111010",
28385=>"100111111",
28386=>"101101111",
28387=>"101101101",
28388=>"000100000",
28389=>"101000101",
28390=>"000000000",
28391=>"111111111",
28392=>"100101001",
28393=>"000100011",
28394=>"010011011",
28395=>"001000000",
28396=>"000000000",
28397=>"000000010",
28398=>"110000000",
28399=>"100000000",
28400=>"001000000",
28401=>"111011011",
28402=>"010000011",
28403=>"000011011",
28404=>"000101111",
28405=>"000111111",
28406=>"000000000",
28407=>"111101111",
28408=>"000101111",
28409=>"001111111",
28410=>"000100100",
28411=>"111100100",
28412=>"011011001",
28413=>"000111111",
28414=>"011001001",
28415=>"100000000",
28416=>"111001100",
28417=>"001000111",
28418=>"000011011",
28419=>"000001000",
28420=>"111111111",
28421=>"101001100",
28422=>"010010000",
28423=>"000011111",
28424=>"111100000",
28425=>"001000010",
28426=>"001011110",
28427=>"011111101",
28428=>"000000000",
28429=>"111100000",
28430=>"110111111",
28431=>"000010111",
28432=>"000000000",
28433=>"000111111",
28434=>"111110010",
28435=>"000100111",
28436=>"010010000",
28437=>"000010111",
28438=>"111111111",
28439=>"111010011",
28440=>"000000000",
28441=>"111000000",
28442=>"001000000",
28443=>"011011010",
28444=>"001001000",
28445=>"000101000",
28446=>"000111100",
28447=>"000000001",
28448=>"111000010",
28449=>"111000111",
28450=>"010000000",
28451=>"111111111",
28452=>"011011011",
28453=>"000001000",
28454=>"110111000",
28455=>"111000111",
28456=>"100000101",
28457=>"100100010",
28458=>"111000000",
28459=>"001101111",
28460=>"010000110",
28461=>"000000100",
28462=>"011000100",
28463=>"000010000",
28464=>"000000010",
28465=>"010111111",
28466=>"111000010",
28467=>"011111111",
28468=>"101111001",
28469=>"000010101",
28470=>"111111011",
28471=>"111111000",
28472=>"001111101",
28473=>"111111010",
28474=>"000000001",
28475=>"111111000",
28476=>"000001001",
28477=>"111111000",
28478=>"001000000",
28479=>"001111011",
28480=>"110111000",
28481=>"000000010",
28482=>"111111111",
28483=>"100100100",
28484=>"101000001",
28485=>"100101111",
28486=>"010111000",
28487=>"001000101",
28488=>"000000110",
28489=>"000001111",
28490=>"110000000",
28491=>"000010000",
28492=>"000000000",
28493=>"110011110",
28494=>"110111010",
28495=>"000010111",
28496=>"110000000",
28497=>"111111110",
28498=>"000000000",
28499=>"001100111",
28500=>"000000000",
28501=>"001011111",
28502=>"111100100",
28503=>"101000001",
28504=>"000000001",
28505=>"100101010",
28506=>"001011011",
28507=>"110110110",
28508=>"011010000",
28509=>"100000011",
28510=>"001111000",
28511=>"101001001",
28512=>"100100000",
28513=>"000101101",
28514=>"000000101",
28515=>"110110110",
28516=>"000111010",
28517=>"000000111",
28518=>"010000000",
28519=>"010010110",
28520=>"101110000",
28521=>"001001101",
28522=>"111111111",
28523=>"000000101",
28524=>"000100110",
28525=>"111011011",
28526=>"000000000",
28527=>"001001111",
28528=>"010000001",
28529=>"111111100",
28530=>"111110110",
28531=>"000000101",
28532=>"111000000",
28533=>"000100101",
28534=>"000111111",
28535=>"111111111",
28536=>"111111011",
28537=>"111000000",
28538=>"111000000",
28539=>"000101101",
28540=>"101000010",
28541=>"100001101",
28542=>"011010011",
28543=>"000000000",
28544=>"011100110",
28545=>"000000000",
28546=>"011111110",
28547=>"001110111",
28548=>"000000110",
28549=>"001101101",
28550=>"000000000",
28551=>"111000110",
28552=>"000101000",
28553=>"101101000",
28554=>"000011011",
28555=>"000101111",
28556=>"000000000",
28557=>"000000000",
28558=>"000111001",
28559=>"001000000",
28560=>"001011111",
28561=>"000011111",
28562=>"111100111",
28563=>"101101111",
28564=>"100010000",
28565=>"001111111",
28566=>"001000000",
28567=>"100010010",
28568=>"000000111",
28569=>"101100111",
28570=>"101101110",
28571=>"011111010",
28572=>"100100111",
28573=>"110000100",
28574=>"111000000",
28575=>"000000000",
28576=>"100011101",
28577=>"111111111",
28578=>"000001111",
28579=>"111111001",
28580=>"011000111",
28581=>"010011111",
28582=>"001000101",
28583=>"101110110",
28584=>"000111111",
28585=>"000000100",
28586=>"111111101",
28587=>"111111111",
28588=>"001101101",
28589=>"010101111",
28590=>"111011010",
28591=>"011111101",
28592=>"000111000",
28593=>"111000101",
28594=>"001111001",
28595=>"011100000",
28596=>"001011111",
28597=>"111111111",
28598=>"100111111",
28599=>"001000000",
28600=>"000110100",
28601=>"101011100",
28602=>"101100000",
28603=>"101000000",
28604=>"001101001",
28605=>"011100111",
28606=>"111011001",
28607=>"111000000",
28608=>"111111000",
28609=>"011111000",
28610=>"010111111",
28611=>"000110000",
28612=>"000000100",
28613=>"001001000",
28614=>"000101111",
28615=>"111000000",
28616=>"111111001",
28617=>"000001000",
28618=>"111111011",
28619=>"010111111",
28620=>"010111011",
28621=>"000001111",
28622=>"111000000",
28623=>"110100000",
28624=>"101010010",
28625=>"100110011",
28626=>"101100100",
28627=>"000000111",
28628=>"000000000",
28629=>"111000000",
28630=>"110111011",
28631=>"101100111",
28632=>"000000000",
28633=>"000000000",
28634=>"011010100",
28635=>"000000100",
28636=>"111110111",
28637=>"000000111",
28638=>"000000000",
28639=>"000000000",
28640=>"000111011",
28641=>"000000100",
28642=>"000000111",
28643=>"111110110",
28644=>"101000000",
28645=>"010110000",
28646=>"101111111",
28647=>"111110010",
28648=>"000000000",
28649=>"010000010",
28650=>"111110011",
28651=>"000000000",
28652=>"000000000",
28653=>"111001101",
28654=>"010011010",
28655=>"100000100",
28656=>"000000100",
28657=>"100100100",
28658=>"001001100",
28659=>"010111111",
28660=>"110010001",
28661=>"111111101",
28662=>"000000101",
28663=>"100000111",
28664=>"111000000",
28665=>"111011111",
28666=>"101000000",
28667=>"010010000",
28668=>"111111011",
28669=>"110000011",
28670=>"101111001",
28671=>"110111111",
28672=>"100100111",
28673=>"000000111",
28674=>"101000000",
28675=>"000010111",
28676=>"000011011",
28677=>"101000001",
28678=>"100000110",
28679=>"001000000",
28680=>"000101000",
28681=>"101101001",
28682=>"110011011",
28683=>"000000000",
28684=>"010000101",
28685=>"000100101",
28686=>"010000010",
28687=>"110001000",
28688=>"010010000",
28689=>"000000110",
28690=>"101000111",
28691=>"000000000",
28692=>"000011111",
28693=>"111000000",
28694=>"000000011",
28695=>"001111111",
28696=>"000101110",
28697=>"000000110",
28698=>"001001001",
28699=>"000111000",
28700=>"110101111",
28701=>"111111011",
28702=>"011011011",
28703=>"110000000",
28704=>"100111111",
28705=>"000010000",
28706=>"110110000",
28707=>"101101111",
28708=>"111001001",
28709=>"000001111",
28710=>"000000111",
28711=>"110111111",
28712=>"011000000",
28713=>"000000110",
28714=>"101000001",
28715=>"011001100",
28716=>"000111111",
28717=>"111101101",
28718=>"111001111",
28719=>"100010001",
28720=>"111100000",
28721=>"010011011",
28722=>"111111001",
28723=>"000010010",
28724=>"000011111",
28725=>"000110111",
28726=>"100000011",
28727=>"111101101",
28728=>"000000100",
28729=>"111111101",
28730=>"001000000",
28731=>"101111010",
28732=>"111011111",
28733=>"111111111",
28734=>"001000111",
28735=>"100111111",
28736=>"011000100",
28737=>"001000000",
28738=>"000100101",
28739=>"011001111",
28740=>"000011010",
28741=>"111100000",
28742=>"000000000",
28743=>"010000000",
28744=>"111111001",
28745=>"000111111",
28746=>"111000000",
28747=>"101101001",
28748=>"101001111",
28749=>"111101000",
28750=>"001110110",
28751=>"010010111",
28752=>"000000001",
28753=>"111001000",
28754=>"110101111",
28755=>"010011011",
28756=>"100010000",
28757=>"000111110",
28758=>"010100100",
28759=>"000110010",
28760=>"110000000",
28761=>"000010011",
28762=>"110000011",
28763=>"001000000",
28764=>"111000001",
28765=>"110000000",
28766=>"111111111",
28767=>"001001101",
28768=>"010111111",
28769=>"111000001",
28770=>"100101111",
28771=>"100000110",
28772=>"001011001",
28773=>"100100011",
28774=>"010101111",
28775=>"110111111",
28776=>"111111000",
28777=>"100011000",
28778=>"010111111",
28779=>"111000000",
28780=>"111000110",
28781=>"010111110",
28782=>"111000000",
28783=>"000100000",
28784=>"000000011",
28785=>"000000000",
28786=>"001010110",
28787=>"110110011",
28788=>"111111111",
28789=>"001000000",
28790=>"111010000",
28791=>"000111111",
28792=>"000010111",
28793=>"100111111",
28794=>"000111111",
28795=>"110111000",
28796=>"110010110",
28797=>"010101000",
28798=>"000111000",
28799=>"001001011",
28800=>"000100000",
28801=>"010101001",
28802=>"000111111",
28803=>"010110000",
28804=>"001001010",
28805=>"000000010",
28806=>"100100110",
28807=>"101001011",
28808=>"100101000",
28809=>"111011011",
28810=>"000000000",
28811=>"111000000",
28812=>"111111000",
28813=>"000000000",
28814=>"000000000",
28815=>"101000000",
28816=>"111111011",
28817=>"110000100",
28818=>"001011000",
28819=>"101011111",
28820=>"101000100",
28821=>"000000000",
28822=>"110111101",
28823=>"010110100",
28824=>"111111111",
28825=>"000000000",
28826=>"111000000",
28827=>"000100011",
28828=>"111110100",
28829=>"111101100",
28830=>"001010100",
28831=>"000111111",
28832=>"011011101",
28833=>"011010000",
28834=>"011000000",
28835=>"110010111",
28836=>"101111111",
28837=>"000000100",
28838=>"000001001",
28839=>"111000001",
28840=>"000101111",
28841=>"000111111",
28842=>"111100000",
28843=>"011000110",
28844=>"101000001",
28845=>"001001001",
28846=>"110011011",
28847=>"110111111",
28848=>"111110000",
28849=>"111111101",
28850=>"000101101",
28851=>"110000100",
28852=>"011000001",
28853=>"000011011",
28854=>"010101011",
28855=>"000010000",
28856=>"111110111",
28857=>"000000110",
28858=>"010000111",
28859=>"001000011",
28860=>"111100111",
28861=>"111101101",
28862=>"001111111",
28863=>"000110111",
28864=>"000010111",
28865=>"111000000",
28866=>"111000101",
28867=>"110110110",
28868=>"000111011",
28869=>"100110110",
28870=>"000000001",
28871=>"000000000",
28872=>"111111110",
28873=>"010110000",
28874=>"000110010",
28875=>"111001000",
28876=>"000111011",
28877=>"001000101",
28878=>"001000110",
28879=>"100110111",
28880=>"000111111",
28881=>"010011001",
28882=>"001010110",
28883=>"110000000",
28884=>"111111011",
28885=>"011001010",
28886=>"100000001",
28887=>"000000000",
28888=>"100111000",
28889=>"010111001",
28890=>"010101100",
28891=>"000000001",
28892=>"000000110",
28893=>"110000000",
28894=>"011000000",
28895=>"000000001",
28896=>"000010010",
28897=>"011000000",
28898=>"111111111",
28899=>"000110110",
28900=>"100111110",
28901=>"000010111",
28902=>"001000101",
28903=>"110100100",
28904=>"111001001",
28905=>"111111111",
28906=>"000110110",
28907=>"000110111",
28908=>"000000000",
28909=>"101000110",
28910=>"111101101",
28911=>"100111101",
28912=>"100111000",
28913=>"101001001",
28914=>"000000111",
28915=>"000110111",
28916=>"101011111",
28917=>"111001001",
28918=>"111000000",
28919=>"000010000",
28920=>"000010000",
28921=>"111111001",
28922=>"111111100",
28923=>"000000111",
28924=>"100000000",
28925=>"000010000",
28926=>"011111110",
28927=>"111000000",
28928=>"000000000",
28929=>"000000010",
28930=>"111101101",
28931=>"110000000",
28932=>"001100100",
28933=>"011101101",
28934=>"000111000",
28935=>"111010010",
28936=>"011101100",
28937=>"000100101",
28938=>"110101111",
28939=>"000011111",
28940=>"000000000",
28941=>"111101111",
28942=>"011000010",
28943=>"010011000",
28944=>"000110110",
28945=>"011000100",
28946=>"100100110",
28947=>"000101101",
28948=>"100101001",
28949=>"101111100",
28950=>"001001010",
28951=>"001000001",
28952=>"101001000",
28953=>"101110111",
28954=>"010101010",
28955=>"000000111",
28956=>"100000000",
28957=>"000011010",
28958=>"010000100",
28959=>"000010010",
28960=>"111001101",
28961=>"111101111",
28962=>"101110101",
28963=>"001010000",
28964=>"101000001",
28965=>"001001100",
28966=>"010000101",
28967=>"000000111",
28968=>"111101111",
28969=>"011100111",
28970=>"000000000",
28971=>"100001000",
28972=>"100111111",
28973=>"111111111",
28974=>"010111101",
28975=>"111111000",
28976=>"111111101",
28977=>"101100001",
28978=>"111111111",
28979=>"111001101",
28980=>"010000011",
28981=>"000111001",
28982=>"011110100",
28983=>"101100101",
28984=>"001111101",
28985=>"111101101",
28986=>"000101000",
28987=>"000111111",
28988=>"110110011",
28989=>"110111111",
28990=>"101101101",
28991=>"011000101",
28992=>"101101101",
28993=>"000111101",
28994=>"110011001",
28995=>"010000000",
28996=>"010101001",
28997=>"000100101",
28998=>"000100101",
28999=>"100111111",
29000=>"111111111",
29001=>"010000010",
29002=>"111101101",
29003=>"011101111",
29004=>"010000000",
29005=>"111000000",
29006=>"111100000",
29007=>"101111111",
29008=>"000000000",
29009=>"110111111",
29010=>"100000101",
29011=>"010011001",
29012=>"000000000",
29013=>"100010110",
29014=>"000001110",
29015=>"101100101",
29016=>"011100110",
29017=>"100010110",
29018=>"010000011",
29019=>"000000100",
29020=>"111101101",
29021=>"010000010",
29022=>"111111011",
29023=>"100000000",
29024=>"011111000",
29025=>"100101010",
29026=>"110101101",
29027=>"001001111",
29028=>"110100000",
29029=>"000010111",
29030=>"111110111",
29031=>"101100000",
29032=>"100101000",
29033=>"111110100",
29034=>"111000101",
29035=>"111111001",
29036=>"000011001",
29037=>"111101111",
29038=>"001000100",
29039=>"000111110",
29040=>"101001001",
29041=>"000001000",
29042=>"000001001",
29043=>"000000111",
29044=>"111111101",
29045=>"000000001",
29046=>"110000001",
29047=>"010111111",
29048=>"110111110",
29049=>"001111110",
29050=>"111000000",
29051=>"111010100",
29052=>"011100000",
29053=>"010110110",
29054=>"000000010",
29055=>"111101000",
29056=>"010011101",
29057=>"111111001",
29058=>"111000101",
29059=>"011110101",
29060=>"000000000",
29061=>"111111111",
29062=>"100101011",
29063=>"111001110",
29064=>"101111110",
29065=>"111001110",
29066=>"000000111",
29067=>"111111101",
29068=>"000101101",
29069=>"111100010",
29070=>"000010000",
29071=>"000000001",
29072=>"011001010",
29073=>"000110111",
29074=>"000010111",
29075=>"011111111",
29076=>"000101000",
29077=>"111100101",
29078=>"000010111",
29079=>"100100000",
29080=>"101111111",
29081=>"111010001",
29082=>"100100100",
29083=>"111100000",
29084=>"010000100",
29085=>"111000000",
29086=>"011000100",
29087=>"010000011",
29088=>"100111011",
29089=>"111100011",
29090=>"000011011",
29091=>"000000101",
29092=>"111000111",
29093=>"111110001",
29094=>"101000101",
29095=>"110101111",
29096=>"000011001",
29097=>"110000000",
29098=>"111101101",
29099=>"111000000",
29100=>"001110101",
29101=>"010101010",
29102=>"001001010",
29103=>"100101110",
29104=>"000101111",
29105=>"100111011",
29106=>"111111100",
29107=>"001001001",
29108=>"000011111",
29109=>"110011000",
29110=>"000011011",
29111=>"011000010",
29112=>"000011010",
29113=>"001101001",
29114=>"010010011",
29115=>"000111111",
29116=>"101011000",
29117=>"111111001",
29118=>"010000000",
29119=>"100101000",
29120=>"010111111",
29121=>"111101100",
29122=>"111100100",
29123=>"110000100",
29124=>"100010110",
29125=>"010011010",
29126=>"000000100",
29127=>"111100110",
29128=>"000000111",
29129=>"111101100",
29130=>"110010100",
29131=>"001001001",
29132=>"111111110",
29133=>"100100011",
29134=>"000100011",
29135=>"111101101",
29136=>"111010001",
29137=>"000111010",
29138=>"100110100",
29139=>"000010000",
29140=>"111000111",
29141=>"001110110",
29142=>"001000010",
29143=>"000110111",
29144=>"000011111",
29145=>"011100100",
29146=>"111111110",
29147=>"101100000",
29148=>"100000000",
29149=>"111101000",
29150=>"000010010",
29151=>"110101101",
29152=>"111101001",
29153=>"011101010",
29154=>"101000000",
29155=>"000001011",
29156=>"010000000",
29157=>"101111011",
29158=>"111000000",
29159=>"000100000",
29160=>"011101001",
29161=>"101000000",
29162=>"111000011",
29163=>"010010111",
29164=>"111100101",
29165=>"111000101",
29166=>"000000111",
29167=>"000110010",
29168=>"000010111",
29169=>"110111110",
29170=>"000000000",
29171=>"000110111",
29172=>"010000000",
29173=>"011000000",
29174=>"010000100",
29175=>"000010010",
29176=>"111100100",
29177=>"000000001",
29178=>"111111000",
29179=>"011110000",
29180=>"110000000",
29181=>"000111001",
29182=>"110111111",
29183=>"111101111",
29184=>"101001000",
29185=>"000011011",
29186=>"000000000",
29187=>"000011111",
29188=>"101101100",
29189=>"011011001",
29190=>"010001000",
29191=>"010011110",
29192=>"001001011",
29193=>"011001001",
29194=>"010011001",
29195=>"010111000",
29196=>"001001001",
29197=>"111110100",
29198=>"101001101",
29199=>"010100110",
29200=>"111011001",
29201=>"000001001",
29202=>"101100101",
29203=>"101011011",
29204=>"010001000",
29205=>"111111111",
29206=>"100101110",
29207=>"100111111",
29208=>"001001000",
29209=>"011011111",
29210=>"011011101",
29211=>"010011011",
29212=>"000100100",
29213=>"111010110",
29214=>"011001001",
29215=>"000010110",
29216=>"000000000",
29217=>"001000011",
29218=>"000100110",
29219=>"000001011",
29220=>"011111110",
29221=>"000000010",
29222=>"001001111",
29223=>"000001000",
29224=>"111110110",
29225=>"000001011",
29226=>"000000101",
29227=>"110110010",
29228=>"111100100",
29229=>"001001001",
29230=>"011010001",
29231=>"100110000",
29232=>"001011111",
29233=>"000000011",
29234=>"000000011",
29235=>"011001001",
29236=>"000001001",
29237=>"000000000",
29238=>"000000000",
29239=>"101001001",
29240=>"011111000",
29241=>"011011011",
29242=>"100100100",
29243=>"011011000",
29244=>"011001111",
29245=>"110110110",
29246=>"000000001",
29247=>"011011000",
29248=>"111011001",
29249=>"011001011",
29250=>"000111010",
29251=>"101000011",
29252=>"011010000",
29253=>"001101000",
29254=>"100011000",
29255=>"000100111",
29256=>"100000110",
29257=>"110111111",
29258=>"111101111",
29259=>"001101001",
29260=>"001000100",
29261=>"001001001",
29262=>"000001001",
29263=>"000000000",
29264=>"000000000",
29265=>"110000110",
29266=>"111111011",
29267=>"010000010",
29268=>"000011110",
29269=>"010000000",
29270=>"100110111",
29271=>"011011000",
29272=>"000000111",
29273=>"010000011",
29274=>"010110110",
29275=>"101101111",
29276=>"011011001",
29277=>"000010111",
29278=>"001011001",
29279=>"010010000",
29280=>"000010010",
29281=>"110110000",
29282=>"011010000",
29283=>"100101100",
29284=>"000010110",
29285=>"000111100",
29286=>"111000111",
29287=>"001000110",
29288=>"011011111",
29289=>"010001001",
29290=>"110110011",
29291=>"010011111",
29292=>"110101111",
29293=>"110110100",
29294=>"001000000",
29295=>"000000100",
29296=>"101000001",
29297=>"011111111",
29298=>"001010001",
29299=>"000000000",
29300=>"011000010",
29301=>"001001001",
29302=>"000011011",
29303=>"111100001",
29304=>"000000000",
29305=>"010100110",
29306=>"000100110",
29307=>"111011111",
29308=>"111011000",
29309=>"111001000",
29310=>"100110111",
29311=>"000110110",
29312=>"001001001",
29313=>"110110011",
29314=>"001001011",
29315=>"001000000",
29316=>"111111110",
29317=>"100110000",
29318=>"011110100",
29319=>"100100100",
29320=>"011011010",
29321=>"100110111",
29322=>"011111001",
29323=>"000001000",
29324=>"001111011",
29325=>"111111000",
29326=>"011000011",
29327=>"000001011",
29328=>"101100101",
29329=>"111101110",
29330=>"000000001",
29331=>"000111011",
29332=>"000101111",
29333=>"001001001",
29334=>"001000010",
29335=>"101100100",
29336=>"000010101",
29337=>"000000111",
29338=>"001000010",
29339=>"001000010",
29340=>"001101111",
29341=>"000000000",
29342=>"000111001",
29343=>"100100001",
29344=>"100000001",
29345=>"011111011",
29346=>"000010110",
29347=>"000000001",
29348=>"110011011",
29349=>"101001111",
29350=>"011111010",
29351=>"100000110",
29352=>"001011001",
29353=>"001101101",
29354=>"101001001",
29355=>"000001000",
29356=>"001111100",
29357=>"101000000",
29358=>"010010000",
29359=>"011010001",
29360=>"011001001",
29361=>"110011001",
29362=>"000000000",
29363=>"000001011",
29364=>"010011011",
29365=>"010100010",
29366=>"101000101",
29367=>"010011000",
29368=>"100100100",
29369=>"010010010",
29370=>"001000110",
29371=>"011110111",
29372=>"110110100",
29373=>"100110110",
29374=>"100010000",
29375=>"000001010",
29376=>"001001001",
29377=>"011000001",
29378=>"011111111",
29379=>"000011010",
29380=>"000001111",
29381=>"000110010",
29382=>"110100111",
29383=>"011000111",
29384=>"100000110",
29385=>"111010010",
29386=>"110000011",
29387=>"000100101",
29388=>"100101101",
29389=>"000000000",
29390=>"001001001",
29391=>"111101100",
29392=>"101000000",
29393=>"100100110",
29394=>"111001001",
29395=>"110110110",
29396=>"001001111",
29397=>"100110110",
29398=>"000011000",
29399=>"011111001",
29400=>"000010010",
29401=>"110010110",
29402=>"011000000",
29403=>"001001001",
29404=>"011111111",
29405=>"100100111",
29406=>"111111111",
29407=>"000111011",
29408=>"000000001",
29409=>"001001001",
29410=>"100110111",
29411=>"110110011",
29412=>"001001001",
29413=>"110110110",
29414=>"111111010",
29415=>"101111010",
29416=>"000100111",
29417=>"100010000",
29418=>"001111101",
29419=>"011011000",
29420=>"001000011",
29421=>"001111110",
29422=>"100000100",
29423=>"000100111",
29424=>"000000000",
29425=>"101100101",
29426=>"001001001",
29427=>"101101100",
29428=>"011000001",
29429=>"100110110",
29430=>"000001110",
29431=>"110110100",
29432=>"001001001",
29433=>"001111010",
29434=>"101100001",
29435=>"111110110",
29436=>"111111111",
29437=>"110110111",
29438=>"001110110",
29439=>"001111000",
29440=>"110110011",
29441=>"001001001",
29442=>"111000000",
29443=>"111010000",
29444=>"001000001",
29445=>"000000000",
29446=>"110010010",
29447=>"010000010",
29448=>"000000000",
29449=>"000110010",
29450=>"001011000",
29451=>"000110100",
29452=>"001000111",
29453=>"000000000",
29454=>"100111011",
29455=>"111111101",
29456=>"001000000",
29457=>"110110011",
29458=>"111000000",
29459=>"000000011",
29460=>"111111010",
29461=>"000100111",
29462=>"100100100",
29463=>"010000000",
29464=>"000000000",
29465=>"000000110",
29466=>"100101011",
29467=>"011000111",
29468=>"100101000",
29469=>"001100000",
29470=>"111110000",
29471=>"101101000",
29472=>"000111100",
29473=>"011011000",
29474=>"110111111",
29475=>"101101000",
29476=>"001001000",
29477=>"000100110",
29478=>"100101111",
29479=>"101111101",
29480=>"101010111",
29481=>"111101101",
29482=>"110111101",
29483=>"111111001",
29484=>"011111111",
29485=>"011100111",
29486=>"111111111",
29487=>"110100000",
29488=>"000011011",
29489=>"010101001",
29490=>"000011010",
29491=>"000111111",
29492=>"001101111",
29493=>"000111000",
29494=>"001001001",
29495=>"000111110",
29496=>"001010111",
29497=>"010000011",
29498=>"011001000",
29499=>"000000101",
29500=>"001001001",
29501=>"111101000",
29502=>"000010001",
29503=>"010110001",
29504=>"101111000",
29505=>"100111011",
29506=>"111000111",
29507=>"001001001",
29508=>"101001011",
29509=>"000000000",
29510=>"000000000",
29511=>"010011010",
29512=>"001001100",
29513=>"000110110",
29514=>"000010110",
29515=>"000110001",
29516=>"001101011",
29517=>"000001001",
29518=>"000000001",
29519=>"011111101",
29520=>"111000000",
29521=>"000000000",
29522=>"000001111",
29523=>"011011101",
29524=>"101000000",
29525=>"101101000",
29526=>"010000001",
29527=>"111111010",
29528=>"111111101",
29529=>"010100101",
29530=>"011001000",
29531=>"000011011",
29532=>"001000000",
29533=>"010011001",
29534=>"000011111",
29535=>"001110100",
29536=>"101111111",
29537=>"111010111",
29538=>"101001000",
29539=>"110010000",
29540=>"010010100",
29541=>"111101111",
29542=>"011011000",
29543=>"011110000",
29544=>"000011111",
29545=>"110110110",
29546=>"010001000",
29547=>"001110010",
29548=>"111101010",
29549=>"110010011",
29550=>"111111010",
29551=>"000000010",
29552=>"000001000",
29553=>"000000111",
29554=>"100100100",
29555=>"000001000",
29556=>"100111000",
29557=>"111010111",
29558=>"111111110",
29559=>"000000000",
29560=>"111011010",
29561=>"011101101",
29562=>"000001101",
29563=>"000111111",
29564=>"000110100",
29565=>"110110001",
29566=>"101111010",
29567=>"000000110",
29568=>"000000101",
29569=>"000000000",
29570=>"111100000",
29571=>"111111001",
29572=>"101001000",
29573=>"000110010",
29574=>"001001011",
29575=>"110000000",
29576=>"001001001",
29577=>"110000110",
29578=>"010010111",
29579=>"000000000",
29580=>"000101111",
29581=>"011111011",
29582=>"010001001",
29583=>"000000000",
29584=>"000100101",
29585=>"101111111",
29586=>"000110111",
29587=>"111111101",
29588=>"000000011",
29589=>"001000000",
29590=>"111111001",
29591=>"000000001",
29592=>"011010011",
29593=>"001001111",
29594=>"101001111",
29595=>"000110000",
29596=>"010110000",
29597=>"001001101",
29598=>"001110000",
29599=>"111100001",
29600=>"101100100",
29601=>"000101111",
29602=>"101111111",
29603=>"000000000",
29604=>"100110011",
29605=>"100100100",
29606=>"000000100",
29607=>"100111100",
29608=>"111000100",
29609=>"000101101",
29610=>"111101110",
29611=>"111101000",
29612=>"001000000",
29613=>"000000001",
29614=>"011011001",
29615=>"010011110",
29616=>"000100000",
29617=>"011010000",
29618=>"000011111",
29619=>"011001000",
29620=>"000001001",
29621=>"001101000",
29622=>"000010011",
29623=>"000110111",
29624=>"100100100",
29625=>"000100110",
29626=>"000100101",
29627=>"010110010",
29628=>"111111111",
29629=>"110010010",
29630=>"000100010",
29631=>"101011111",
29632=>"001101011",
29633=>"111011000",
29634=>"010000010",
29635=>"001011001",
29636=>"000000011",
29637=>"110110101",
29638=>"001000000",
29639=>"110111110",
29640=>"111000000",
29641=>"100000111",
29642=>"000110010",
29643=>"101000111",
29644=>"100111010",
29645=>"001011000",
29646=>"111101001",
29647=>"011111001",
29648=>"011101111",
29649=>"000000011",
29650=>"000000110",
29651=>"101101110",
29652=>"111000110",
29653=>"111010000",
29654=>"111111001",
29655=>"110111100",
29656=>"000000111",
29657=>"000000000",
29658=>"111011011",
29659=>"000000110",
29660=>"001001001",
29661=>"001000000",
29662=>"001111111",
29663=>"011111110",
29664=>"000000000",
29665=>"101001111",
29666=>"101101111",
29667=>"011111101",
29668=>"000000000",
29669=>"101010000",
29670=>"000000010",
29671=>"100100100",
29672=>"010110010",
29673=>"110111101",
29674=>"100110000",
29675=>"111111011",
29676=>"000000110",
29677=>"000000111",
29678=>"100000010",
29679=>"001000111",
29680=>"001101001",
29681=>"101111101",
29682=>"101101111",
29683=>"111111001",
29684=>"011001110",
29685=>"010110101",
29686=>"010000000",
29687=>"011111111",
29688=>"101001000",
29689=>"101101111",
29690=>"011111000",
29691=>"010000101",
29692=>"010111101",
29693=>"001000000",
29694=>"010000100",
29695=>"111111000",
29696=>"000000011",
29697=>"100000000",
29698=>"010010000",
29699=>"010000011",
29700=>"100101111",
29701=>"110110000",
29702=>"111011111",
29703=>"000010110",
29704=>"000001101",
29705=>"000111111",
29706=>"100100101",
29707=>"101110110",
29708=>"111001000",
29709=>"110111000",
29710=>"000011010",
29711=>"000010000",
29712=>"000001000",
29713=>"000010000",
29714=>"000000000",
29715=>"101111111",
29716=>"001100010",
29717=>"000110010",
29718=>"010000000",
29719=>"001011110",
29720=>"000000000",
29721=>"101001111",
29722=>"001001111",
29723=>"000000000",
29724=>"000000111",
29725=>"101001111",
29726=>"000000000",
29727=>"000001111",
29728=>"111000000",
29729=>"000101000",
29730=>"000000000",
29731=>"000000000",
29732=>"101111111",
29733=>"001000110",
29734=>"111010000",
29735=>"111000011",
29736=>"010111111",
29737=>"000100110",
29738=>"110111101",
29739=>"111111111",
29740=>"001001111",
29741=>"000000011",
29742=>"101001000",
29743=>"010001001",
29744=>"010000101",
29745=>"111111111",
29746=>"000101000",
29747=>"000000000",
29748=>"111110011",
29749=>"111010110",
29750=>"110001001",
29751=>"000111111",
29752=>"111000000",
29753=>"000000000",
29754=>"001000000",
29755=>"111000000",
29756=>"101111111",
29757=>"111111000",
29758=>"000000010",
29759=>"110110110",
29760=>"001000000",
29761=>"100101101",
29762=>"111000010",
29763=>"110111111",
29764=>"010000111",
29765=>"000001000",
29766=>"001101100",
29767=>"111111001",
29768=>"101111111",
29769=>"000001000",
29770=>"000000001",
29771=>"000000001",
29772=>"001011111",
29773=>"111011111",
29774=>"011111111",
29775=>"110000000",
29776=>"001100000",
29777=>"111000000",
29778=>"111000111",
29779=>"011001101",
29780=>"101000010",
29781=>"101100111",
29782=>"011011001",
29783=>"110111100",
29784=>"001011001",
29785=>"111101111",
29786=>"100100000",
29787=>"101101101",
29788=>"000000100",
29789=>"000000001",
29790=>"111111111",
29791=>"110111011",
29792=>"010110010",
29793=>"000000000",
29794=>"000000000",
29795=>"010111000",
29796=>"000000000",
29797=>"111101000",
29798=>"111001111",
29799=>"101111111",
29800=>"010000000",
29801=>"000101111",
29802=>"000000011",
29803=>"111111110",
29804=>"110000110",
29805=>"110010000",
29806=>"001001111",
29807=>"000100000",
29808=>"101011011",
29809=>"001101101",
29810=>"011100101",
29811=>"010000000",
29812=>"111111111",
29813=>"000000101",
29814=>"111111101",
29815=>"111111000",
29816=>"110111100",
29817=>"001000000",
29818=>"100000110",
29819=>"111001001",
29820=>"100000110",
29821=>"100000000",
29822=>"111000010",
29823=>"001001001",
29824=>"001000100",
29825=>"111101000",
29826=>"000100110",
29827=>"111101110",
29828=>"001000010",
29829=>"111001010",
29830=>"101101111",
29831=>"010001101",
29832=>"001001001",
29833=>"111100000",
29834=>"101000001",
29835=>"001000100",
29836=>"010111111",
29837=>"000000110",
29838=>"110111011",
29839=>"001000000",
29840=>"001001011",
29841=>"110010110",
29842=>"110000001",
29843=>"010100110",
29844=>"000010010",
29845=>"111111110",
29846=>"110011110",
29847=>"000001001",
29848=>"111111111",
29849=>"111101111",
29850=>"111111111",
29851=>"010000100",
29852=>"100111010",
29853=>"111111011",
29854=>"000010111",
29855=>"101000101",
29856=>"111100100",
29857=>"000000000",
29858=>"110111010",
29859=>"111101111",
29860=>"101000101",
29861=>"001001100",
29862=>"000000000",
29863=>"111101001",
29864=>"101010011",
29865=>"000000000",
29866=>"111001000",
29867=>"000000000",
29868=>"000001000",
29869=>"000110000",
29870=>"000000100",
29871=>"010001011",
29872=>"111110110",
29873=>"110100001",
29874=>"111111101",
29875=>"000000100",
29876=>"100100100",
29877=>"000000000",
29878=>"111111111",
29879=>"000101101",
29880=>"001011111",
29881=>"100100100",
29882=>"110110011",
29883=>"000000110",
29884=>"100111111",
29885=>"111111111",
29886=>"011011011",
29887=>"011000000",
29888=>"000010010",
29889=>"000000000",
29890=>"101110100",
29891=>"011101101",
29892=>"001111000",
29893=>"101000001",
29894=>"000000111",
29895=>"001000000",
29896=>"101111110",
29897=>"110010101",
29898=>"011111011",
29899=>"111011111",
29900=>"011111000",
29901=>"010011011",
29902=>"000000000",
29903=>"111111111",
29904=>"000000000",
29905=>"110000010",
29906=>"001001110",
29907=>"001011110",
29908=>"101010000",
29909=>"001000000",
29910=>"000000000",
29911=>"101111111",
29912=>"111111111",
29913=>"000100111",
29914=>"111001001",
29915=>"001000000",
29916=>"000000000",
29917=>"101001001",
29918=>"101111111",
29919=>"110000111",
29920=>"000000001",
29921=>"000000000",
29922=>"111111111",
29923=>"100000000",
29924=>"001000000",
29925=>"001000000",
29926=>"101111111",
29927=>"100010000",
29928=>"111111111",
29929=>"101000001",
29930=>"000000001",
29931=>"110010010",
29932=>"000000000",
29933=>"101111111",
29934=>"000000000",
29935=>"000000111",
29936=>"101111111",
29937=>"111011000",
29938=>"000000100",
29939=>"001001001",
29940=>"000000100",
29941=>"000000000",
29942=>"001000111",
29943=>"111111101",
29944=>"101100111",
29945=>"001010010",
29946=>"101111011",
29947=>"100010001",
29948=>"000000000",
29949=>"111111111",
29950=>"000000101",
29951=>"111110000",
29952=>"000001001",
29953=>"100111111",
29954=>"000000100",
29955=>"101101101",
29956=>"110011101",
29957=>"100010110",
29958=>"111011011",
29959=>"100111111",
29960=>"000000000",
29961=>"000000110",
29962=>"000000100",
29963=>"110100010",
29964=>"011000000",
29965=>"110010011",
29966=>"001001110",
29967=>"001101001",
29968=>"100000000",
29969=>"111000110",
29970=>"000000000",
29971=>"011000111",
29972=>"100100111",
29973=>"000011000",
29974=>"010110011",
29975=>"001001011",
29976=>"001101000",
29977=>"010100100",
29978=>"100000111",
29979=>"000000100",
29980=>"110000011",
29981=>"100111110",
29982=>"000010000",
29983=>"101101100",
29984=>"111100011",
29985=>"100110010",
29986=>"000010001",
29987=>"111111011",
29988=>"001001110",
29989=>"011100111",
29990=>"011000100",
29991=>"001100111",
29992=>"000000101",
29993=>"110010011",
29994=>"001100001",
29995=>"101100010",
29996=>"001111011",
29997=>"110111111",
29998=>"100101111",
29999=>"000100011",
30000=>"000111111",
30001=>"110010001",
30002=>"110110100",
30003=>"000011111",
30004=>"000000000",
30005=>"000111011",
30006=>"000001111",
30007=>"000011111",
30008=>"011111010",
30009=>"101000011",
30010=>"000100001",
30011=>"111011111",
30012=>"010001100",
30013=>"111111000",
30014=>"000000101",
30015=>"001100001",
30016=>"111111001",
30017=>"001000010",
30018=>"011011001",
30019=>"110000100",
30020=>"011011000",
30021=>"000010101",
30022=>"000100111",
30023=>"011111110",
30024=>"001111111",
30025=>"000000011",
30026=>"101100101",
30027=>"111100111",
30028=>"000000100",
30029=>"110110011",
30030=>"011001010",
30031=>"011111111",
30032=>"000010111",
30033=>"000100100",
30034=>"001000000",
30035=>"000110110",
30036=>"110100000",
30037=>"111101100",
30038=>"010001011",
30039=>"111000110",
30040=>"000100100",
30041=>"110010000",
30042=>"110111110",
30043=>"001100000",
30044=>"011010000",
30045=>"000000101",
30046=>"011011000",
30047=>"001100100",
30048=>"011000000",
30049=>"000000110",
30050=>"111000000",
30051=>"100101001",
30052=>"100110011",
30053=>"100100011",
30054=>"000101111",
30055=>"000100111",
30056=>"000011000",
30057=>"100000000",
30058=>"110111000",
30059=>"000011110",
30060=>"111110100",
30061=>"101000111",
30062=>"000000001",
30063=>"011001111",
30064=>"110100111",
30065=>"100100110",
30066=>"100110110",
30067=>"011011000",
30068=>"111110001",
30069=>"000000011",
30070=>"100111000",
30071=>"011000000",
30072=>"000000000",
30073=>"011000101",
30074=>"100110000",
30075=>"111101011",
30076=>"100111111",
30077=>"100100111",
30078=>"111001000",
30079=>"000000100",
30080=>"001011011",
30081=>"000011111",
30082=>"011000011",
30083=>"001000010",
30084=>"000010111",
30085=>"001101011",
30086=>"010000001",
30087=>"010001000",
30088=>"101111000",
30089=>"100011011",
30090=>"100100011",
30091=>"100011000",
30092=>"001000111",
30093=>"000111111",
30094=>"001000000",
30095=>"000000000",
30096=>"110111111",
30097=>"000011001",
30098=>"000000010",
30099=>"010000000",
30100=>"001101010",
30101=>"001000100",
30102=>"011111000",
30103=>"001001011",
30104=>"100001111",
30105=>"001100000",
30106=>"000100111",
30107=>"000000110",
30108=>"011000011",
30109=>"000000011",
30110=>"000111011",
30111=>"101000100",
30112=>"000111111",
30113=>"100100111",
30114=>"000000111",
30115=>"100100000",
30116=>"100000000",
30117=>"000011110",
30118=>"100010000",
30119=>"011110110",
30120=>"111001111",
30121=>"111111111",
30122=>"111100111",
30123=>"011000000",
30124=>"101000011",
30125=>"000100100",
30126=>"001101100",
30127=>"111011011",
30128=>"000000011",
30129=>"000101110",
30130=>"000100110",
30131=>"100000000",
30132=>"110101100",
30133=>"111011111",
30134=>"011000001",
30135=>"011011000",
30136=>"101000000",
30137=>"110101101",
30138=>"000010000",
30139=>"011100000",
30140=>"111010001",
30141=>"111111101",
30142=>"110100100",
30143=>"000000111",
30144=>"000100101",
30145=>"100000000",
30146=>"001111011",
30147=>"110110001",
30148=>"000110110",
30149=>"010111111",
30150=>"110010110",
30151=>"001001111",
30152=>"111111011",
30153=>"011011000",
30154=>"000101010",
30155=>"111001100",
30156=>"000000100",
30157=>"011001010",
30158=>"000001000",
30159=>"111011000",
30160=>"111100100",
30161=>"111110100",
30162=>"010000001",
30163=>"000000000",
30164=>"000100111",
30165=>"100110111",
30166=>"101011001",
30167=>"100111111",
30168=>"111101011",
30169=>"011000100",
30170=>"111101111",
30171=>"001000111",
30172=>"111000110",
30173=>"111000100",
30174=>"011000000",
30175=>"000111110",
30176=>"011011000",
30177=>"000100000",
30178=>"100000000",
30179=>"010100111",
30180=>"111000000",
30181=>"001010000",
30182=>"111101011",
30183=>"100100111",
30184=>"011000010",
30185=>"101001000",
30186=>"010000001",
30187=>"111011000",
30188=>"011011000",
30189=>"011011011",
30190=>"000010000",
30191=>"111100100",
30192=>"100111011",
30193=>"000101001",
30194=>"011010000",
30195=>"001101101",
30196=>"100110110",
30197=>"000001011",
30198=>"000000000",
30199=>"100100111",
30200=>"000111010",
30201=>"000101011",
30202=>"100000111",
30203=>"100100010",
30204=>"111100001",
30205=>"101000000",
30206=>"000000001",
30207=>"100100011",
30208=>"000100000",
30209=>"001001010",
30210=>"100000000",
30211=>"000101101",
30212=>"110111011",
30213=>"001001101",
30214=>"101111111",
30215=>"111000000",
30216=>"000001001",
30217=>"100000000",
30218=>"100100111",
30219=>"000111111",
30220=>"101111111",
30221=>"000011111",
30222=>"100010101",
30223=>"111110111",
30224=>"100010111",
30225=>"111000111",
30226=>"010000110",
30227=>"111000000",
30228=>"101111001",
30229=>"000000110",
30230=>"110110101",
30231=>"110111011",
30232=>"000000000",
30233=>"100000000",
30234=>"001100100",
30235=>"000010111",
30236=>"000000011",
30237=>"010101000",
30238=>"101010000",
30239=>"001000101",
30240=>"111101111",
30241=>"110111111",
30242=>"001000000",
30243=>"000000000",
30244=>"110011100",
30245=>"100000000",
30246=>"111000111",
30247=>"111000101",
30248=>"111111000",
30249=>"101111011",
30250=>"100000101",
30251=>"111000000",
30252=>"101100010",
30253=>"111000110",
30254=>"101000000",
30255=>"111111111",
30256=>"000111111",
30257=>"011111001",
30258=>"111101111",
30259=>"100000000",
30260=>"111001000",
30261=>"000111111",
30262=>"110100011",
30263=>"000111111",
30264=>"110000000",
30265=>"000000001",
30266=>"001000000",
30267=>"111111111",
30268=>"001011101",
30269=>"000010001",
30270=>"000000101",
30271=>"000001101",
30272=>"101011111",
30273=>"111010010",
30274=>"000011110",
30275=>"000000000",
30276=>"111101000",
30277=>"000101011",
30278=>"000110011",
30279=>"111000111",
30280=>"000001101",
30281=>"000000100",
30282=>"101000000",
30283=>"000001011",
30284=>"111000001",
30285=>"111000000",
30286=>"111111110",
30287=>"000000001",
30288=>"100000000",
30289=>"000111001",
30290=>"100100000",
30291=>"100000000",
30292=>"000000000",
30293=>"011110111",
30294=>"111000000",
30295=>"110000010",
30296=>"101000001",
30297=>"111000001",
30298=>"101111111",
30299=>"010100100",
30300=>"000000000",
30301=>"100100000",
30302=>"111111111",
30303=>"100000000",
30304=>"111101101",
30305=>"000000000",
30306=>"000000000",
30307=>"110110111",
30308=>"000001101",
30309=>"011001011",
30310=>"000000000",
30311=>"000000000",
30312=>"001001000",
30313=>"111111011",
30314=>"111000000",
30315=>"000100011",
30316=>"011000110",
30317=>"111111100",
30318=>"000100111",
30319=>"010101111",
30320=>"100110000",
30321=>"000000111",
30322=>"011000110",
30323=>"111000000",
30324=>"011011111",
30325=>"100000000",
30326=>"110111111",
30327=>"000111101",
30328=>"101010101",
30329=>"111001001",
30330=>"110111110",
30331=>"111101000",
30332=>"001001001",
30333=>"001000000",
30334=>"111111111",
30335=>"000100000",
30336=>"001000100",
30337=>"000011011",
30338=>"000001111",
30339=>"001001100",
30340=>"000000010",
30341=>"010000000",
30342=>"010011000",
30343=>"000000100",
30344=>"001111110",
30345=>"011000100",
30346=>"111111000",
30347=>"100111111",
30348=>"011111000",
30349=>"000000000",
30350=>"111111111",
30351=>"101000101",
30352=>"001101001",
30353=>"111011111",
30354=>"010111111",
30355=>"000011101",
30356=>"000000100",
30357=>"000000000",
30358=>"111111100",
30359=>"110111111",
30360=>"111001000",
30361=>"001000000",
30362=>"010000001",
30363=>"110000111",
30364=>"000000000",
30365=>"010111000",
30366=>"001100101",
30367=>"111000111",
30368=>"110100011",
30369=>"111000101",
30370=>"001000011",
30371=>"000000000",
30372=>"101001101",
30373=>"011000001",
30374=>"101100111",
30375=>"111111101",
30376=>"000000000",
30377=>"111011101",
30378=>"000000000",
30379=>"111000000",
30380=>"000101110",
30381=>"000000000",
30382=>"101010110",
30383=>"001000010",
30384=>"000110111",
30385=>"100000110",
30386=>"100000011",
30387=>"000000100",
30388=>"100110001",
30389=>"010100111",
30390=>"111100100",
30391=>"011111101",
30392=>"000000000",
30393=>"010110001",
30394=>"101000000",
30395=>"000001111",
30396=>"000101010",
30397=>"011111010",
30398=>"111110101",
30399=>"111000000",
30400=>"000000001",
30401=>"000000111",
30402=>"110010110",
30403=>"011111111",
30404=>"111111111",
30405=>"001011111",
30406=>"110110011",
30407=>"111000001",
30408=>"111100110",
30409=>"000010110",
30410=>"101111111",
30411=>"100000000",
30412=>"100000000",
30413=>"000000000",
30414=>"111111111",
30415=>"010111101",
30416=>"001000001",
30417=>"111111001",
30418=>"000100111",
30419=>"111111100",
30420=>"000000000",
30421=>"001011011",
30422=>"000000000",
30423=>"000000111",
30424=>"111111111",
30425=>"011000000",
30426=>"011000000",
30427=>"111111000",
30428=>"000001111",
30429=>"111000001",
30430=>"111000100",
30431=>"000000111",
30432=>"000000100",
30433=>"000010010",
30434=>"000111111",
30435=>"111100000",
30436=>"000000101",
30437=>"101111011",
30438=>"000000111",
30439=>"011101001",
30440=>"111001000",
30441=>"111111011",
30442=>"111100111",
30443=>"000000001",
30444=>"011111111",
30445=>"111001110",
30446=>"000000000",
30447=>"100001111",
30448=>"011000010",
30449=>"000010110",
30450=>"000001011",
30451=>"001000001",
30452=>"101001000",
30453=>"010110111",
30454=>"100000000",
30455=>"000010111",
30456=>"110111000",
30457=>"111011011",
30458=>"000000000",
30459=>"111111111",
30460=>"111000101",
30461=>"001110111",
30462=>"000000000",
30463=>"110000000",
30464=>"011111100",
30465=>"010111111",
30466=>"000000101",
30467=>"101111000",
30468=>"000000010",
30469=>"000000000",
30470=>"000000010",
30471=>"111111111",
30472=>"111111111",
30473=>"111100000",
30474=>"111010100",
30475=>"101011001",
30476=>"001011000",
30477=>"000000000",
30478=>"000000100",
30479=>"111111110",
30480=>"111110101",
30481=>"101101000",
30482=>"111111111",
30483=>"111101000",
30484=>"110110010",
30485=>"111000001",
30486=>"000010110",
30487=>"110100001",
30488=>"100100111",
30489=>"100111001",
30490=>"000001011",
30491=>"111111111",
30492=>"110101010",
30493=>"000010000",
30494=>"111001011",
30495=>"110000000",
30496=>"000010110",
30497=>"111111000",
30498=>"111010001",
30499=>"000000000",
30500=>"100100101",
30501=>"111111011",
30502=>"000101011",
30503=>"001110010",
30504=>"111111111",
30505=>"111010111",
30506=>"000000000",
30507=>"001110000",
30508=>"000110000",
30509=>"111111000",
30510=>"010010000",
30511=>"001000010",
30512=>"000000110",
30513=>"101011011",
30514=>"101000011",
30515=>"111111000",
30516=>"000000010",
30517=>"110110010",
30518=>"001011011",
30519=>"111101100",
30520=>"110011011",
30521=>"000000001",
30522=>"011001001",
30523=>"100111111",
30524=>"111111011",
30525=>"111111111",
30526=>"000000000",
30527=>"000000110",
30528=>"010000101",
30529=>"101100101",
30530=>"001101111",
30531=>"010000001",
30532=>"111111111",
30533=>"010000000",
30534=>"010111110",
30535=>"010000000",
30536=>"111110001",
30537=>"011010011",
30538=>"000111111",
30539=>"011111011",
30540=>"000000101",
30541=>"000000110",
30542=>"000110111",
30543=>"111110111",
30544=>"110101111",
30545=>"111111110",
30546=>"111111111",
30547=>"111001001",
30548=>"110111011",
30549=>"111110100",
30550=>"111110101",
30551=>"110100111",
30552=>"100001000",
30553=>"011011000",
30554=>"000101011",
30555=>"000011011",
30556=>"000000111",
30557=>"001001011",
30558=>"111000111",
30559=>"111000100",
30560=>"110100000",
30561=>"111011110",
30562=>"000000000",
30563=>"000001101",
30564=>"000101111",
30565=>"100011010",
30566=>"010111011",
30567=>"111000110",
30568=>"010111111",
30569=>"010000000",
30570=>"000001110",
30571=>"010000100",
30572=>"110110111",
30573=>"001000000",
30574=>"010010000",
30575=>"000101111",
30576=>"000100110",
30577=>"000011101",
30578=>"110110110",
30579=>"110000111",
30580=>"111111000",
30581=>"100000011",
30582=>"000000000",
30583=>"110000000",
30584=>"111111000",
30585=>"000110010",
30586=>"111111111",
30587=>"101111111",
30588=>"110110101",
30589=>"100000000",
30590=>"101000100",
30591=>"100000110",
30592=>"000101000",
30593=>"111000000",
30594=>"100000000",
30595=>"001001111",
30596=>"111111111",
30597=>"101111111",
30598=>"100010000",
30599=>"001000000",
30600=>"000010110",
30601=>"000010101",
30602=>"111101110",
30603=>"010000000",
30604=>"111000111",
30605=>"000000000",
30606=>"111010111",
30607=>"001000100",
30608=>"000111111",
30609=>"111000010",
30610=>"000100111",
30611=>"001010000",
30612=>"000110000",
30613=>"011111000",
30614=>"000000101",
30615=>"111111111",
30616=>"010110011",
30617=>"111000000",
30618=>"101000001",
30619=>"011111110",
30620=>"111111100",
30621=>"111011110",
30622=>"111010000",
30623=>"000001000",
30624=>"100010000",
30625=>"001000111",
30626=>"000000000",
30627=>"001010011",
30628=>"000000000",
30629=>"100101100",
30630=>"110101011",
30631=>"000100010",
30632=>"011111110",
30633=>"011111101",
30634=>"101111110",
30635=>"111111101",
30636=>"000000010",
30637=>"010000111",
30638=>"101111101",
30639=>"000111010",
30640=>"000101111",
30641=>"011101101",
30642=>"001000000",
30643=>"101101111",
30644=>"000011011",
30645=>"000000010",
30646=>"010000011",
30647=>"010000000",
30648=>"111100110",
30649=>"111010011",
30650=>"110110111",
30651=>"000000000",
30652=>"000111010",
30653=>"111010000",
30654=>"111100110",
30655=>"000000010",
30656=>"010001111",
30657=>"000000000",
30658=>"110111100",
30659=>"000001011",
30660=>"011010000",
30661=>"101111100",
30662=>"011111010",
30663=>"100000111",
30664=>"111100000",
30665=>"110000100",
30666=>"000010000",
30667=>"111000001",
30668=>"010000000",
30669=>"011111110",
30670=>"000000101",
30671=>"000000010",
30672=>"111111000",
30673=>"100111111",
30674=>"111011011",
30675=>"111111111",
30676=>"111111111",
30677=>"000011111",
30678=>"000100101",
30679=>"110010100",
30680=>"010000000",
30681=>"001110001",
30682=>"101110000",
30683=>"101100101",
30684=>"110110010",
30685=>"000111000",
30686=>"010010110",
30687=>"100000101",
30688=>"111101111",
30689=>"000001100",
30690=>"101010010",
30691=>"000101111",
30692=>"111111011",
30693=>"010000000",
30694=>"000000000",
30695=>"100000000",
30696=>"010110000",
30697=>"000000100",
30698=>"101011001",
30699=>"111111111",
30700=>"110000000",
30701=>"011110100",
30702=>"111001000",
30703=>"111001001",
30704=>"111111000",
30705=>"111111001",
30706=>"110111011",
30707=>"111111110",
30708=>"110001011",
30709=>"000100101",
30710=>"001001001",
30711=>"101111111",
30712=>"111110001",
30713=>"111111100",
30714=>"111111110",
30715=>"000111010",
30716=>"001001101",
30717=>"000101010",
30718=>"001011011",
30719=>"000101001",
30720=>"010111101",
30721=>"101111111",
30722=>"000101010",
30723=>"000000010",
30724=>"100111000",
30725=>"000111101",
30726=>"111011011",
30727=>"011011000",
30728=>"001000100",
30729=>"010010111",
30730=>"011110100",
30731=>"101011101",
30732=>"101101101",
30733=>"101101101",
30734=>"011011010",
30735=>"111111111",
30736=>"000000000",
30737=>"000000011",
30738=>"101101111",
30739=>"000011000",
30740=>"111111111",
30741=>"110100001",
30742=>"000001001",
30743=>"000000000",
30744=>"010000000",
30745=>"100101111",
30746=>"101101010",
30747=>"010010000",
30748=>"100000101",
30749=>"011110010",
30750=>"100111011",
30751=>"000000101",
30752=>"101100100",
30753=>"101100111",
30754=>"101010001",
30755=>"000000000",
30756=>"110100100",
30757=>"100111111",
30758=>"100101100",
30759=>"101010101",
30760=>"101101100",
30761=>"011011000",
30762=>"000000000",
30763=>"010000001",
30764=>"011011011",
30765=>"110010010",
30766=>"000101111",
30767=>"111111101",
30768=>"010101000",
30769=>"100011011",
30770=>"000000000",
30771=>"010111010",
30772=>"011111101",
30773=>"010111101",
30774=>"001001100",
30775=>"011111101",
30776=>"001101100",
30777=>"001000000",
30778=>"100100110",
30779=>"010010010",
30780=>"000001001",
30781=>"111111101",
30782=>"010000001",
30783=>"000100000",
30784=>"001001000",
30785=>"110110100",
30786=>"000110110",
30787=>"000010110",
30788=>"111001010",
30789=>"011101001",
30790=>"111010100",
30791=>"000000000",
30792=>"101100010",
30793=>"010101010",
30794=>"011101111",
30795=>"010011011",
30796=>"000100101",
30797=>"101001000",
30798=>"000100100",
30799=>"010010010",
30800=>"001000111",
30801=>"000000111",
30802=>"111010101",
30803=>"001001000",
30804=>"001001000",
30805=>"001011100",
30806=>"011000100",
30807=>"101100000",
30808=>"000111100",
30809=>"110011000",
30810=>"000000001",
30811=>"001111111",
30812=>"000000000",
30813=>"001001001",
30814=>"000100111",
30815=>"001110101",
30816=>"111111111",
30817=>"111000000",
30818=>"000100001",
30819=>"110000000",
30820=>"110111100",
30821=>"001110100",
30822=>"111010101",
30823=>"110110010",
30824=>"000010110",
30825=>"010110111",
30826=>"001010111",
30827=>"110110010",
30828=>"010010011",
30829=>"010110000",
30830=>"010010000",
30831=>"110101101",
30832=>"001001111",
30833=>"111111110",
30834=>"000000101",
30835=>"111100000",
30836=>"111111111",
30837=>"100101101",
30838=>"101000100",
30839=>"111101111",
30840=>"000100100",
30841=>"010000000",
30842=>"111110111",
30843=>"000000000",
30844=>"110111011",
30845=>"100100001",
30846=>"000000000",
30847=>"001000111",
30848=>"000000110",
30849=>"000101000",
30850=>"010011100",
30851=>"111111111",
30852=>"111111001",
30853=>"110010101",
30854=>"001110111",
30855=>"100001011",
30856=>"101101111",
30857=>"110111111",
30858=>"010010000",
30859=>"100000000",
30860=>"000001001",
30861=>"010110010",
30862=>"111001000",
30863=>"101101101",
30864=>"111101111",
30865=>"101111101",
30866=>"000001101",
30867=>"101100000",
30868=>"011011011",
30869=>"000010111",
30870=>"111100101",
30871=>"100100110",
30872=>"010010111",
30873=>"000111000",
30874=>"010010000",
30875=>"000000000",
30876=>"111111000",
30877=>"000001001",
30878=>"010000100",
30879=>"011101001",
30880=>"111011001",
30881=>"100000000",
30882=>"001000010",
30883=>"000000000",
30884=>"000010000",
30885=>"101101111",
30886=>"000001011",
30887=>"010010011",
30888=>"011000111",
30889=>"001001000",
30890=>"000101111",
30891=>"011001001",
30892=>"110011101",
30893=>"010000000",
30894=>"111111111",
30895=>"010011010",
30896=>"000000111",
30897=>"011111001",
30898=>"101101100",
30899=>"100110010",
30900=>"100101000",
30901=>"010011110",
30902=>"111100100",
30903=>"100101101",
30904=>"000100100",
30905=>"111110110",
30906=>"000000011",
30907=>"111111000",
30908=>"111111010",
30909=>"000000000",
30910=>"101001110",
30911=>"010101110",
30912=>"101001101",
30913=>"011010000",
30914=>"000110101",
30915=>"111011011",
30916=>"011001000",
30917=>"110100100",
30918=>"000001000",
30919=>"000000000",
30920=>"001101111",
30921=>"101101001",
30922=>"100111100",
30923=>"111110100",
30924=>"101000111",
30925=>"001011110",
30926=>"010001101",
30927=>"100111111",
30928=>"000000101",
30929=>"111011000",
30930=>"111110110",
30931=>"111110101",
30932=>"101111111",
30933=>"100000100",
30934=>"101100000",
30935=>"010110111",
30936=>"101011010",
30937=>"001011001",
30938=>"110000000",
30939=>"010000000",
30940=>"000001000",
30941=>"000100000",
30942=>"111111011",
30943=>"000000100",
30944=>"000100011",
30945=>"000001110",
30946=>"100000001",
30947=>"111111111",
30948=>"000100010",
30949=>"101011111",
30950=>"111110101",
30951=>"011111111",
30952=>"000010001",
30953=>"111000101",
30954=>"110111001",
30955=>"100000000",
30956=>"111101101",
30957=>"101000000",
30958=>"000000000",
30959=>"000011111",
30960=>"111111111",
30961=>"101001101",
30962=>"000010010",
30963=>"000000000",
30964=>"010001001",
30965=>"110011101",
30966=>"100000110",
30967=>"000000011",
30968=>"000000000",
30969=>"111010110",
30970=>"111111111",
30971=>"000000100",
30972=>"111111000",
30973=>"101011101",
30974=>"011011000",
30975=>"011110111",
30976=>"011001001",
30977=>"000000111",
30978=>"000000111",
30979=>"111100010",
30980=>"000000100",
30981=>"010000000",
30982=>"111011110",
30983=>"111111110",
30984=>"011100100",
30985=>"100001101",
30986=>"110111000",
30987=>"000000011",
30988=>"101001110",
30989=>"001110000",
30990=>"111001001",
30991=>"100000000",
30992=>"110110010",
30993=>"000101000",
30994=>"000000000",
30995=>"000000011",
30996=>"111111000",
30997=>"001001000",
30998=>"000001000",
30999=>"000000010",
31000=>"110010000",
31001=>"010111000",
31002=>"011000000",
31003=>"000111110",
31004=>"111110110",
31005=>"000000000",
31006=>"111001000",
31007=>"000101111",
31008=>"010110010",
31009=>"001001111",
31010=>"111001101",
31011=>"100000100",
31012=>"000101100",
31013=>"100011110",
31014=>"111111000",
31015=>"101110100",
31016=>"110110111",
31017=>"111111111",
31018=>"000010011",
31019=>"110001000",
31020=>"000000100",
31021=>"111111110",
31022=>"110000111",
31023=>"000001001",
31024=>"000000000",
31025=>"000011001",
31026=>"111100000",
31027=>"000001010",
31028=>"111111000",
31029=>"111111010",
31030=>"000000100",
31031=>"011000000",
31032=>"110001111",
31033=>"111001101",
31034=>"000000100",
31035=>"111111100",
31036=>"100111111",
31037=>"100111111",
31038=>"001000101",
31039=>"110110000",
31040=>"010011101",
31041=>"000001111",
31042=>"111111000",
31043=>"110110000",
31044=>"000000101",
31045=>"011001000",
31046=>"010000111",
31047=>"101101101",
31048=>"101111111",
31049=>"110110000",
31050=>"101100000",
31051=>"111110111",
31052=>"001000111",
31053=>"001111011",
31054=>"100101101",
31055=>"101101111",
31056=>"001000001",
31057=>"010000000",
31058=>"111110100",
31059=>"100001000",
31060=>"000000101",
31061=>"110000011",
31062=>"100101110",
31063=>"111111000",
31064=>"110100111",
31065=>"110100110",
31066=>"001000001",
31067=>"000001001",
31068=>"001011011",
31069=>"001001011",
31070=>"001101111",
31071=>"011010000",
31072=>"000001101",
31073=>"110110000",
31074=>"101000100",
31075=>"100010100",
31076=>"100000100",
31077=>"001000001",
31078=>"110110000",
31079=>"010111110",
31080=>"111101000",
31081=>"000111100",
31082=>"111000100",
31083=>"110001101",
31084=>"100110111",
31085=>"000110000",
31086=>"111000000",
31087=>"001101111",
31088=>"100110101",
31089=>"111001000",
31090=>"100000000",
31091=>"011000000",
31092=>"111111000",
31093=>"011000000",
31094=>"001000010",
31095=>"000010010",
31096=>"000100111",
31097=>"000100111",
31098=>"000001000",
31099=>"101000000",
31100=>"110010110",
31101=>"100101000",
31102=>"110110010",
31103=>"110110110",
31104=>"001000000",
31105=>"010000000",
31106=>"011110101",
31107=>"010011111",
31108=>"111010000",
31109=>"110000000",
31110=>"011100111",
31111=>"000000011",
31112=>"011011010",
31113=>"001101001",
31114=>"011111010",
31115=>"111000000",
31116=>"000000000",
31117=>"000000111",
31118=>"000000000",
31119=>"000000110",
31120=>"010011001",
31121=>"110000001",
31122=>"001001001",
31123=>"111011111",
31124=>"011100011",
31125=>"010000110",
31126=>"111000000",
31127=>"100100110",
31128=>"011100101",
31129=>"101111111",
31130=>"001001111",
31131=>"010110010",
31132=>"111101111",
31133=>"101111000",
31134=>"111100011",
31135=>"000000000",
31136=>"001101110",
31137=>"001000000",
31138=>"001101010",
31139=>"110111100",
31140=>"010000101",
31141=>"101100101",
31142=>"000000001",
31143=>"001000100",
31144=>"110000001",
31145=>"110111000",
31146=>"111111111",
31147=>"111000000",
31148=>"001000010",
31149=>"101100101",
31150=>"000000100",
31151=>"111111010",
31152=>"000000010",
31153=>"001001110",
31154=>"000111111",
31155=>"100000010",
31156=>"011111010",
31157=>"111111111",
31158=>"000000100",
31159=>"000000000",
31160=>"001111111",
31161=>"010101110",
31162=>"011010011",
31163=>"100010000",
31164=>"110110111",
31165=>"011010000",
31166=>"011011001",
31167=>"111111101",
31168=>"110010111",
31169=>"000000111",
31170=>"000111110",
31171=>"110111100",
31172=>"000111000",
31173=>"100100011",
31174=>"000000010",
31175=>"100000111",
31176=>"111001001",
31177=>"001000001",
31178=>"001001001",
31179=>"011111101",
31180=>"000010111",
31181=>"011000011",
31182=>"010000111",
31183=>"000100000",
31184=>"000000100",
31185=>"111111111",
31186=>"001001000",
31187=>"010100000",
31188=>"000001111",
31189=>"100101111",
31190=>"111000000",
31191=>"111000100",
31192=>"100100111",
31193=>"001110000",
31194=>"101100100",
31195=>"010010000",
31196=>"001100011",
31197=>"111101000",
31198=>"010101001",
31199=>"000000010",
31200=>"101000111",
31201=>"111000000",
31202=>"000000000",
31203=>"101100101",
31204=>"010010000",
31205=>"101101111",
31206=>"000101111",
31207=>"100000010",
31208=>"001000000",
31209=>"001110010",
31210=>"011111001",
31211=>"010110001",
31212=>"101001000",
31213=>"001111000",
31214=>"000000000",
31215=>"111101111",
31216=>"000010010",
31217=>"011010111",
31218=>"111111000",
31219=>"111101000",
31220=>"111101110",
31221=>"111000000",
31222=>"000000001",
31223=>"000000101",
31224=>"111000110",
31225=>"101000000",
31226=>"011111110",
31227=>"100101110",
31228=>"000000101",
31229=>"001111110",
31230=>"000000001",
31231=>"000011111",
31232=>"001101100",
31233=>"111000001",
31234=>"000110000",
31235=>"110101010",
31236=>"111110010",
31237=>"100001110",
31238=>"001001111",
31239=>"110100010",
31240=>"100101111",
31241=>"000001101",
31242=>"000000001",
31243=>"000101101",
31244=>"111110010",
31245=>"010011010",
31246=>"011011011",
31247=>"000001000",
31248=>"110110000",
31249=>"000100000",
31250=>"000110111",
31251=>"111111000",
31252=>"111010000",
31253=>"111111101",
31254=>"011100011",
31255=>"100110010",
31256=>"111111101",
31257=>"001000000",
31258=>"000000101",
31259=>"000001000",
31260=>"000001010",
31261=>"001101111",
31262=>"001101110",
31263=>"010000000",
31264=>"000101011",
31265=>"100111111",
31266=>"000001000",
31267=>"000000000",
31268=>"011011000",
31269=>"100100101",
31270=>"000000000",
31271=>"000001010",
31272=>"111111111",
31273=>"110110010",
31274=>"000000000",
31275=>"001000100",
31276=>"111011011",
31277=>"000100100",
31278=>"000001001",
31279=>"001011001",
31280=>"000101101",
31281=>"111111111",
31282=>"000001000",
31283=>"001001000",
31284=>"000000011",
31285=>"110000110",
31286=>"000000001",
31287=>"010111101",
31288=>"001000001",
31289=>"000110010",
31290=>"100100011",
31291=>"111111000",
31292=>"100110000",
31293=>"000001111",
31294=>"000000000",
31295=>"011001011",
31296=>"110111110",
31297=>"111001101",
31298=>"111011010",
31299=>"011001001",
31300=>"000000000",
31301=>"100010010",
31302=>"000001001",
31303=>"000101111",
31304=>"011100111",
31305=>"010011011",
31306=>"000000000",
31307=>"111000011",
31308=>"000000100",
31309=>"111111101",
31310=>"111111011",
31311=>"111111000",
31312=>"001010000",
31313=>"110110111",
31314=>"100111010",
31315=>"011110101",
31316=>"000010110",
31317=>"110100011",
31318=>"000100000",
31319=>"000000111",
31320=>"011101011",
31321=>"101100000",
31322=>"111000010",
31323=>"110110000",
31324=>"000101001",
31325=>"001001000",
31326=>"111111001",
31327=>"000000000",
31328=>"111111110",
31329=>"000000100",
31330=>"001111110",
31331=>"111010010",
31332=>"100110110",
31333=>"000000100",
31334=>"000001101",
31335=>"001101111",
31336=>"000001100",
31337=>"001000101",
31338=>"000000111",
31339=>"111111101",
31340=>"000001000",
31341=>"111110101",
31342=>"001100001",
31343=>"100010000",
31344=>"101011110",
31345=>"000001101",
31346=>"010000100",
31347=>"000010000",
31348=>"010000101",
31349=>"000101000",
31350=>"010110111",
31351=>"110110001",
31352=>"000000000",
31353=>"111110100",
31354=>"100001011",
31355=>"001101000",
31356=>"110110101",
31357=>"100100101",
31358=>"000000111",
31359=>"000010110",
31360=>"111000000",
31361=>"110110111",
31362=>"000101101",
31363=>"111111001",
31364=>"100111110",
31365=>"100010010",
31366=>"011001001",
31367=>"111110010",
31368=>"011011111",
31369=>"111001111",
31370=>"101100000",
31371=>"001011101",
31372=>"011001001",
31373=>"011001111",
31374=>"000000000",
31375=>"000001110",
31376=>"101011010",
31377=>"000001111",
31378=>"100011101",
31379=>"110111101",
31380=>"111111101",
31381=>"000000111",
31382=>"011010110",
31383=>"011011000",
31384=>"000000100",
31385=>"110000010",
31386=>"000000101",
31387=>"000000000",
31388=>"011000000",
31389=>"111111100",
31390=>"001111111",
31391=>"010010010",
31392=>"111010111",
31393=>"000000001",
31394=>"111111000",
31395=>"000000000",
31396=>"001011100",
31397=>"110110111",
31398=>"100111110",
31399=>"011000001",
31400=>"111000000",
31401=>"110110110",
31402=>"101101101",
31403=>"110110111",
31404=>"111111111",
31405=>"001001101",
31406=>"001011001",
31407=>"101111111",
31408=>"000000000",
31409=>"011011011",
31410=>"101101101",
31411=>"100000000",
31412=>"111110110",
31413=>"101111111",
31414=>"101110000",
31415=>"001001001",
31416=>"011011011",
31417=>"111110100",
31418=>"000000100",
31419=>"000001000",
31420=>"001001101",
31421=>"000010000",
31422=>"000000000",
31423=>"000001111",
31424=>"000001111",
31425=>"000100111",
31426=>"000010011",
31427=>"100100100",
31428=>"111011001",
31429=>"100111111",
31430=>"000111010",
31431=>"000000000",
31432=>"000000000",
31433=>"111010000",
31434=>"000111111",
31435=>"111110000",
31436=>"001000100",
31437=>"011011001",
31438=>"000110110",
31439=>"111111101",
31440=>"000000111",
31441=>"111110011",
31442=>"000110110",
31443=>"111111111",
31444=>"000111111",
31445=>"000000000",
31446=>"000001001",
31447=>"010101101",
31448=>"110111011",
31449=>"000101101",
31450=>"111110111",
31451=>"101001000",
31452=>"110111111",
31453=>"011001100",
31454=>"000101000",
31455=>"000001111",
31456=>"011010010",
31457=>"001001011",
31458=>"101111110",
31459=>"111100100",
31460=>"000010010",
31461=>"110011000",
31462=>"101100011",
31463=>"110100100",
31464=>"000101000",
31465=>"110111000",
31466=>"000000000",
31467=>"000001000",
31468=>"111110000",
31469=>"100111110",
31470=>"000000000",
31471=>"001001000",
31472=>"101101100",
31473=>"111100100",
31474=>"000101001",
31475=>"001001111",
31476=>"011101110",
31477=>"000000000",
31478=>"001000000",
31479=>"100101110",
31480=>"000000000",
31481=>"000000000",
31482=>"111111101",
31483=>"010111111",
31484=>"000101101",
31485=>"000000001",
31486=>"110110101",
31487=>"101111110",
31488=>"000000000",
31489=>"001101101",
31490=>"111111001",
31491=>"001000000",
31492=>"010010001",
31493=>"000111111",
31494=>"011110111",
31495=>"111000000",
31496=>"000000000",
31497=>"101000111",
31498=>"000100011",
31499=>"000000000",
31500=>"001001011",
31501=>"111101101",
31502=>"011011011",
31503=>"101111010",
31504=>"000000000",
31505=>"000000000",
31506=>"110110000",
31507=>"000000100",
31508=>"111111011",
31509=>"111111111",
31510=>"010111111",
31511=>"111111110",
31512=>"001110000",
31513=>"111001101",
31514=>"111011100",
31515=>"000111111",
31516=>"111111110",
31517=>"111111111",
31518=>"000001111",
31519=>"000010000",
31520=>"000000000",
31521=>"000001011",
31522=>"001111111",
31523=>"011001001",
31524=>"111100100",
31525=>"100001000",
31526=>"001000000",
31527=>"111110101",
31528=>"111111111",
31529=>"110110111",
31530=>"000000001",
31531=>"111111101",
31532=>"011110010",
31533=>"110000101",
31534=>"000000000",
31535=>"110011111",
31536=>"000000000",
31537=>"110000011",
31538=>"000001001",
31539=>"000010000",
31540=>"101010000",
31541=>"010111110",
31542=>"110111110",
31543=>"000001001",
31544=>"000000000",
31545=>"000000000",
31546=>"100000111",
31547=>"111111111",
31548=>"100011011",
31549=>"101101000",
31550=>"000000111",
31551=>"011111111",
31552=>"000000000",
31553=>"101000001",
31554=>"010010011",
31555=>"000000000",
31556=>"111101111",
31557=>"000110000",
31558=>"101000000",
31559=>"111111100",
31560=>"111101100",
31561=>"011111101",
31562=>"101010010",
31563=>"000000111",
31564=>"000000110",
31565=>"000000000",
31566=>"100000100",
31567=>"101000111",
31568=>"001000000",
31569=>"100010000",
31570=>"000000111",
31571=>"001001001",
31572=>"111111111",
31573=>"110101111",
31574=>"111111111",
31575=>"001000001",
31576=>"001010110",
31577=>"111111001",
31578=>"111111111",
31579=>"000001000",
31580=>"000000000",
31581=>"000001001",
31582=>"111000000",
31583=>"000000001",
31584=>"000001011",
31585=>"000000111",
31586=>"011011000",
31587=>"110111110",
31588=>"000000000",
31589=>"111001011",
31590=>"010000011",
31591=>"111111111",
31592=>"000010000",
31593=>"001000000",
31594=>"000010000",
31595=>"010010001",
31596=>"011111011",
31597=>"111110010",
31598=>"110111101",
31599=>"110101111",
31600=>"000000000",
31601=>"000000000",
31602=>"001111011",
31603=>"000000110",
31604=>"000110110",
31605=>"111000001",
31606=>"000000000",
31607=>"110111101",
31608=>"111111001",
31609=>"000001100",
31610=>"000000000",
31611=>"111111000",
31612=>"000000000",
31613=>"100100000",
31614=>"111111110",
31615=>"001000000",
31616=>"111010111",
31617=>"001000000",
31618=>"111111000",
31619=>"111100111",
31620=>"011001000",
31621=>"111111111",
31622=>"111101011",
31623=>"011011111",
31624=>"000000000",
31625=>"111001111",
31626=>"000000000",
31627=>"000101101",
31628=>"111101110",
31629=>"101111111",
31630=>"000000010",
31631=>"000000001",
31632=>"110011000",
31633=>"000111001",
31634=>"111011000",
31635=>"000001001",
31636=>"000010010",
31637=>"000000011",
31638=>"010000000",
31639=>"000000000",
31640=>"000111001",
31641=>"111111101",
31642=>"110110000",
31643=>"000110010",
31644=>"000000000",
31645=>"000000101",
31646=>"000000000",
31647=>"000000000",
31648=>"111111011",
31649=>"100111111",
31650=>"111000000",
31651=>"011111111",
31652=>"000000111",
31653=>"111101000",
31654=>"000000000",
31655=>"000000011",
31656=>"111100110",
31657=>"000001000",
31658=>"000001000",
31659=>"000000000",
31660=>"110100101",
31661=>"000000000",
31662=>"000110000",
31663=>"111111111",
31664=>"001101111",
31665=>"010000100",
31666=>"110110110",
31667=>"100100111",
31668=>"111111111",
31669=>"010110111",
31670=>"111100101",
31671=>"000000110",
31672=>"001110110",
31673=>"010100000",
31674=>"001111111",
31675=>"000001001",
31676=>"111111111",
31677=>"111010000",
31678=>"000110111",
31679=>"000000101",
31680=>"111111100",
31681=>"111111111",
31682=>"110111111",
31683=>"000001111",
31684=>"111000000",
31685=>"001010111",
31686=>"000000100",
31687=>"111111100",
31688=>"111000000",
31689=>"111001000",
31690=>"000100011",
31691=>"001000000",
31692=>"000010011",
31693=>"000100100",
31694=>"111111111",
31695=>"101111111",
31696=>"010110110",
31697=>"011011000",
31698=>"000001000",
31699=>"010010000",
31700=>"000000000",
31701=>"000000011",
31702=>"000010000",
31703=>"000000100",
31704=>"111101111",
31705=>"000000000",
31706=>"111111111",
31707=>"111000000",
31708=>"000000010",
31709=>"000000001",
31710=>"111000101",
31711=>"100000000",
31712=>"111111111",
31713=>"000000000",
31714=>"110111110",
31715=>"010100110",
31716=>"000000000",
31717=>"000100111",
31718=>"000000000",
31719=>"010111111",
31720=>"000010000",
31721=>"001100110",
31722=>"000000101",
31723=>"001111000",
31724=>"000000001",
31725=>"000000111",
31726=>"000000000",
31727=>"000000111",
31728=>"111111111",
31729=>"100111111",
31730=>"000000000",
31731=>"001011000",
31732=>"101100111",
31733=>"111111111",
31734=>"000011001",
31735=>"111111111",
31736=>"000000111",
31737=>"101111111",
31738=>"100100000",
31739=>"000100001",
31740=>"111111111",
31741=>"111101001",
31742=>"010010000",
31743=>"111110110",
31744=>"010110010",
31745=>"001001001",
31746=>"110110110",
31747=>"000011111",
31748=>"101111111",
31749=>"000000110",
31750=>"000101001",
31751=>"001001001",
31752=>"000001001",
31753=>"000000111",
31754=>"110110100",
31755=>"001000011",
31756=>"110110111",
31757=>"010000010",
31758=>"100101000",
31759=>"110111111",
31760=>"010001011",
31761=>"110000111",
31762=>"000110000",
31763=>"000001001",
31764=>"011011011",
31765=>"001100100",
31766=>"001000000",
31767=>"110110100",
31768=>"110110010",
31769=>"010110110",
31770=>"000000010",
31771=>"000001011",
31772=>"010011110",
31773=>"100000000",
31774=>"001111111",
31775=>"001000000",
31776=>"110110110",
31777=>"001001000",
31778=>"101010000",
31779=>"000010000",
31780=>"000001001",
31781=>"100010010",
31782=>"011110110",
31783=>"011011011",
31784=>"111111101",
31785=>"000000110",
31786=>"011000011",
31787=>"010111011",
31788=>"001010010",
31789=>"111001100",
31790=>"010000001",
31791=>"011011011",
31792=>"011001000",
31793=>"100100101",
31794=>"101000000",
31795=>"111111010",
31796=>"111000001",
31797=>"011000010",
31798=>"111111001",
31799=>"011011011",
31800=>"001011001",
31801=>"011001000",
31802=>"001111000",
31803=>"011011010",
31804=>"000011001",
31805=>"111011101",
31806=>"100100011",
31807=>"000001001",
31808=>"111110110",
31809=>"010011111",
31810=>"110100000",
31811=>"010110100",
31812=>"000100111",
31813=>"001111110",
31814=>"011000001",
31815=>"100100100",
31816=>"011111111",
31817=>"001001001",
31818=>"011010111",
31819=>"001011000",
31820=>"110100000",
31821=>"011011010",
31822=>"010010110",
31823=>"111011010",
31824=>"011000000",
31825=>"001110000",
31826=>"001001000",
31827=>"001000000",
31828=>"001000111",
31829=>"110010011",
31830=>"101111011",
31831=>"100100110",
31832=>"100100110",
31833=>"000000000",
31834=>"000011001",
31835=>"001000000",
31836=>"000001011",
31837=>"000100000",
31838=>"101101100",
31839=>"110100110",
31840=>"111100110",
31841=>"111111010",
31842=>"100110110",
31843=>"001011011",
31844=>"011011001",
31845=>"011001001",
31846=>"000001001",
31847=>"011001001",
31848=>"001001011",
31849=>"101100111",
31850=>"111111000",
31851=>"100111100",
31852=>"110111000",
31853=>"100110100",
31854=>"011100001",
31855=>"011001011",
31856=>"011111000",
31857=>"011000011",
31858=>"011001111",
31859=>"100110110",
31860=>"111010010",
31861=>"000110001",
31862=>"011000000",
31863=>"001101000",
31864=>"001111011",
31865=>"001001001",
31866=>"111001000",
31867=>"100100110",
31868=>"111011100",
31869=>"000000001",
31870=>"110101001",
31871=>"001000100",
31872=>"011110100",
31873=>"111110110",
31874=>"001001001",
31875=>"000111011",
31876=>"011011011",
31877=>"011011111",
31878=>"011001011",
31879=>"000000000",
31880=>"000000000",
31881=>"000011000",
31882=>"000001011",
31883=>"100000010",
31884=>"111110100",
31885=>"011001100",
31886=>"000001001",
31887=>"010000011",
31888=>"010010010",
31889=>"010111011",
31890=>"011000000",
31891=>"010000010",
31892=>"000001001",
31893=>"110110110",
31894=>"000001000",
31895=>"001111011",
31896=>"111011000",
31897=>"101001001",
31898=>"100100111",
31899=>"111111111",
31900=>"001001001",
31901=>"000000111",
31902=>"001001001",
31903=>"110110111",
31904=>"010000000",
31905=>"111000111",
31906=>"111111110",
31907=>"000010010",
31908=>"111011001",
31909=>"111111100",
31910=>"010000011",
31911=>"011001000",
31912=>"110000010",
31913=>"000001000",
31914=>"111110111",
31915=>"100110110",
31916=>"111000000",
31917=>"000001001",
31918=>"001001011",
31919=>"001101101",
31920=>"111011001",
31921=>"111111000",
31922=>"111100100",
31923=>"110001100",
31924=>"100000101",
31925=>"101001001",
31926=>"000010010",
31927=>"001010011",
31928=>"001001000",
31929=>"000011010",
31930=>"010011001",
31931=>"100100001",
31932=>"001001000",
31933=>"110110110",
31934=>"000000000",
31935=>"001110111",
31936=>"010011001",
31937=>"000000001",
31938=>"111100000",
31939=>"100101001",
31940=>"001000000",
31941=>"111011111",
31942=>"000010011",
31943=>"100110010",
31944=>"010001000",
31945=>"100100110",
31946=>"100100000",
31947=>"000101101",
31948=>"001001011",
31949=>"001001001",
31950=>"001000001",
31951=>"111110100",
31952=>"111110110",
31953=>"100001101",
31954=>"010001011",
31955=>"100000011",
31956=>"111111011",
31957=>"111010111",
31958=>"101100110",
31959=>"000001011",
31960=>"011011001",
31961=>"000011001",
31962=>"111111111",
31963=>"110110110",
31964=>"111111011",
31965=>"111110110",
31966=>"001001000",
31967=>"011001001",
31968=>"100100111",
31969=>"111110110",
31970=>"100101100",
31971=>"000000000",
31972=>"000001000",
31973=>"100100100",
31974=>"001000100",
31975=>"101111001",
31976=>"100101111",
31977=>"100110110",
31978=>"110100100",
31979=>"110100000",
31980=>"100100110",
31981=>"001000011",
31982=>"000110010",
31983=>"001011011",
31984=>"000110010",
31985=>"010000111",
31986=>"000011011",
31987=>"011011111",
31988=>"000000011",
31989=>"000101000",
31990=>"100100011",
31991=>"000001011",
31992=>"011110111",
31993=>"001001011",
31994=>"110110110",
31995=>"011110100",
31996=>"011011111",
31997=>"100001101",
31998=>"001001000",
31999=>"001101001",
32000=>"011001000",
32001=>"000000111",
32002=>"000000000",
32003=>"000110111",
32004=>"000000100",
32005=>"000011010",
32006=>"001001101",
32007=>"101000110",
32008=>"000001011",
32009=>"000001111",
32010=>"010100110",
32011=>"110101101",
32012=>"011011100",
32013=>"110001000",
32014=>"101001001",
32015=>"000000011",
32016=>"110111000",
32017=>"110000000",
32018=>"001000010",
32019=>"101111111",
32020=>"001111010",
32021=>"111111111",
32022=>"011100001",
32023=>"111111010",
32024=>"000100100",
32025=>"101000000",
32026=>"000000000",
32027=>"011010100",
32028=>"000100111",
32029=>"000111111",
32030=>"111000000",
32031=>"001111111",
32032=>"110111000",
32033=>"000100000",
32034=>"111000101",
32035=>"110110111",
32036=>"110111111",
32037=>"110100000",
32038=>"010111010",
32039=>"010000001",
32040=>"111111000",
32041=>"111111000",
32042=>"101001000",
32043=>"101000101",
32044=>"110100111",
32045=>"000000110",
32046=>"000111110",
32047=>"001001011",
32048=>"101101011",
32049=>"001101001",
32050=>"000110111",
32051=>"101000001",
32052=>"001000101",
32053=>"000101110",
32054=>"110111111",
32055=>"000000111",
32056=>"110010101",
32057=>"001110100",
32058=>"100100100",
32059=>"111101111",
32060=>"000010000",
32061=>"111111000",
32062=>"011000001",
32063=>"011111111",
32064=>"100000000",
32065=>"100000000",
32066=>"101111111",
32067=>"101110100",
32068=>"100100010",
32069=>"011000010",
32070=>"001000110",
32071=>"100111100",
32072=>"000000011",
32073=>"110111010",
32074=>"000000000",
32075=>"001000001",
32076=>"001000111",
32077=>"011111010",
32078=>"101101110",
32079=>"000000111",
32080=>"111111000",
32081=>"001011000",
32082=>"011111010",
32083=>"011000100",
32084=>"101101000",
32085=>"001000011",
32086=>"011001001",
32087=>"111110010",
32088=>"110100100",
32089=>"111111111",
32090=>"100101001",
32091=>"111011110",
32092=>"000000000",
32093=>"001001001",
32094=>"111111110",
32095=>"110011011",
32096=>"000000000",
32097=>"011010010",
32098=>"010000000",
32099=>"100111001",
32100=>"110111000",
32101=>"010011011",
32102=>"000001111",
32103=>"000101111",
32104=>"000010001",
32105=>"000110010",
32106=>"010000111",
32107=>"010000000",
32108=>"000000000",
32109=>"000000000",
32110=>"001001010",
32111=>"000001010",
32112=>"100100101",
32113=>"010000101",
32114=>"000111111",
32115=>"101000101",
32116=>"010010111",
32117=>"000000000",
32118=>"000110111",
32119=>"111111111",
32120=>"000000010",
32121=>"111001000",
32122=>"000000110",
32123=>"110111000",
32124=>"000110111",
32125=>"110100100",
32126=>"010101101",
32127=>"111111001",
32128=>"100000111",
32129=>"111000000",
32130=>"111000010",
32131=>"001010010",
32132=>"011010010",
32133=>"111101001",
32134=>"000011000",
32135=>"011000000",
32136=>"101101011",
32137=>"111000000",
32138=>"000010110",
32139=>"110000111",
32140=>"001000000",
32141=>"101111011",
32142=>"011111010",
32143=>"101001101",
32144=>"100111110",
32145=>"010000000",
32146=>"101000101",
32147=>"111000000",
32148=>"111111001",
32149=>"110110000",
32150=>"010111101",
32151=>"111011011",
32152=>"000000111",
32153=>"000000010",
32154=>"000001101",
32155=>"111111111",
32156=>"111011010",
32157=>"100111010",
32158=>"000010111",
32159=>"001000101",
32160=>"100110110",
32161=>"111010100",
32162=>"110111000",
32163=>"011100101",
32164=>"111000000",
32165=>"111001011",
32166=>"111110110",
32167=>"010000111",
32168=>"010100000",
32169=>"101000110",
32170=>"110111111",
32171=>"000000000",
32172=>"001000000",
32173=>"111110000",
32174=>"110101110",
32175=>"010111110",
32176=>"000000000",
32177=>"110000000",
32178=>"111000000",
32179=>"000100110",
32180=>"011011111",
32181=>"101100010",
32182=>"010000000",
32183=>"011010000",
32184=>"000010010",
32185=>"110110100",
32186=>"111101000",
32187=>"110011111",
32188=>"000000000",
32189=>"100110000",
32190=>"110110110",
32191=>"000110100",
32192=>"000010010",
32193=>"000000001",
32194=>"110110100",
32195=>"100110110",
32196=>"101000000",
32197=>"001001011",
32198=>"000100000",
32199=>"101000000",
32200=>"011110001",
32201=>"101000001",
32202=>"000000100",
32203=>"000111000",
32204=>"000000000",
32205=>"000011011",
32206=>"011101111",
32207=>"111110000",
32208=>"010010010",
32209=>"110110110",
32210=>"111111101",
32211=>"000000111",
32212=>"011000001",
32213=>"000000110",
32214=>"000110011",
32215=>"000111111",
32216=>"000000111",
32217=>"011111111",
32218=>"011001000",
32219=>"100000000",
32220=>"000001100",
32221=>"001000011",
32222=>"000000000",
32223=>"110100000",
32224=>"001001111",
32225=>"000000001",
32226=>"110111010",
32227=>"110010000",
32228=>"101000001",
32229=>"000000111",
32230=>"000000100",
32231=>"010011001",
32232=>"000001100",
32233=>"000000000",
32234=>"100001001",
32235=>"111001001",
32236=>"010010010",
32237=>"111000000",
32238=>"000000000",
32239=>"001000000",
32240=>"111111111",
32241=>"100100000",
32242=>"011101100",
32243=>"001001110",
32244=>"110000001",
32245=>"000111000",
32246=>"110000000",
32247=>"101101111",
32248=>"011000111",
32249=>"010000110",
32250=>"000010010",
32251=>"000000010",
32252=>"011111010",
32253=>"100111110",
32254=>"110111111",
32255=>"111000000",
32256=>"000000110",
32257=>"111000010",
32258=>"000100110",
32259=>"111000100",
32260=>"111011011",
32261=>"000010011",
32262=>"000000111",
32263=>"110111011",
32264=>"000101001",
32265=>"101000000",
32266=>"100001000",
32267=>"101001011",
32268=>"000110111",
32269=>"011001111",
32270=>"100011001",
32271=>"000000000",
32272=>"100010110",
32273=>"001000000",
32274=>"000111000",
32275=>"111111001",
32276=>"000100011",
32277=>"111111010",
32278=>"100111001",
32279=>"010010010",
32280=>"111001101",
32281=>"111111111",
32282=>"000101111",
32283=>"101101101",
32284=>"101101101",
32285=>"000000000",
32286=>"000000000",
32287=>"000000000",
32288=>"110111000",
32289=>"101101111",
32290=>"000010000",
32291=>"001011010",
32292=>"001101111",
32293=>"101101110",
32294=>"011001000",
32295=>"110000001",
32296=>"101101011",
32297=>"110011000",
32298=>"000000000",
32299=>"111111101",
32300=>"001111110",
32301=>"000000110",
32302=>"000111111",
32303=>"111101010",
32304=>"000111010",
32305=>"001100101",
32306=>"000010100",
32307=>"000000010",
32308=>"000000000",
32309=>"111111110",
32310=>"100000000",
32311=>"011110000",
32312=>"000011101",
32313=>"000000101",
32314=>"111010000",
32315=>"000001011",
32316=>"110110111",
32317=>"000111011",
32318=>"100000101",
32319=>"100000111",
32320=>"000000000",
32321=>"111101111",
32322=>"111101111",
32323=>"101000000",
32324=>"000000011",
32325=>"000010000",
32326=>"000000001",
32327=>"001000101",
32328=>"000100111",
32329=>"000101111",
32330=>"010111101",
32331=>"010011000",
32332=>"000001101",
32333=>"110100110",
32334=>"101001011",
32335=>"111110111",
32336=>"001000000",
32337=>"011111111",
32338=>"100101001",
32339=>"001111111",
32340=>"101000000",
32341=>"001111110",
32342=>"000011011",
32343=>"111000010",
32344=>"000001000",
32345=>"000100100",
32346=>"111110000",
32347=>"111101001",
32348=>"000000101",
32349=>"000000000",
32350=>"000001010",
32351=>"000011001",
32352=>"111101101",
32353=>"000000111",
32354=>"101101101",
32355=>"111000000",
32356=>"000100000",
32357=>"101100110",
32358=>"010010000",
32359=>"111101000",
32360=>"111000001",
32361=>"000000100",
32362=>"000100101",
32363=>"000001111",
32364=>"110111011",
32365=>"001100110",
32366=>"000100010",
32367=>"011010001",
32368=>"001001111",
32369=>"000000100",
32370=>"001000001",
32371=>"110010000",
32372=>"001000000",
32373=>"000000001",
32374=>"010101101",
32375=>"001110111",
32376=>"111000000",
32377=>"000111111",
32378=>"000000000",
32379=>"000000001",
32380=>"001110100",
32381=>"000001111",
32382=>"000000011",
32383=>"100110111",
32384=>"111000010",
32385=>"000111111",
32386=>"001111111",
32387=>"111000001",
32388=>"000000100",
32389=>"111001111",
32390=>"101101011",
32391=>"111100011",
32392=>"100100110",
32393=>"000101000",
32394=>"111011011",
32395=>"000001111",
32396=>"000000000",
32397=>"111010000",
32398=>"000100100",
32399=>"001000000",
32400=>"100111010",
32401=>"111101000",
32402=>"000000101",
32403=>"000000000",
32404=>"110100100",
32405=>"000000111",
32406=>"000010110",
32407=>"010011000",
32408=>"111111001",
32409=>"111101000",
32410=>"100000100",
32411=>"111000000",
32412=>"000111011",
32413=>"111100000",
32414=>"100101011",
32415=>"010111101",
32416=>"101111111",
32417=>"010100000",
32418=>"000111111",
32419=>"111101101",
32420=>"111011000",
32421=>"101111111",
32422=>"111110100",
32423=>"111001011",
32424=>"111000011",
32425=>"000000100",
32426=>"111100010",
32427=>"000000000",
32428=>"011010000",
32429=>"101101101",
32430=>"100001001",
32431=>"000111111",
32432=>"110100000",
32433=>"111111110",
32434=>"101111111",
32435=>"001001000",
32436=>"001011001",
32437=>"010010000",
32438=>"111111111",
32439=>"101001100",
32440=>"111111111",
32441=>"111011110",
32442=>"111110011",
32443=>"010000010",
32444=>"101101111",
32445=>"111111010",
32446=>"000001011",
32447=>"110100000",
32448=>"000000100",
32449=>"000000101",
32450=>"101101111",
32451=>"100100110",
32452=>"000111110",
32453=>"100100001",
32454=>"000000011",
32455=>"000010101",
32456=>"000000111",
32457=>"110011010",
32458=>"111111111",
32459=>"111111010",
32460=>"111111000",
32461=>"100101001",
32462=>"100010000",
32463=>"111101001",
32464=>"100110100",
32465=>"111111010",
32466=>"011000101",
32467=>"000111111",
32468=>"000000000",
32469=>"110110110",
32470=>"000000101",
32471=>"101111000",
32472=>"010000000",
32473=>"000000101",
32474=>"101110111",
32475=>"010000000",
32476=>"100100001",
32477=>"111111010",
32478=>"111101001",
32479=>"000000111",
32480=>"111000011",
32481=>"101101101",
32482=>"101001000",
32483=>"001001110",
32484=>"010111111",
32485=>"000110010",
32486=>"000000000",
32487=>"010111000",
32488=>"000100100",
32489=>"010111101",
32490=>"000000000",
32491=>"000010111",
32492=>"100111111",
32493=>"111101111",
32494=>"000000001",
32495=>"000110000",
32496=>"000110000",
32497=>"000000100",
32498=>"110011001",
32499=>"100000010",
32500=>"000011000",
32501=>"101101000",
32502=>"010000100",
32503=>"111101000",
32504=>"001101110",
32505=>"111000000",
32506=>"111101111",
32507=>"000110101",
32508=>"000100111",
32509=>"101101010",
32510=>"011011011",
32511=>"110111111",
32512=>"000001001",
32513=>"111000000",
32514=>"001000001",
32515=>"000000001",
32516=>"110111111",
32517=>"111111110",
32518=>"000010011",
32519=>"110101000",
32520=>"111111111",
32521=>"101001000",
32522=>"110110010",
32523=>"101010110",
32524=>"000000000",
32525=>"000000101",
32526=>"100111111",
32527=>"100000000",
32528=>"111100000",
32529=>"000111111",
32530=>"000100101",
32531=>"111001100",
32532=>"111111000",
32533=>"101001111",
32534=>"000010000",
32535=>"110111111",
32536=>"101000111",
32537=>"111110001",
32538=>"101101111",
32539=>"000000000",
32540=>"110101000",
32541=>"110000001",
32542=>"001101110",
32543=>"010010000",
32544=>"010110000",
32545=>"000010000",
32546=>"010010111",
32547=>"111111111",
32548=>"011111110",
32549=>"001011001",
32550=>"100001000",
32551=>"001111011",
32552=>"000010000",
32553=>"000001001",
32554=>"111000010",
32555=>"111111110",
32556=>"111110111",
32557=>"111110001",
32558=>"010110010",
32559=>"010010010",
32560=>"011010111",
32561=>"111111100",
32562=>"000000000",
32563=>"010011000",
32564=>"110111101",
32565=>"001100011",
32566=>"111111000",
32567=>"000000000",
32568=>"111111111",
32569=>"000001111",
32570=>"010000101",
32571=>"011111111",
32572=>"110111011",
32573=>"110111111",
32574=>"001000101",
32575=>"000111111",
32576=>"000101001",
32577=>"101001111",
32578=>"000101000",
32579=>"100111011",
32580=>"001000101",
32581=>"000101101",
32582=>"110101111",
32583=>"000000100",
32584=>"000001111",
32585=>"011110111",
32586=>"001101111",
32587=>"101000000",
32588=>"000000000",
32589=>"010101001",
32590=>"001111111",
32591=>"010000000",
32592=>"101100101",
32593=>"010111111",
32594=>"010011111",
32595=>"011001000",
32596=>"101000000",
32597=>"111000000",
32598=>"110111011",
32599=>"101110101",
32600=>"101001101",
32601=>"001001000",
32602=>"111111101",
32603=>"111111011",
32604=>"000000001",
32605=>"000000111",
32606=>"000000000",
32607=>"011111100",
32608=>"101101111",
32609=>"000010110",
32610=>"000000000",
32611=>"110111100",
32612=>"000110010",
32613=>"000000011",
32614=>"110111111",
32615=>"111111000",
32616=>"010010111",
32617=>"000010111",
32618=>"000100000",
32619=>"110110111",
32620=>"000110111",
32621=>"010111010",
32622=>"000000111",
32623=>"000011111",
32624=>"010110010",
32625=>"001000111",
32626=>"111111001",
32627=>"100111000",
32628=>"111011010",
32629=>"000000000",
32630=>"101101111",
32631=>"000000111",
32632=>"001001000",
32633=>"000001111",
32634=>"111111111",
32635=>"111000111",
32636=>"011011111",
32637=>"010100000",
32638=>"001010010",
32639=>"111010101",
32640=>"110101010",
32641=>"111100110",
32642=>"111110000",
32643=>"001000111",
32644=>"000000000",
32645=>"011111111",
32646=>"101110100",
32647=>"000110111",
32648=>"011111101",
32649=>"010111001",
32650=>"000000000",
32651=>"000111001",
32652=>"000110111",
32653=>"010110110",
32654=>"101100100",
32655=>"000001011",
32656=>"111001101",
32657=>"011010110",
32658=>"011111010",
32659=>"100100111",
32660=>"111111010",
32661=>"111110001",
32662=>"000000000",
32663=>"110110110",
32664=>"111001111",
32665=>"001000001",
32666=>"111010000",
32667=>"111111000",
32668=>"110101001",
32669=>"100110101",
32670=>"110000010",
32671=>"101000101",
32672=>"101100010",
32673=>"000000110",
32674=>"101000101",
32675=>"000000001",
32676=>"000000000",
32677=>"110111111",
32678=>"011011011",
32679=>"000000101",
32680=>"111111011",
32681=>"000100111",
32682=>"101000100",
32683=>"111000000",
32684=>"101010000",
32685=>"000101111",
32686=>"000000100",
32687=>"000000000",
32688=>"000101101",
32689=>"000011111",
32690=>"000100000",
32691=>"100111111",
32692=>"110110111",
32693=>"000000000",
32694=>"111111101",
32695=>"000101000",
32696=>"110110110",
32697=>"110011011",
32698=>"011010100",
32699=>"000110111",
32700=>"010111111",
32701=>"111111100",
32702=>"000101111",
32703=>"001000111",
32704=>"000011110",
32705=>"001000111",
32706=>"001111110",
32707=>"000010010",
32708=>"010111111",
32709=>"011000000",
32710=>"111111111",
32711=>"001000000",
32712=>"111101111",
32713=>"100001000",
32714=>"111111011",
32715=>"001101111",
32716=>"000010000",
32717=>"010111101",
32718=>"111111111",
32719=>"111110100",
32720=>"010000000",
32721=>"111011011",
32722=>"110011011",
32723=>"001001000",
32724=>"111110000",
32725=>"000001011",
32726=>"100000001",
32727=>"111111110",
32728=>"001111011",
32729=>"000111000",
32730=>"100000000",
32731=>"000000110",
32732=>"000000000",
32733=>"101101111",
32734=>"111111011",
32735=>"001000111",
32736=>"000000000",
32737=>"100001101",
32738=>"000010000",
32739=>"101101111",
32740=>"011111011",
32741=>"000111011",
32742=>"010111111",
32743=>"000000000",
32744=>"000011111",
32745=>"111110000",
32746=>"001011011",
32747=>"001111111",
32748=>"101100101",
32749=>"101100101",
32750=>"000010010",
32751=>"111010110",
32752=>"111111111",
32753=>"111001000",
32754=>"000010010",
32755=>"110100000",
32756=>"010010110",
32757=>"111011111",
32758=>"110000011",
32759=>"111111111",
32760=>"101100011",
32761=>"010010000",
32762=>"011111111",
32763=>"010011101",
32764=>"000000000",
32765=>"110111100",
32766=>"001000001",
32767=>"010101000",
32768=>"010010101",
32769=>"010111011",
32770=>"111000001",
32771=>"111111001",
32772=>"001001001",
32773=>"111110001",
32774=>"000010000",
32775=>"000111111",
32776=>"000000110",
32777=>"000100100",
32778=>"101101111",
32779=>"101000001",
32780=>"000100100",
32781=>"010000000",
32782=>"111111101",
32783=>"110110001",
32784=>"100110110",
32785=>"110000000",
32786=>"000000000",
32787=>"101101101",
32788=>"111100000",
32789=>"000000000",
32790=>"110111011",
32791=>"110010000",
32792=>"000000000",
32793=>"010100000",
32794=>"110111111",
32795=>"111111010",
32796=>"000000000",
32797=>"000010000",
32798=>"111111111",
32799=>"000000000",
32800=>"100001000",
32801=>"111111101",
32802=>"000000001",
32803=>"010011111",
32804=>"001011001",
32805=>"100111001",
32806=>"010111110",
32807=>"111101111",
32808=>"101111101",
32809=>"000111111",
32810=>"111111110",
32811=>"000000000",
32812=>"111111110",
32813=>"001000000",
32814=>"010010111",
32815=>"011001101",
32816=>"111011111",
32817=>"100100100",
32818=>"000110110",
32819=>"110110111",
32820=>"111111011",
32821=>"000000000",
32822=>"000111101",
32823=>"111111010",
32824=>"111000000",
32825=>"000000010",
32826=>"000001000",
32827=>"111101100",
32828=>"010000001",
32829=>"101111111",
32830=>"001000001",
32831=>"100111000",
32832=>"111000110",
32833=>"110101111",
32834=>"011111111",
32835=>"011011110",
32836=>"000000110",
32837=>"000000010",
32838=>"101000001",
32839=>"111000000",
32840=>"000001000",
32841=>"101001000",
32842=>"000000000",
32843=>"111111110",
32844=>"111000000",
32845=>"000000100",
32846=>"001000000",
32847=>"111000000",
32848=>"110110000",
32849=>"000111111",
32850=>"000001100",
32851=>"000000000",
32852=>"010010000",
32853=>"100111100",
32854=>"011001100",
32855=>"000001000",
32856=>"000000001",
32857=>"010100100",
32858=>"111111001",
32859=>"100100100",
32860=>"010110110",
32861=>"111001001",
32862=>"111000000",
32863=>"110100111",
32864=>"010110110",
32865=>"110000000",
32866=>"000001000",
32867=>"110110000",
32868=>"101101110",
32869=>"000000001",
32870=>"101101111",
32871=>"111111000",
32872=>"111110111",
32873=>"000000111",
32874=>"111111010",
32875=>"010100110",
32876=>"010111111",
32877=>"111111111",
32878=>"111000101",
32879=>"111111011",
32880=>"001001001",
32881=>"111001111",
32882=>"000111111",
32883=>"001001000",
32884=>"010111000",
32885=>"000000111",
32886=>"111111101",
32887=>"010000000",
32888=>"111101001",
32889=>"110000000",
32890=>"001111101",
32891=>"000000101",
32892=>"101001100",
32893=>"000100010",
32894=>"101000000",
32895=>"011110110",
32896=>"000000000",
32897=>"000000000",
32898=>"100000111",
32899=>"111111000",
32900=>"000110110",
32901=>"000000110",
32902=>"011111000",
32903=>"000001000",
32904=>"100100100",
32905=>"000000101",
32906=>"111101111",
32907=>"010111111",
32908=>"111000000",
32909=>"000000000",
32910=>"011011000",
32911=>"110011100",
32912=>"010111011",
32913=>"100110110",
32914=>"110010010",
32915=>"110010111",
32916=>"010010111",
32917=>"101001000",
32918=>"110111111",
32919=>"111010011",
32920=>"111111111",
32921=>"110010001",
32922=>"101101011",
32923=>"001001100",
32924=>"111010000",
32925=>"000001000",
32926=>"111111011",
32927=>"100111110",
32928=>"110100010",
32929=>"111000010",
32930=>"010110111",
32931=>"110001001",
32932=>"100001111",
32933=>"000000000",
32934=>"010111000",
32935=>"111111111",
32936=>"110000100",
32937=>"111111111",
32938=>"001000101",
32939=>"111010001",
32940=>"111100000",
32941=>"110111000",
32942=>"000000011",
32943=>"111001000",
32944=>"111111111",
32945=>"100110101",
32946=>"011010000",
32947=>"011001100",
32948=>"110010000",
32949=>"111101111",
32950=>"000000000",
32951=>"011111111",
32952=>"001000000",
32953=>"100110100",
32954=>"111000000",
32955=>"111011000",
32956=>"011000110",
32957=>"000110111",
32958=>"110110010",
32959=>"000000000",
32960=>"000000000",
32961=>"111001010",
32962=>"111010111",
32963=>"100101110",
32964=>"000000010",
32965=>"011010001",
32966=>"000000000",
32967=>"101000000",
32968=>"000000000",
32969=>"000000000",
32970=>"000000001",
32971=>"100001101",
32972=>"111111110",
32973=>"011000000",
32974=>"110110001",
32975=>"000000000",
32976=>"010000000",
32977=>"110110010",
32978=>"010000000",
32979=>"000000000",
32980=>"011001000",
32981=>"111110000",
32982=>"111110100",
32983=>"000000101",
32984=>"000000000",
32985=>"001000100",
32986=>"011001010",
32987=>"111111000",
32988=>"010101000",
32989=>"000000000",
32990=>"000000000",
32991=>"111111000",
32992=>"111000000",
32993=>"000000000",
32994=>"000001000",
32995=>"011001001",
32996=>"101101000",
32997=>"000010000",
32998=>"000010010",
32999=>"000100010",
33000=>"000111111",
33001=>"110010001",
33002=>"001011100",
33003=>"011000101",
33004=>"000010010",
33005=>"000000000",
33006=>"000000000",
33007=>"000000000",
33008=>"000000111",
33009=>"111000000",
33010=>"011001111",
33011=>"011010010",
33012=>"000100011",
33013=>"111111111",
33014=>"100000000",
33015=>"000001000",
33016=>"111000000",
33017=>"001111111",
33018=>"111100100",
33019=>"000010001",
33020=>"001000000",
33021=>"000111111",
33022=>"011111111",
33023=>"100111111",
33024=>"011011111",
33025=>"011010100",
33026=>"100000111",
33027=>"000000111",
33028=>"000100101",
33029=>"111000000",
33030=>"100100111",
33031=>"000111110",
33032=>"000000000",
33033=>"001000000",
33034=>"011010011",
33035=>"000100000",
33036=>"111111101",
33037=>"000011111",
33038=>"100100111",
33039=>"101000000",
33040=>"000000011",
33041=>"000111111",
33042=>"100000100",
33043=>"110000000",
33044=>"001000011",
33045=>"000111000",
33046=>"011001000",
33047=>"010111111",
33048=>"011010000",
33049=>"011101001",
33050=>"001011010",
33051=>"001000000",
33052=>"111000111",
33053=>"101010000",
33054=>"110010000",
33055=>"100101100",
33056=>"000111010",
33057=>"001101000",
33058=>"000000000",
33059=>"000101011",
33060=>"111111110",
33061=>"110110001",
33062=>"000011010",
33063=>"101000010",
33064=>"000010010",
33065=>"010111000",
33066=>"100000000",
33067=>"111111000",
33068=>"111111100",
33069=>"111000000",
33070=>"111011111",
33071=>"001000010",
33072=>"010011010",
33073=>"000010011",
33074=>"101111010",
33075=>"111111000",
33076=>"000010000",
33077=>"000100000",
33078=>"111110100",
33079=>"000000110",
33080=>"011010011",
33081=>"000000000",
33082=>"000000010",
33083=>"101010011",
33084=>"100100000",
33085=>"010101000",
33086=>"000101101",
33087=>"000001011",
33088=>"011110001",
33089=>"111001000",
33090=>"010011000",
33091=>"001001011",
33092=>"111111100",
33093=>"000000000",
33094=>"111010000",
33095=>"100111111",
33096=>"000001110",
33097=>"000110011",
33098=>"000101100",
33099=>"001000001",
33100=>"100000010",
33101=>"100100110",
33102=>"001001111",
33103=>"111100110",
33104=>"010000100",
33105=>"010000000",
33106=>"111001101",
33107=>"011011011",
33108=>"000011111",
33109=>"011111001",
33110=>"001111011",
33111=>"000000000",
33112=>"111000001",
33113=>"010000001",
33114=>"000000010",
33115=>"011011001",
33116=>"111111111",
33117=>"000001000",
33118=>"111101000",
33119=>"100000011",
33120=>"111111011",
33121=>"001000111",
33122=>"111101001",
33123=>"110010000",
33124=>"001101101",
33125=>"000000000",
33126=>"000010111",
33127=>"000000000",
33128=>"111111111",
33129=>"010000010",
33130=>"111000001",
33131=>"110000101",
33132=>"000111000",
33133=>"100111111",
33134=>"000000100",
33135=>"000000000",
33136=>"000100110",
33137=>"111011000",
33138=>"011011000",
33139=>"011110100",
33140=>"110100111",
33141=>"001000000",
33142=>"010000010",
33143=>"111101000",
33144=>"111111010",
33145=>"110000111",
33146=>"111101000",
33147=>"001011111",
33148=>"010001111",
33149=>"010110010",
33150=>"001111111",
33151=>"000011111",
33152=>"111011000",
33153=>"010010010",
33154=>"000000010",
33155=>"101001000",
33156=>"000000000",
33157=>"100010111",
33158=>"011001100",
33159=>"011000110",
33160=>"100001011",
33161=>"000010111",
33162=>"000011011",
33163=>"000111110",
33164=>"000000110",
33165=>"000111111",
33166=>"111101000",
33167=>"111001001",
33168=>"001001001",
33169=>"101111010",
33170=>"100111111",
33171=>"000001010",
33172=>"111111111",
33173=>"100000000",
33174=>"111100000",
33175=>"000110110",
33176=>"010111000",
33177=>"101010101",
33178=>"000010010",
33179=>"111111010",
33180=>"111100111",
33181=>"111111000",
33182=>"011111000",
33183=>"001001010",
33184=>"001000000",
33185=>"111110000",
33186=>"000011100",
33187=>"000011011",
33188=>"110111000",
33189=>"110100000",
33190=>"010000001",
33191=>"110110100",
33192=>"111000000",
33193=>"001011010",
33194=>"001101110",
33195=>"000001101",
33196=>"111101100",
33197=>"101001011",
33198=>"010101001",
33199=>"011000000",
33200=>"001101000",
33201=>"110110110",
33202=>"100000000",
33203=>"000000000",
33204=>"000111111",
33205=>"010000100",
33206=>"010011101",
33207=>"111000100",
33208=>"001000001",
33209=>"010111011",
33210=>"111010000",
33211=>"000011011",
33212=>"001001101",
33213=>"111111111",
33214=>"000110111",
33215=>"111111000",
33216=>"100100100",
33217=>"010011111",
33218=>"111111000",
33219=>"110111110",
33220=>"111011010",
33221=>"100111001",
33222=>"110011010",
33223=>"001111111",
33224=>"111000000",
33225=>"000010000",
33226=>"111010100",
33227=>"010011101",
33228=>"000010011",
33229=>"110100010",
33230=>"000101000",
33231=>"010000111",
33232=>"000000010",
33233=>"110111010",
33234=>"010010000",
33235=>"111100100",
33236=>"111111010",
33237=>"011011011",
33238=>"111111111",
33239=>"000000011",
33240=>"101001000",
33241=>"000011111",
33242=>"100100000",
33243=>"000000010",
33244=>"111100000",
33245=>"000100110",
33246=>"011011101",
33247=>"001000000",
33248=>"001001111",
33249=>"111011000",
33250=>"100000000",
33251=>"011110110",
33252=>"111011011",
33253=>"111111000",
33254=>"000000000",
33255=>"000011000",
33256=>"000111001",
33257=>"110110101",
33258=>"010011110",
33259=>"101101001",
33260=>"011001000",
33261=>"111111110",
33262=>"000000010",
33263=>"000000000",
33264=>"000111011",
33265=>"011001100",
33266=>"111011000",
33267=>"100111111",
33268=>"010111011",
33269=>"111101111",
33270=>"000000001",
33271=>"100000000",
33272=>"001001101",
33273=>"011100000",
33274=>"010111101",
33275=>"111110111",
33276=>"111000000",
33277=>"000110111",
33278=>"001101100",
33279=>"010000000",
33280=>"111000000",
33281=>"000000100",
33282=>"000100111",
33283=>"000000000",
33284=>"100110101",
33285=>"000000111",
33286=>"000010111",
33287=>"100110111",
33288=>"001001001",
33289=>"111000000",
33290=>"100110000",
33291=>"000000000",
33292=>"111001000",
33293=>"000000000",
33294=>"110011000",
33295=>"001000000",
33296=>"111010110",
33297=>"000010110",
33298=>"100010111",
33299=>"000111111",
33300=>"000010011",
33301=>"000100111",
33302=>"111001110",
33303=>"010010000",
33304=>"101000000",
33305=>"011010011",
33306=>"100100000",
33307=>"000110111",
33308=>"110000111",
33309=>"110110110",
33310=>"111010110",
33311=>"000100100",
33312=>"000000010",
33313=>"000000000",
33314=>"000000111",
33315=>"111101111",
33316=>"011000000",
33317=>"011000000",
33318=>"101111100",
33319=>"111111111",
33320=>"111111010",
33321=>"100100000",
33322=>"101111001",
33323=>"110111111",
33324=>"010011001",
33325=>"110101111",
33326=>"111111111",
33327=>"000011001",
33328=>"000000000",
33329=>"110010110",
33330=>"000001111",
33331=>"011000000",
33332=>"000111111",
33333=>"000101000",
33334=>"011011011",
33335=>"000000111",
33336=>"000000000",
33337=>"000001011",
33338=>"000011011",
33339=>"011000000",
33340=>"111100100",
33341=>"010000001",
33342=>"111100000",
33343=>"000011001",
33344=>"111000111",
33345=>"010010011",
33346=>"000111111",
33347=>"000000000",
33348=>"000011010",
33349=>"111100000",
33350=>"010000011",
33351=>"110001101",
33352=>"110101110",
33353=>"111111100",
33354=>"100110001",
33355=>"101110010",
33356=>"111000000",
33357=>"110000011",
33358=>"011000001",
33359=>"010100111",
33360=>"111001111",
33361=>"111001101",
33362=>"000010011",
33363=>"011001000",
33364=>"101000000",
33365=>"111011000",
33366=>"100110011",
33367=>"000001111",
33368=>"111011010",
33369=>"111100000",
33370=>"001010000",
33371=>"000000100",
33372=>"111011000",
33373=>"011110000",
33374=>"011111111",
33375=>"001100101",
33376=>"001001000",
33377=>"011110111",
33378=>"101000000",
33379=>"100000100",
33380=>"011111000",
33381=>"000101001",
33382=>"000110010",
33383=>"000110100",
33384=>"111010000",
33385=>"000100110",
33386=>"111111010",
33387=>"000010111",
33388=>"000111000",
33389=>"000011111",
33390=>"000000111",
33391=>"000000000",
33392=>"111100000",
33393=>"000000100",
33394=>"110110110",
33395=>"001000110",
33396=>"011111111",
33397=>"100000000",
33398=>"000010000",
33399=>"100000101",
33400=>"000000010",
33401=>"111111111",
33402=>"000111101",
33403=>"011010000",
33404=>"001010001",
33405=>"111110000",
33406=>"100111111",
33407=>"000000010",
33408=>"110110000",
33409=>"000000000",
33410=>"100100100",
33411=>"000110111",
33412=>"011001000",
33413=>"000100110",
33414=>"110000001",
33415=>"000100100",
33416=>"010010010",
33417=>"000011011",
33418=>"110011010",
33419=>"000100111",
33420=>"000101101",
33421=>"000000000",
33422=>"111000000",
33423=>"010001001",
33424=>"110011111",
33425=>"111010110",
33426=>"100000010",
33427=>"111111100",
33428=>"010111011",
33429=>"111000000",
33430=>"111011000",
33431=>"111000000",
33432=>"101111000",
33433=>"101000111",
33434=>"000000000",
33435=>"011001001",
33436=>"111101100",
33437=>"111011000",
33438=>"000000000",
33439=>"110111010",
33440=>"011010010",
33441=>"110100010",
33442=>"000111111",
33443=>"101010111",
33444=>"111011111",
33445=>"110011011",
33446=>"110000101",
33447=>"000111111",
33448=>"010110111",
33449=>"000100000",
33450=>"111000000",
33451=>"000010100",
33452=>"000000011",
33453=>"111101001",
33454=>"111010001",
33455=>"000000010",
33456=>"111000000",
33457=>"010110111",
33458=>"111000000",
33459=>"100101001",
33460=>"111100100",
33461=>"000100000",
33462=>"001000000",
33463=>"000000000",
33464=>"011001011",
33465=>"100001010",
33466=>"111100000",
33467=>"000101000",
33468=>"010010111",
33469=>"111011111",
33470=>"110100100",
33471=>"000100011",
33472=>"000111111",
33473=>"010001101",
33474=>"101101101",
33475=>"110011111",
33476=>"000100100",
33477=>"011011100",
33478=>"000100000",
33479=>"111111111",
33480=>"110001111",
33481=>"000000000",
33482=>"000010111",
33483=>"111000000",
33484=>"000100010",
33485=>"010011001",
33486=>"110110000",
33487=>"111000000",
33488=>"000111111",
33489=>"111110001",
33490=>"000100000",
33491=>"011111101",
33492=>"000000110",
33493=>"001001001",
33494=>"111101111",
33495=>"000100001",
33496=>"100111000",
33497=>"000011000",
33498=>"010010001",
33499=>"111000000",
33500=>"111100001",
33501=>"011000101",
33502=>"001001001",
33503=>"000000000",
33504=>"000100111",
33505=>"000110111",
33506=>"010000000",
33507=>"001011111",
33508=>"100000000",
33509=>"000000001",
33510=>"000011111",
33511=>"111101000",
33512=>"111110100",
33513=>"000110010",
33514=>"001011110",
33515=>"000000111",
33516=>"000101111",
33517=>"000000000",
33518=>"000000101",
33519=>"111001000",
33520=>"101110000",
33521=>"111010100",
33522=>"110000100",
33523=>"111001000",
33524=>"011100100",
33525=>"000000111",
33526=>"111101101",
33527=>"011111000",
33528=>"100111110",
33529=>"010111011",
33530=>"111000111",
33531=>"000001001",
33532=>"111000000",
33533=>"010000000",
33534=>"011010010",
33535=>"011111111",
33536=>"100001010",
33537=>"110011011",
33538=>"111001001",
33539=>"000000110",
33540=>"110000000",
33541=>"010110000",
33542=>"100110110",
33543=>"000001111",
33544=>"001111011",
33545=>"011001001",
33546=>"000100000",
33547=>"110100100",
33548=>"000100110",
33549=>"011001000",
33550=>"101001000",
33551=>"111100100",
33552=>"001001001",
33553=>"000000111",
33554=>"110011000",
33555=>"110110010",
33556=>"110001101",
33557=>"001100110",
33558=>"011000011",
33559=>"110011001",
33560=>"011001001",
33561=>"001000011",
33562=>"000010010",
33563=>"000011111",
33564=>"000010010",
33565=>"010111110",
33566=>"101111000",
33567=>"001110110",
33568=>"001001101",
33569=>"011111010",
33570=>"111101110",
33571=>"000110110",
33572=>"100100000",
33573=>"001001011",
33574=>"001110110",
33575=>"000000011",
33576=>"001111110",
33577=>"000100110",
33578=>"001110011",
33579=>"001001001",
33580=>"000101110",
33581=>"100100111",
33582=>"010111001",
33583=>"000001111",
33584=>"100110110",
33585=>"001111111",
33586=>"011011010",
33587=>"111001000",
33588=>"101001110",
33589=>"110110110",
33590=>"101001001",
33591=>"110001111",
33592=>"111001100",
33593=>"111001011",
33594=>"000111100",
33595=>"000011011",
33596=>"001110101",
33597=>"111111000",
33598=>"000000001",
33599=>"000110110",
33600=>"001001001",
33601=>"001001011",
33602=>"111001000",
33603=>"001111111",
33604=>"011001010",
33605=>"000110011",
33606=>"110000110",
33607=>"110110000",
33608=>"111100100",
33609=>"110011100",
33610=>"000000111",
33611=>"001001000",
33612=>"111001111",
33613=>"000101100",
33614=>"000100100",
33615=>"001101101",
33616=>"011001001",
33617=>"010101000",
33618=>"110000110",
33619=>"110011011",
33620=>"111001001",
33621=>"110000011",
33622=>"111110110",
33623=>"111001001",
33624=>"010110100",
33625=>"110111111",
33626=>"000001001",
33627=>"000100000",
33628=>"000001000",
33629=>"000010011",
33630=>"111001011",
33631=>"000101000",
33632=>"000110110",
33633=>"010110111",
33634=>"001001001",
33635=>"111111001",
33636=>"010001110",
33637=>"000000100",
33638=>"110100000",
33639=>"011000011",
33640=>"000100110",
33641=>"110110001",
33642=>"000101101",
33643=>"010001110",
33644=>"110011111",
33645=>"000000001",
33646=>"001001100",
33647=>"000111111",
33648=>"111111011",
33649=>"000000000",
33650=>"000001001",
33651=>"000110000",
33652=>"001001011",
33653=>"010001001",
33654=>"101000000",
33655=>"001001001",
33656=>"000011001",
33657=>"111110010",
33658=>"111001000",
33659=>"000111100",
33660=>"111000011",
33661=>"101000000",
33662=>"001001001",
33663=>"001100100",
33664=>"110111001",
33665=>"000110000",
33666=>"000110100",
33667=>"000110001",
33668=>"000110010",
33669=>"110001000",
33670=>"000001111",
33671=>"111001101",
33672=>"110110110",
33673=>"001000000",
33674=>"000001001",
33675=>"110100001",
33676=>"011001001",
33677=>"011001001",
33678=>"100000000",
33679=>"001001111",
33680=>"101101110",
33681=>"001000111",
33682=>"001001000",
33683=>"111110011",
33684=>"101000000",
33685=>"011001100",
33686=>"001110010",
33687=>"000110111",
33688=>"000110000",
33689=>"001111000",
33690=>"100110100",
33691=>"111011001",
33692=>"111111000",
33693=>"111001001",
33694=>"111110111",
33695=>"001110000",
33696=>"111111101",
33697=>"011001001",
33698=>"011001001",
33699=>"110111011",
33700=>"110110000",
33701=>"000000111",
33702=>"100100000",
33703=>"000000100",
33704=>"110100110",
33705=>"110100110",
33706=>"000100100",
33707=>"001111001",
33708=>"110110010",
33709=>"011001000",
33710=>"010000011",
33711=>"101001001",
33712=>"000010100",
33713=>"000010111",
33714=>"000011001",
33715=>"101011001",
33716=>"010110100",
33717=>"111011111",
33718=>"110110101",
33719=>"001001011",
33720=>"000110100",
33721=>"110010011",
33722=>"010011000",
33723=>"110110001",
33724=>"110110110",
33725=>"111111110",
33726=>"000111101",
33727=>"000111001",
33728=>"111001001",
33729=>"101001011",
33730=>"111110110",
33731=>"001100100",
33732=>"000100010",
33733=>"000110110",
33734=>"110001001",
33735=>"000110001",
33736=>"000110001",
33737=>"000000110",
33738=>"110011011",
33739=>"000000110",
33740=>"011001001",
33741=>"111001001",
33742=>"011001001",
33743=>"010111111",
33744=>"100100000",
33745=>"000100100",
33746=>"111100011",
33747=>"000100010",
33748=>"001001001",
33749=>"011001100",
33750=>"011000101",
33751=>"000111110",
33752=>"100100110",
33753=>"110110110",
33754=>"001101001",
33755=>"110001001",
33756=>"001001000",
33757=>"001111010",
33758=>"110111110",
33759=>"010101001",
33760=>"001001111",
33761=>"111011001",
33762=>"101100000",
33763=>"011111111",
33764=>"101001101",
33765=>"011001001",
33766=>"000110110",
33767=>"000110011",
33768=>"010010000",
33769=>"100100111",
33770=>"001000000",
33771=>"100001011",
33772=>"001010100",
33773=>"000110110",
33774=>"010001111",
33775=>"000110110",
33776=>"110110110",
33777=>"110000101",
33778=>"100101000",
33779=>"100100000",
33780=>"000110101",
33781=>"111001001",
33782=>"000000010",
33783=>"110000000",
33784=>"111001011",
33785=>"110000010",
33786=>"110001001",
33787=>"000111110",
33788=>"000110110",
33789=>"011001001",
33790=>"110101001",
33791=>"111001001",
33792=>"000001100",
33793=>"010000000",
33794=>"001001111",
33795=>"000000110",
33796=>"001001101",
33797=>"010001011",
33798=>"110101111",
33799=>"000000001",
33800=>"000010100",
33801=>"001100111",
33802=>"010101001",
33803=>"110100010",
33804=>"000000001",
33805=>"001001001",
33806=>"011011011",
33807=>"111001000",
33808=>"010110100",
33809=>"000000100",
33810=>"001111110",
33811=>"000110110",
33812=>"111111111",
33813=>"010010110",
33814=>"000000001",
33815=>"000110110",
33816=>"110111111",
33817=>"111111011",
33818=>"000000000",
33819=>"000000001",
33820=>"110110000",
33821=>"000101110",
33822=>"000000011",
33823=>"001001101",
33824=>"001101111",
33825=>"000001010",
33826=>"001000000",
33827=>"001000100",
33828=>"101100100",
33829=>"111101010",
33830=>"000101111",
33831=>"111000101",
33832=>"001001111",
33833=>"011100011",
33834=>"000000000",
33835=>"001000100",
33836=>"010001000",
33837=>"111111111",
33838=>"010100011",
33839=>"110001010",
33840=>"000000000",
33841=>"101111011",
33842=>"000001111",
33843=>"001001011",
33844=>"110110100",
33845=>"111101110",
33846=>"111011111",
33847=>"110111000",
33848=>"011000110",
33849=>"001001000",
33850=>"111111100",
33851=>"000000100",
33852=>"010000000",
33853=>"111011010",
33854=>"000000011",
33855=>"100101111",
33856=>"110111111",
33857=>"110110000",
33858=>"001000000",
33859=>"011000100",
33860=>"000001000",
33861=>"001101111",
33862=>"110110000",
33863=>"001111111",
33864=>"101011010",
33865=>"111101001",
33866=>"000001011",
33867=>"110110000",
33868=>"111001111",
33869=>"011111011",
33870=>"100111101",
33871=>"001010110",
33872=>"000010010",
33873=>"101000111",
33874=>"011111111",
33875=>"011011010",
33876=>"010110000",
33877=>"000001010",
33878=>"010011010",
33879=>"000010111",
33880=>"011011000",
33881=>"000001001",
33882=>"000101000",
33883=>"011111000",
33884=>"000000000",
33885=>"001000001",
33886=>"110010110",
33887=>"100001011",
33888=>"101101111",
33889=>"000000000",
33890=>"001000101",
33891=>"000001110",
33892=>"000000000",
33893=>"111111101",
33894=>"100101011",
33895=>"001101111",
33896=>"111101111",
33897=>"000111111",
33898=>"001111111",
33899=>"000000100",
33900=>"000001000",
33901=>"110110111",
33902=>"000100110",
33903=>"010000000",
33904=>"001011001",
33905=>"000000000",
33906=>"001000100",
33907=>"111111000",
33908=>"000000000",
33909=>"101001000",
33910=>"111010010",
33911=>"111000001",
33912=>"001000110",
33913=>"011111111",
33914=>"111010000",
33915=>"110001011",
33916=>"110010010",
33917=>"100000010",
33918=>"111110110",
33919=>"001001001",
33920=>"111100000",
33921=>"010000000",
33922=>"111000100",
33923=>"110010111",
33924=>"001001100",
33925=>"111111101",
33926=>"011011001",
33927=>"011001000",
33928=>"000000000",
33929=>"000000001",
33930=>"010111101",
33931=>"000000110",
33932=>"000000100",
33933=>"110110110",
33934=>"111011000",
33935=>"111000000",
33936=>"111010110",
33937=>"011111100",
33938=>"000000010",
33939=>"000110111",
33940=>"110111101",
33941=>"001000110",
33942=>"111111000",
33943=>"100100010",
33944=>"111101111",
33945=>"010001111",
33946=>"111010111",
33947=>"111111111",
33948=>"011111111",
33949=>"010010000",
33950=>"110110000",
33951=>"000100111",
33952=>"101100110",
33953=>"111001111",
33954=>"000000010",
33955=>"101111001",
33956=>"010110110",
33957=>"110111000",
33958=>"000000111",
33959=>"111101000",
33960=>"010110010",
33961=>"101010110",
33962=>"111111010",
33963=>"001000110",
33964=>"111111111",
33965=>"000000010",
33966=>"110000000",
33967=>"111111110",
33968=>"110000011",
33969=>"010111001",
33970=>"111001001",
33971=>"001000100",
33972=>"000001010",
33973=>"000011000",
33974=>"111101000",
33975=>"100000000",
33976=>"011010010",
33977=>"110110010",
33978=>"111101110",
33979=>"101111111",
33980=>"000100101",
33981=>"111111111",
33982=>"010011111",
33983=>"000000000",
33984=>"110110110",
33985=>"010110000",
33986=>"110000000",
33987=>"011110100",
33988=>"110001001",
33989=>"001101001",
33990=>"000111110",
33991=>"000000001",
33992=>"111100110",
33993=>"001001001",
33994=>"001000000",
33995=>"111111000",
33996=>"000101000",
33997=>"011101100",
33998=>"000010000",
33999=>"101101111",
34000=>"010110010",
34001=>"011011111",
34002=>"110000000",
34003=>"111110000",
34004=>"010000101",
34005=>"000000010",
34006=>"001001111",
34007=>"110011010",
34008=>"000100110",
34009=>"000110110",
34010=>"011001001",
34011=>"000110000",
34012=>"000000001",
34013=>"101101010",
34014=>"111111000",
34015=>"001101100",
34016=>"001001101",
34017=>"101001001",
34018=>"010000000",
34019=>"110110001",
34020=>"001001111",
34021=>"000000001",
34022=>"110110111",
34023=>"010110111",
34024=>"001001111",
34025=>"010110110",
34026=>"010100100",
34027=>"011110010",
34028=>"000001101",
34029=>"110100000",
34030=>"000000000",
34031=>"000000001",
34032=>"000000000",
34033=>"000011100",
34034=>"001000011",
34035=>"000001111",
34036=>"000111011",
34037=>"011000000",
34038=>"110100010",
34039=>"010000010",
34040=>"110010000",
34041=>"000001111",
34042=>"010110000",
34043=>"010111110",
34044=>"111111110",
34045=>"010111111",
34046=>"111111011",
34047=>"111111001",
34048=>"000000000",
34049=>"000000000",
34050=>"111000111",
34051=>"010000111",
34052=>"000000000",
34053=>"111111011",
34054=>"000000100",
34055=>"000000000",
34056=>"000010011",
34057=>"000000111",
34058=>"000000100",
34059=>"011100100",
34060=>"011011111",
34061=>"101000101",
34062=>"110000100",
34063=>"110000000",
34064=>"111011011",
34065=>"101111000",
34066=>"100000110",
34067=>"011111000",
34068=>"111011001",
34069=>"000001001",
34070=>"000000000",
34071=>"111111100",
34072=>"000010011",
34073=>"101000000",
34074=>"000000010",
34075=>"000000111",
34076=>"011111011",
34077=>"000101000",
34078=>"100111010",
34079=>"101100100",
34080=>"111000101",
34081=>"000000000",
34082=>"000100001",
34083=>"111100111",
34084=>"100110110",
34085=>"100000010",
34086=>"111110000",
34087=>"000101011",
34088=>"111111111",
34089=>"001111111",
34090=>"000000000",
34091=>"001111111",
34092=>"000011011",
34093=>"111010100",
34094=>"100111000",
34095=>"000000000",
34096=>"101111010",
34097=>"011000100",
34098=>"000000000",
34099=>"101111000",
34100=>"000000111",
34101=>"100110000",
34102=>"010000011",
34103=>"000100111",
34104=>"100111111",
34105=>"000000000",
34106=>"111000000",
34107=>"100111111",
34108=>"100001101",
34109=>"111101101",
34110=>"000110010",
34111=>"000010011",
34112=>"001111011",
34113=>"000001010",
34114=>"001011000",
34115=>"000100110",
34116=>"101000000",
34117=>"000111111",
34118=>"000000000",
34119=>"100100000",
34120=>"010011111",
34121=>"100000011",
34122=>"110010110",
34123=>"010111011",
34124=>"011111111",
34125=>"000001011",
34126=>"100000000",
34127=>"111111100",
34128=>"000000111",
34129=>"101100101",
34130=>"000111000",
34131=>"100010110",
34132=>"110000100",
34133=>"001001111",
34134=>"011110100",
34135=>"101101101",
34136=>"001001000",
34137=>"000011001",
34138=>"011011011",
34139=>"000111011",
34140=>"000111010",
34141=>"111000100",
34142=>"101000101",
34143=>"100000011",
34144=>"111011111",
34145=>"100100000",
34146=>"010010111",
34147=>"111110110",
34148=>"010111101",
34149=>"010010010",
34150=>"100000000",
34151=>"100100111",
34152=>"001000110",
34153=>"000000110",
34154=>"000111111",
34155=>"010000010",
34156=>"111111000",
34157=>"000111000",
34158=>"111111010",
34159=>"000000000",
34160=>"010011011",
34161=>"111111011",
34162=>"001000110",
34163=>"000100000",
34164=>"000111111",
34165=>"110100111",
34166=>"000000000",
34167=>"111111111",
34168=>"101001000",
34169=>"000111111",
34170=>"111111000",
34171=>"101000100",
34172=>"011001100",
34173=>"000001001",
34174=>"101100111",
34175=>"011100111",
34176=>"100011111",
34177=>"111111000",
34178=>"000011010",
34179=>"100100111",
34180=>"000010000",
34181=>"111111111",
34182=>"001010110",
34183=>"110100001",
34184=>"111010010",
34185=>"000000000",
34186=>"111111101",
34187=>"001001111",
34188=>"111111011",
34189=>"000111010",
34190=>"000110111",
34191=>"011000000",
34192=>"001000011",
34193=>"100111111",
34194=>"101000000",
34195=>"000000000",
34196=>"010000010",
34197=>"001111011",
34198=>"111000001",
34199=>"110111111",
34200=>"000111011",
34201=>"101101101",
34202=>"111000100",
34203=>"100011111",
34204=>"000011011",
34205=>"100111000",
34206=>"010111111",
34207=>"111111111",
34208=>"101111111",
34209=>"111111000",
34210=>"010000111",
34211=>"111000000",
34212=>"000111110",
34213=>"000110110",
34214=>"000111011",
34215=>"010111011",
34216=>"000111111",
34217=>"111011111",
34218=>"101000001",
34219=>"010111111",
34220=>"101101001",
34221=>"010110011",
34222=>"100101101",
34223=>"111111000",
34224=>"100111101",
34225=>"110011100",
34226=>"000010000",
34227=>"011011000",
34228=>"100010110",
34229=>"000010000",
34230=>"000000100",
34231=>"010000011",
34232=>"100100101",
34233=>"010000000",
34234=>"100001000",
34235=>"001111111",
34236=>"100111000",
34237=>"111100101",
34238=>"000010000",
34239=>"101000111",
34240=>"111111011",
34241=>"010110010",
34242=>"111001000",
34243=>"111110111",
34244=>"001100000",
34245=>"110111011",
34246=>"100111000",
34247=>"001000001",
34248=>"001000000",
34249=>"011011111",
34250=>"000000000",
34251=>"111000000",
34252=>"111111111",
34253=>"111100101",
34254=>"010000000",
34255=>"001111110",
34256=>"110111011",
34257=>"001011011",
34258=>"111111000",
34259=>"111110010",
34260=>"000000000",
34261=>"001000001",
34262=>"011010010",
34263=>"011011011",
34264=>"001000100",
34265=>"100011111",
34266=>"111010010",
34267=>"010111010",
34268=>"000000110",
34269=>"100111001",
34270=>"000010000",
34271=>"100000110",
34272=>"000101010",
34273=>"111111110",
34274=>"100000100",
34275=>"100110111",
34276=>"010000001",
34277=>"000101100",
34278=>"010011010",
34279=>"000001101",
34280=>"011010000",
34281=>"110000111",
34282=>"000000000",
34283=>"000000001",
34284=>"111111111",
34285=>"000100000",
34286=>"100111111",
34287=>"111000100",
34288=>"000000000",
34289=>"001110011",
34290=>"000101111",
34291=>"000011011",
34292=>"000100000",
34293=>"010010010",
34294=>"010011010",
34295=>"011000000",
34296=>"101101101",
34297=>"100000100",
34298=>"111111011",
34299=>"000100101",
34300=>"101111101",
34301=>"000011010",
34302=>"000010110",
34303=>"111011111",
34304=>"111001100",
34305=>"000000000",
34306=>"111101100",
34307=>"101010100",
34308=>"000000010",
34309=>"001011100",
34310=>"000001001",
34311=>"000000001",
34312=>"000000000",
34313=>"010100000",
34314=>"000100110",
34315=>"000011110",
34316=>"110010000",
34317=>"100001001",
34318=>"100010000",
34319=>"101010011",
34320=>"101000000",
34321=>"111000100",
34322=>"001110100",
34323=>"011001111",
34324=>"111100110",
34325=>"111000110",
34326=>"001110111",
34327=>"111101111",
34328=>"111010000",
34329=>"100000011",
34330=>"000110011",
34331=>"000100110",
34332=>"000000011",
34333=>"000000100",
34334=>"010111100",
34335=>"111100011",
34336=>"001000111",
34337=>"001001001",
34338=>"110000011",
34339=>"000000000",
34340=>"000000101",
34341=>"100001001",
34342=>"111100100",
34343=>"000000011",
34344=>"111110100",
34345=>"111011110",
34346=>"000011111",
34347=>"111111100",
34348=>"000010011",
34349=>"000010000",
34350=>"000000110",
34351=>"000001011",
34352=>"110100100",
34353=>"101011011",
34354=>"111000100",
34355=>"101111111",
34356=>"001011111",
34357=>"110111111",
34358=>"000110000",
34359=>"100110100",
34360=>"000011011",
34361=>"111100000",
34362=>"111100000",
34363=>"001110110",
34364=>"100100001",
34365=>"010011111",
34366=>"111100100",
34367=>"000001000",
34368=>"100100100",
34369=>"010111111",
34370=>"000011011",
34371=>"010110100",
34372=>"111000000",
34373=>"000001001",
34374=>"001100100",
34375=>"111001001",
34376=>"000110111",
34377=>"000011111",
34378=>"001111110",
34379=>"010110111",
34380=>"010100110",
34381=>"110111010",
34382=>"110100101",
34383=>"100001111",
34384=>"111110001",
34385=>"011100111",
34386=>"111011110",
34387=>"001011001",
34388=>"000000000",
34389=>"001000111",
34390=>"100000010",
34391=>"010011000",
34392=>"100100111",
34393=>"010001011",
34394=>"100111101",
34395=>"010000101",
34396=>"000000000",
34397=>"010100100",
34398=>"111010110",
34399=>"111100100",
34400=>"110100000",
34401=>"100110111",
34402=>"111110100",
34403=>"000000110",
34404=>"100010001",
34405=>"100100110",
34406=>"000000001",
34407=>"111011000",
34408=>"011110100",
34409=>"000000111",
34410=>"011010000",
34411=>"111110111",
34412=>"111110100",
34413=>"010111111",
34414=>"010001001",
34415=>"011011111",
34416=>"000011111",
34417=>"000100000",
34418=>"111000100",
34419=>"000101001",
34420=>"010100111",
34421=>"101100100",
34422=>"000010011",
34423=>"100111100",
34424=>"101000010",
34425=>"010001111",
34426=>"011111111",
34427=>"000000101",
34428=>"110011011",
34429=>"100101010",
34430=>"001100100",
34431=>"011010000",
34432=>"110011000",
34433=>"001011100",
34434=>"011001001",
34435=>"000001000",
34436=>"000100111",
34437=>"011110000",
34438=>"010010011",
34439=>"000000010",
34440=>"110101110",
34441=>"111000000",
34442=>"101111000",
34443=>"000001111",
34444=>"111110100",
34445=>"000000000",
34446=>"100111001",
34447=>"000100000",
34448=>"110010011",
34449=>"101111011",
34450=>"100000011",
34451=>"111111100",
34452=>"000100011",
34453=>"011100100",
34454=>"110010111",
34455=>"110111111",
34456=>"001111111",
34457=>"100110011",
34458=>"000010011",
34459=>"111100101",
34460=>"000000000",
34461=>"111110000",
34462=>"000011000",
34463=>"111110000",
34464=>"000010001",
34465=>"111111111",
34466=>"100101011",
34467=>"010010000",
34468=>"000000011",
34469=>"000100111",
34470=>"100000000",
34471=>"000001011",
34472=>"111111100",
34473=>"001011001",
34474=>"110100100",
34475=>"111011000",
34476=>"100011111",
34477=>"000011011",
34478=>"111111110",
34479=>"011101000",
34480=>"001011000",
34481=>"000100100",
34482=>"001111110",
34483=>"000001000",
34484=>"100000011",
34485=>"010111011",
34486=>"000011011",
34487=>"010011011",
34488=>"000111001",
34489=>"000000111",
34490=>"000011011",
34491=>"010011001",
34492=>"000111011",
34493=>"011110111",
34494=>"000001010",
34495=>"010000001",
34496=>"111100100",
34497=>"000001001",
34498=>"000011011",
34499=>"000011011",
34500=>"000000011",
34501=>"100100111",
34502=>"111011011",
34503=>"000001111",
34504=>"000001010",
34505=>"011111000",
34506=>"100110011",
34507=>"111100100",
34508=>"110111110",
34509=>"011110011",
34510=>"001001001",
34511=>"100001000",
34512=>"010110000",
34513=>"000010110",
34514=>"110100000",
34515=>"010110111",
34516=>"111100100",
34517=>"110100010",
34518=>"001001100",
34519=>"110011011",
34520=>"000010011",
34521=>"110000000",
34522=>"100110111",
34523=>"011100100",
34524=>"110111010",
34525=>"011000111",
34526=>"000011011",
34527=>"000000100",
34528=>"111000001",
34529=>"111110100",
34530=>"011000100",
34531=>"111011110",
34532=>"010111010",
34533=>"001000011",
34534=>"000011011",
34535=>"111111110",
34536=>"000100110",
34537=>"000100011",
34538=>"000100000",
34539=>"101011011",
34540=>"110011011",
34541=>"011111110",
34542=>"010000000",
34543=>"000001100",
34544=>"110100100",
34545=>"000010111",
34546=>"011001100",
34547=>"000010010",
34548=>"001001110",
34549=>"100100100",
34550=>"011100000",
34551=>"000000000",
34552=>"000000111",
34553=>"000001001",
34554=>"011011111",
34555=>"011000111",
34556=>"111100100",
34557=>"001000110",
34558=>"000011111",
34559=>"010111100",
34560=>"111110110",
34561=>"000000001",
34562=>"111111110",
34563=>"100111001",
34564=>"111111100",
34565=>"110010001",
34566=>"000010110",
34567=>"110111110",
34568=>"111111000",
34569=>"111001001",
34570=>"001001011",
34571=>"111111001",
34572=>"111010000",
34573=>"000101000",
34574=>"111011000",
34575=>"000000010",
34576=>"000110010",
34577=>"000000000",
34578=>"000000001",
34579=>"010000010",
34580=>"000011010",
34581=>"111111110",
34582=>"000000110",
34583=>"111110010",
34584=>"010000011",
34585=>"000100111",
34586=>"001000000",
34587=>"000000011",
34588=>"101011111",
34589=>"101000011",
34590=>"111011101",
34591=>"101000000",
34592=>"000111111",
34593=>"111011001",
34594=>"111011000",
34595=>"111000111",
34596=>"011101100",
34597=>"101011010",
34598=>"000000101",
34599=>"000000000",
34600=>"000100110",
34601=>"111111111",
34602=>"111000000",
34603=>"000110111",
34604=>"011011000",
34605=>"100111101",
34606=>"000000000",
34607=>"001101111",
34608=>"011111111",
34609=>"101101001",
34610=>"000101000",
34611=>"000111111",
34612=>"010110000",
34613=>"111111111",
34614=>"000001010",
34615=>"111001100",
34616=>"110111111",
34617=>"111001000",
34618=>"101011000",
34619=>"000111110",
34620=>"011000011",
34621=>"001011011",
34622=>"000000000",
34623=>"101000000",
34624=>"110010110",
34625=>"110011001",
34626=>"010010101",
34627=>"001000100",
34628=>"010000000",
34629=>"010010001",
34630=>"011000000",
34631=>"000001100",
34632=>"111011111",
34633=>"000011111",
34634=>"110111101",
34635=>"111111000",
34636=>"111111111",
34637=>"101001000",
34638=>"111101010",
34639=>"111110000",
34640=>"001001001",
34641=>"100111010",
34642=>"111000000",
34643=>"111100111",
34644=>"000000001",
34645=>"100101001",
34646=>"000010011",
34647=>"000001111",
34648=>"111101001",
34649=>"001001000",
34650=>"111000001",
34651=>"001010000",
34652=>"100010110",
34653=>"100000100",
34654=>"011111110",
34655=>"000011111",
34656=>"010000000",
34657=>"001000000",
34658=>"100000000",
34659=>"011000000",
34660=>"111000000",
34661=>"111001000",
34662=>"001111111",
34663=>"001111111",
34664=>"110011111",
34665=>"000000101",
34666=>"001001011",
34667=>"111111000",
34668=>"000110100",
34669=>"000011111",
34670=>"000000101",
34671=>"000000000",
34672=>"011111110",
34673=>"001111111",
34674=>"000100111",
34675=>"111010011",
34676=>"101000110",
34677=>"001101001",
34678=>"011111100",
34679=>"111111100",
34680=>"000000111",
34681=>"000000111",
34682=>"001101010",
34683=>"101111000",
34684=>"101100010",
34685=>"110100011",
34686=>"000111111",
34687=>"110000000",
34688=>"000010001",
34689=>"111111000",
34690=>"000010110",
34691=>"111111000",
34692=>"111000011",
34693=>"101111111",
34694=>"010100001",
34695=>"011011010",
34696=>"011111011",
34697=>"000001101",
34698=>"000111111",
34699=>"010010011",
34700=>"000101111",
34701=>"000011111",
34702=>"001000100",
34703=>"001000000",
34704=>"000001011",
34705=>"101000000",
34706=>"000111011",
34707=>"111101000",
34708=>"111101100",
34709=>"000101001",
34710=>"110000000",
34711=>"100111100",
34712=>"111101100",
34713=>"000000111",
34714=>"000100111",
34715=>"100000000",
34716=>"111111000",
34717=>"101000000",
34718=>"000001001",
34719=>"110110000",
34720=>"000000010",
34721=>"000111011",
34722=>"000111000",
34723=>"110000101",
34724=>"110111101",
34725=>"001000000",
34726=>"111110000",
34727=>"000010110",
34728=>"000111111",
34729=>"000010101",
34730=>"011111101",
34731=>"010000000",
34732=>"001111000",
34733=>"110100000",
34734=>"101011011",
34735=>"011110000",
34736=>"111100110",
34737=>"111101010",
34738=>"100011000",
34739=>"001001100",
34740=>"100111001",
34741=>"111110110",
34742=>"111111000",
34743=>"111111111",
34744=>"100000110",
34745=>"001000001",
34746=>"111011011",
34747=>"000001110",
34748=>"111101101",
34749=>"111000111",
34750=>"111100000",
34751=>"001111111",
34752=>"111010000",
34753=>"011000000",
34754=>"011011101",
34755=>"111001100",
34756=>"100000111",
34757=>"001100111",
34758=>"110100111",
34759=>"111011000",
34760=>"011111100",
34761=>"111001001",
34762=>"110000001",
34763=>"111000001",
34764=>"000000000",
34765=>"010001010",
34766=>"001000000",
34767=>"100000100",
34768=>"010000001",
34769=>"001001000",
34770=>"111000001",
34771=>"100111011",
34772=>"111000000",
34773=>"001000010",
34774=>"110000000",
34775=>"000000100",
34776=>"110111111",
34777=>"100000111",
34778=>"001000001",
34779=>"001100111",
34780=>"000111110",
34781=>"111111101",
34782=>"111111000",
34783=>"111110100",
34784=>"111000000",
34785=>"111011000",
34786=>"111011000",
34787=>"110000000",
34788=>"101000010",
34789=>"111111000",
34790=>"100110000",
34791=>"110110010",
34792=>"000000000",
34793=>"000110111",
34794=>"100000010",
34795=>"011000000",
34796=>"110111000",
34797=>"000000000",
34798=>"010010000",
34799=>"111000000",
34800=>"000000111",
34801=>"001001010",
34802=>"111001001",
34803=>"011000000",
34804=>"111010111",
34805=>"001000101",
34806=>"111000000",
34807=>"001000111",
34808=>"010111000",
34809=>"001111110",
34810=>"000000000",
34811=>"001000101",
34812=>"111010111",
34813=>"001111111",
34814=>"111000000",
34815=>"011000000",
34816=>"001100100",
34817=>"011100000",
34818=>"110100100",
34819=>"111111111",
34820=>"011000000",
34821=>"001111111",
34822=>"000111000",
34823=>"110111111",
34824=>"000000000",
34825=>"000001010",
34826=>"000000111",
34827=>"101000000",
34828=>"111010000",
34829=>"000000000",
34830=>"101000000",
34831=>"000000110",
34832=>"000000000",
34833=>"011111000",
34834=>"111000000",
34835=>"111111000",
34836=>"001000000",
34837=>"111000010",
34838=>"010000111",
34839=>"111111001",
34840=>"001010000",
34841=>"000000000",
34842=>"011000100",
34843=>"101100110",
34844=>"100000001",
34845=>"000000000",
34846=>"001100111",
34847=>"000111110",
34848=>"111111111",
34849=>"010000100",
34850=>"001101000",
34851=>"011111111",
34852=>"110111111",
34853=>"000101001",
34854=>"010111001",
34855=>"110110000",
34856=>"000001110",
34857=>"111000000",
34858=>"100000000",
34859=>"010100101",
34860=>"001010000",
34861=>"011000001",
34862=>"111100100",
34863=>"000110111",
34864=>"111000010",
34865=>"111111110",
34866=>"000000110",
34867=>"100110011",
34868=>"101000110",
34869=>"111111000",
34870=>"000001111",
34871=>"000000111",
34872=>"001111111",
34873=>"101100000",
34874=>"000010111",
34875=>"111111111",
34876=>"111100100",
34877=>"111111111",
34878=>"000000000",
34879=>"111010011",
34880=>"010001111",
34881=>"000101011",
34882=>"000111111",
34883=>"000000001",
34884=>"111000000",
34885=>"111000000",
34886=>"000000000",
34887=>"011011000",
34888=>"001111111",
34889=>"110110000",
34890=>"000000000",
34891=>"111010000",
34892=>"111000111",
34893=>"011000110",
34894=>"110111011",
34895=>"101111000",
34896=>"111110110",
34897=>"100111010",
34898=>"111111111",
34899=>"000000000",
34900=>"110000001",
34901=>"111110110",
34902=>"111011000",
34903=>"010111001",
34904=>"010011001",
34905=>"101011110",
34906=>"000010110",
34907=>"001011000",
34908=>"001111000",
34909=>"000000010",
34910=>"000111111",
34911=>"000000010",
34912=>"000000101",
34913=>"111000000",
34914=>"100000111",
34915=>"001011001",
34916=>"110100010",
34917=>"100000010",
34918=>"111000100",
34919=>"111111000",
34920=>"000100111",
34921=>"100110010",
34922=>"001001000",
34923=>"000100111",
34924=>"100100111",
34925=>"111111111",
34926=>"011011100",
34927=>"111100000",
34928=>"100100011",
34929=>"000000000",
34930=>"000000011",
34931=>"110000000",
34932=>"000111100",
34933=>"100000000",
34934=>"100101001",
34935=>"000000000",
34936=>"000001011",
34937=>"111111111",
34938=>"000000000",
34939=>"111111111",
34940=>"100100100",
34941=>"000000000",
34942=>"000011110",
34943=>"010000000",
34944=>"011100000",
34945=>"010101011",
34946=>"010000000",
34947=>"011111111",
34948=>"111001000",
34949=>"000000010",
34950=>"010111100",
34951=>"111110010",
34952=>"111100110",
34953=>"111000000",
34954=>"111011000",
34955=>"000000000",
34956=>"000000011",
34957=>"110000111",
34958=>"000111011",
34959=>"111000000",
34960=>"111110001",
34961=>"000000111",
34962=>"000111111",
34963=>"000000000",
34964=>"000011000",
34965=>"000111011",
34966=>"000000000",
34967=>"110000011",
34968=>"000111101",
34969=>"010011000",
34970=>"000010000",
34971=>"000000000",
34972=>"111111000",
34973=>"101101000",
34974=>"001100000",
34975=>"000100000",
34976=>"011100011",
34977=>"000000111",
34978=>"010000000",
34979=>"111111111",
34980=>"000000111",
34981=>"111001000",
34982=>"111000110",
34983=>"000111110",
34984=>"111000000",
34985=>"000000111",
34986=>"000000000",
34987=>"000100110",
34988=>"110011000",
34989=>"110000000",
34990=>"100001011",
34991=>"111111111",
34992=>"100000100",
34993=>"001000111",
34994=>"100000110",
34995=>"000000000",
34996=>"011001011",
34997=>"010000000",
34998=>"001100010",
34999=>"001000000",
35000=>"111100010",
35001=>"001000000",
35002=>"010101111",
35003=>"100010000",
35004=>"111111010",
35005=>"100001111",
35006=>"111111100",
35007=>"111010000",
35008=>"111000100",
35009=>"110100101",
35010=>"000000000",
35011=>"001011100",
35012=>"000000000",
35013=>"010000000",
35014=>"000110000",
35015=>"111111111",
35016=>"111111101",
35017=>"000000110",
35018=>"110110101",
35019=>"111110100",
35020=>"011110000",
35021=>"110101000",
35022=>"000000100",
35023=>"101111111",
35024=>"111101000",
35025=>"001110110",
35026=>"000100000",
35027=>"001000000",
35028=>"110111110",
35029=>"100000101",
35030=>"100100111",
35031=>"000000010",
35032=>"111111100",
35033=>"000000011",
35034=>"110010001",
35035=>"100000000",
35036=>"111101100",
35037=>"111111000",
35038=>"000001000",
35039=>"001110110",
35040=>"000100000",
35041=>"000000000",
35042=>"011001011",
35043=>"111011011",
35044=>"010010100",
35045=>"111000000",
35046=>"010101101",
35047=>"000110110",
35048=>"000001000",
35049=>"111110001",
35050=>"010000100",
35051=>"000100111",
35052=>"000100111",
35053=>"100000000",
35054=>"010110000",
35055=>"000000000",
35056=>"111100000",
35057=>"011000000",
35058=>"011000000",
35059=>"000110000",
35060=>"001001000",
35061=>"100000000",
35062=>"100000000",
35063=>"000011111",
35064=>"000000000",
35065=>"001011100",
35066=>"111010000",
35067=>"000000010",
35068=>"111011000",
35069=>"010111111",
35070=>"000000001",
35071=>"100111101",
35072=>"011111011",
35073=>"000111111",
35074=>"001000101",
35075=>"000000000",
35076=>"001011011",
35077=>"000000100",
35078=>"000000000",
35079=>"000111111",
35080=>"110010111",
35081=>"000000000",
35082=>"110111000",
35083=>"000001111",
35084=>"000000011",
35085=>"000000001",
35086=>"111111010",
35087=>"000001011",
35088=>"111001000",
35089=>"011111000",
35090=>"101000100",
35091=>"000111111",
35092=>"101010100",
35093=>"000101100",
35094=>"111001100",
35095=>"000010010",
35096=>"010010000",
35097=>"111001101",
35098=>"110011000",
35099=>"000000000",
35100=>"000000100",
35101=>"000010010",
35102=>"111110000",
35103=>"000010111",
35104=>"111000111",
35105=>"110110000",
35106=>"000000000",
35107=>"011000000",
35108=>"000000000",
35109=>"011011110",
35110=>"010011000",
35111=>"111110001",
35112=>"111001101",
35113=>"010010000",
35114=>"001000000",
35115=>"000110101",
35116=>"001011011",
35117=>"110000011",
35118=>"111011000",
35119=>"000001001",
35120=>"010000100",
35121=>"011011001",
35122=>"111101001",
35123=>"000000000",
35124=>"111010000",
35125=>"000000001",
35126=>"011111100",
35127=>"000000101",
35128=>"000111111",
35129=>"111111111",
35130=>"101000100",
35131=>"000000111",
35132=>"100110000",
35133=>"111111000",
35134=>"000000101",
35135=>"110011011",
35136=>"111000000",
35137=>"011111111",
35138=>"111111000",
35139=>"000100110",
35140=>"111011010",
35141=>"000111111",
35142=>"001101000",
35143=>"111100111",
35144=>"000011011",
35145=>"110010010",
35146=>"101000111",
35147=>"000010000",
35148=>"001111111",
35149=>"101111000",
35150=>"110110110",
35151=>"000111111",
35152=>"110111111",
35153=>"011111111",
35154=>"011000001",
35155=>"001000000",
35156=>"000000010",
35157=>"010000011",
35158=>"111110010",
35159=>"001001000",
35160=>"000110000",
35161=>"001000011",
35162=>"000011011",
35163=>"110110110",
35164=>"111101000",
35165=>"001011010",
35166=>"010000111",
35167=>"000001110",
35168=>"110010000",
35169=>"100100101",
35170=>"111001110",
35171=>"000110100",
35172=>"101110000",
35173=>"111100111",
35174=>"111111001",
35175=>"110000111",
35176=>"001100000",
35177=>"000111000",
35178=>"111010000",
35179=>"000001000",
35180=>"100110111",
35181=>"110110101",
35182=>"101101111",
35183=>"000010111",
35184=>"011011000",
35185=>"010000000",
35186=>"110111011",
35187=>"000001111",
35188=>"111110000",
35189=>"110111100",
35190=>"111111111",
35191=>"011000001",
35192=>"000101111",
35193=>"111000000",
35194=>"111101000",
35195=>"000100001",
35196=>"100110111",
35197=>"110100000",
35198=>"000010110",
35199=>"110000010",
35200=>"111111101",
35201=>"000000000",
35202=>"001010111",
35203=>"110000101",
35204=>"111110010",
35205=>"111101111",
35206=>"100110111",
35207=>"111110000",
35208=>"111110000",
35209=>"000110000",
35210=>"100000001",
35211=>"110111001",
35212=>"100100001",
35213=>"000000011",
35214=>"001000101",
35215=>"110111001",
35216=>"011011000",
35217=>"010011010",
35218=>"000000100",
35219=>"010000000",
35220=>"111011001",
35221=>"111111000",
35222=>"010010001",
35223=>"011000001",
35224=>"111011101",
35225=>"000111111",
35226=>"000000101",
35227=>"100000111",
35228=>"101100111",
35229=>"110100111",
35230=>"010000111",
35231=>"000000011",
35232=>"001100100",
35233=>"101000111",
35234=>"111011000",
35235=>"111101101",
35236=>"111010000",
35237=>"111111110",
35238=>"110111111",
35239=>"010111111",
35240=>"000111111",
35241=>"001111111",
35242=>"000000111",
35243=>"010111111",
35244=>"111101111",
35245=>"111000111",
35246=>"100010010",
35247=>"110100101",
35248=>"000101001",
35249=>"000011000",
35250=>"000110100",
35251=>"100110010",
35252=>"110010011",
35253=>"111111010",
35254=>"011010100",
35255=>"011110000",
35256=>"001001111",
35257=>"110110001",
35258=>"010010000",
35259=>"010010000",
35260=>"100100000",
35261=>"111111000",
35262=>"010000010",
35263=>"111110000",
35264=>"001001101",
35265=>"001101100",
35266=>"111111000",
35267=>"100100100",
35268=>"111101101",
35269=>"110011000",
35270=>"000111111",
35271=>"111101000",
35272=>"011111001",
35273=>"000100111",
35274=>"011011000",
35275=>"101101110",
35276=>"011110011",
35277=>"011011111",
35278=>"000000100",
35279=>"110110000",
35280=>"000111000",
35281=>"100100000",
35282=>"000000101",
35283=>"111101111",
35284=>"101101011",
35285=>"110110110",
35286=>"000001111",
35287=>"000111111",
35288=>"000000111",
35289=>"101111111",
35290=>"001001001",
35291=>"000000111",
35292=>"011100010",
35293=>"000111111",
35294=>"010010000",
35295=>"000110111",
35296=>"111001010",
35297=>"011000000",
35298=>"110000000",
35299=>"101111000",
35300=>"010000110",
35301=>"010010000",
35302=>"111110111",
35303=>"011100110",
35304=>"111000000",
35305=>"001111111",
35306=>"011111001",
35307=>"111111000",
35308=>"111101111",
35309=>"000000111",
35310=>"101100000",
35311=>"001100000",
35312=>"000000111",
35313=>"011010000",
35314=>"000101111",
35315=>"000000000",
35316=>"110011100",
35317=>"010010010",
35318=>"111000111",
35319=>"111100111",
35320=>"111001010",
35321=>"000001001",
35322=>"110010000",
35323=>"101011000",
35324=>"100101110",
35325=>"100000100",
35326=>"100100000",
35327=>"100111000",
35328=>"110111111",
35329=>"101000000",
35330=>"101000000",
35331=>"000000000",
35332=>"001111101",
35333=>"111011111",
35334=>"000000000",
35335=>"101111111",
35336=>"000111001",
35337=>"001001000",
35338=>"100000100",
35339=>"101001111",
35340=>"110110111",
35341=>"000000000",
35342=>"110100011",
35343=>"000101110",
35344=>"010110111",
35345=>"000000000",
35346=>"010100001",
35347=>"111100000",
35348=>"111111101",
35349=>"111101001",
35350=>"011100000",
35351=>"111000000",
35352=>"100000101",
35353=>"001110011",
35354=>"000111101",
35355=>"000000111",
35356=>"010111110",
35357=>"010000001",
35358=>"111011111",
35359=>"110111001",
35360=>"000000110",
35361=>"010111001",
35362=>"111101100",
35363=>"010110111",
35364=>"110111101",
35365=>"011111111",
35366=>"111001001",
35367=>"100011110",
35368=>"111111111",
35369=>"001111111",
35370=>"001000010",
35371=>"011000000",
35372=>"111111100",
35373=>"101101100",
35374=>"000000000",
35375=>"000000000",
35376=>"000111111",
35377=>"000110111",
35378=>"111111111",
35379=>"000111111",
35380=>"101000000",
35381=>"000000000",
35382=>"001010011",
35383=>"111111010",
35384=>"111111111",
35385=>"010100110",
35386=>"001000000",
35387=>"000000000",
35388=>"011011001",
35389=>"000111101",
35390=>"000000100",
35391=>"000001110",
35392=>"111001111",
35393=>"101011111",
35394=>"011011010",
35395=>"011011001",
35396=>"000000000",
35397=>"101110000",
35398=>"111000101",
35399=>"011000000",
35400=>"101110111",
35401=>"110111111",
35402=>"000010101",
35403=>"100111011",
35404=>"111000101",
35405=>"010110001",
35406=>"000110111",
35407=>"000000010",
35408=>"101000100",
35409=>"101111111",
35410=>"111111111",
35411=>"000000110",
35412=>"000000100",
35413=>"111110110",
35414=>"000111111",
35415=>"111000010",
35416=>"000000000",
35417=>"011111101",
35418=>"011111100",
35419=>"111111111",
35420=>"000000100",
35421=>"100000000",
35422=>"111111111",
35423=>"000110000",
35424=>"000011000",
35425=>"110111111",
35426=>"000000000",
35427=>"100000000",
35428=>"011111111",
35429=>"011011111",
35430=>"110011111",
35431=>"000011101",
35432=>"011001000",
35433=>"111011110",
35434=>"000001100",
35435=>"111111101",
35436=>"000000001",
35437=>"000000000",
35438=>"010011000",
35439=>"101010111",
35440=>"000011001",
35441=>"001001101",
35442=>"100000100",
35443=>"100111111",
35444=>"010001100",
35445=>"111111000",
35446=>"110000000",
35447=>"101110111",
35448=>"010000000",
35449=>"000000000",
35450=>"001111101",
35451=>"000101111",
35452=>"001110100",
35453=>"000100000",
35454=>"100000010",
35455=>"001101111",
35456=>"000010010",
35457=>"000110000",
35458=>"000001101",
35459=>"110010101",
35460=>"101001111",
35461=>"001000000",
35462=>"110100101",
35463=>"000000100",
35464=>"000101100",
35465=>"001001000",
35466=>"111000000",
35467=>"100000100",
35468=>"000111000",
35469=>"111000000",
35470=>"000001111",
35471=>"001001010",
35472=>"111101000",
35473=>"111101101",
35474=>"000000011",
35475=>"000000110",
35476=>"000000010",
35477=>"100111111",
35478=>"111101111",
35479=>"100111101",
35480=>"111111110",
35481=>"111001000",
35482=>"100000000",
35483=>"001000000",
35484=>"110110010",
35485=>"000000000",
35486=>"010111001",
35487=>"101001101",
35488=>"000001111",
35489=>"001000000",
35490=>"000000000",
35491=>"111101111",
35492=>"010111111",
35493=>"110110000",
35494=>"111110110",
35495=>"111110111",
35496=>"111011100",
35497=>"010000000",
35498=>"101101111",
35499=>"110001101",
35500=>"000000100",
35501=>"101011111",
35502=>"001101000",
35503=>"111101011",
35504=>"000001100",
35505=>"001111011",
35506=>"000100011",
35507=>"001001111",
35508=>"110011101",
35509=>"111111000",
35510=>"100100010",
35511=>"111010101",
35512=>"110111110",
35513=>"000000110",
35514=>"111000111",
35515=>"110001001",
35516=>"100111001",
35517=>"101111110",
35518=>"111111111",
35519=>"111000100",
35520=>"111000011",
35521=>"101000000",
35522=>"111111101",
35523=>"010110100",
35524=>"111010000",
35525=>"000000000",
35526=>"111111011",
35527=>"100111110",
35528=>"000000101",
35529=>"000101000",
35530=>"100000000",
35531=>"000010000",
35532=>"000000000",
35533=>"000011111",
35534=>"101000000",
35535=>"010100100",
35536=>"110111000",
35537=>"010111101",
35538=>"101000001",
35539=>"100111000",
35540=>"111101100",
35541=>"001011001",
35542=>"001001001",
35543=>"111111111",
35544=>"111001000",
35545=>"000000000",
35546=>"000000000",
35547=>"001000100",
35548=>"111011001",
35549=>"110000101",
35550=>"101111110",
35551=>"111111111",
35552=>"100010001",
35553=>"111111111",
35554=>"001001011",
35555=>"000001100",
35556=>"010100000",
35557=>"111111101",
35558=>"111001000",
35559=>"000011011",
35560=>"000001011",
35561=>"100011110",
35562=>"101000001",
35563=>"101101001",
35564=>"111111101",
35565=>"101110111",
35566=>"000011000",
35567=>"000100110",
35568=>"101000100",
35569=>"001000010",
35570=>"111111111",
35571=>"000111111",
35572=>"000110011",
35573=>"000000001",
35574=>"100001001",
35575=>"110000111",
35576=>"101111111",
35577=>"111111111",
35578=>"000111101",
35579=>"000000000",
35580=>"000111111",
35581=>"000000100",
35582=>"101101111",
35583=>"011000000",
35584=>"001010011",
35585=>"000100000",
35586=>"101000000",
35587=>"001111010",
35588=>"010011111",
35589=>"110110000",
35590=>"110110110",
35591=>"111001001",
35592=>"000110111",
35593=>"000000001",
35594=>"111001111",
35595=>"001001001",
35596=>"000110110",
35597=>"000111111",
35598=>"100000100",
35599=>"110111110",
35600=>"111001001",
35601=>"111101111",
35602=>"010110010",
35603=>"111101100",
35604=>"111101101",
35605=>"001000110",
35606=>"101000111",
35607=>"101101000",
35608=>"110101111",
35609=>"010001001",
35610=>"000001001",
35611=>"000000100",
35612=>"000101111",
35613=>"110111111",
35614=>"000000000",
35615=>"110000010",
35616=>"110111100",
35617=>"010110111",
35618=>"000000111",
35619=>"000110110",
35620=>"111011001",
35621=>"101000000",
35622=>"000001011",
35623=>"111001111",
35624=>"000000000",
35625=>"001001001",
35626=>"100000000",
35627=>"110111000",
35628=>"100001001",
35629=>"111000111",
35630=>"111000001",
35631=>"000000000",
35632=>"001100111",
35633=>"011111011",
35634=>"000110111",
35635=>"101101111",
35636=>"000000101",
35637=>"000001110",
35638=>"000110111",
35639=>"111101001",
35640=>"111111101",
35641=>"111000000",
35642=>"111000000",
35643=>"111000000",
35644=>"011100000",
35645=>"110110111",
35646=>"001000000",
35647=>"000110010",
35648=>"001000011",
35649=>"000001000",
35650=>"000111111",
35651=>"010110000",
35652=>"000110110",
35653=>"111110000",
35654=>"000110110",
35655=>"110100000",
35656=>"110110111",
35657=>"001000101",
35658=>"110001101",
35659=>"111101001",
35660=>"101101111",
35661=>"110111010",
35662=>"110111001",
35663=>"011000001",
35664=>"000011111",
35665=>"111010000",
35666=>"111000000",
35667=>"011001001",
35668=>"001000001",
35669=>"111110110",
35670=>"101011111",
35671=>"101000000",
35672=>"110010000",
35673=>"011110111",
35674=>"111000000",
35675=>"101100100",
35676=>"100000000",
35677=>"011000010",
35678=>"111111110",
35679=>"010110100",
35680=>"000000111",
35681=>"000000000",
35682=>"001001001",
35683=>"111011001",
35684=>"111000000",
35685=>"000011111",
35686=>"101001000",
35687=>"001000001",
35688=>"111001001",
35689=>"111010111",
35690=>"000010000",
35691=>"110100001",
35692=>"111111101",
35693=>"111001000",
35694=>"110110010",
35695=>"001001111",
35696=>"011100101",
35697=>"001000111",
35698=>"001010111",
35699=>"111001111",
35700=>"110001000",
35701=>"000001001",
35702=>"111111001",
35703=>"000111110",
35704=>"101001001",
35705=>"110111001",
35706=>"001001101",
35707=>"010111111",
35708=>"111100000",
35709=>"100100000",
35710=>"111110001",
35711=>"000110110",
35712=>"000000111",
35713=>"111000000",
35714=>"000111111",
35715=>"000100000",
35716=>"011001000",
35717=>"000001001",
35718=>"011111011",
35719=>"111001000",
35720=>"110011011",
35721=>"111001001",
35722=>"111001000",
35723=>"111110000",
35724=>"000110110",
35725=>"011111111",
35726=>"010010010",
35727=>"111001001",
35728=>"110110100",
35729=>"001111111",
35730=>"000111111",
35731=>"000000001",
35732=>"111010000",
35733=>"001111110",
35734=>"110001001",
35735=>"000011011",
35736=>"010110001",
35737=>"110000000",
35738=>"011111111",
35739=>"010010110",
35740=>"000110110",
35741=>"111111010",
35742=>"001001111",
35743=>"001001001",
35744=>"011110111",
35745=>"000001000",
35746=>"010000000",
35747=>"000000110",
35748=>"000110111",
35749=>"100001011",
35750=>"001000000",
35751=>"000010110",
35752=>"111111111",
35753=>"001010100",
35754=>"101101000",
35755=>"001001000",
35756=>"101100001",
35757=>"111111010",
35758=>"111100100",
35759=>"111110110",
35760=>"111110000",
35761=>"100010000",
35762=>"111000000",
35763=>"110000000",
35764=>"011001111",
35765=>"000000110",
35766=>"000000110",
35767=>"000110011",
35768=>"000100111",
35769=>"010010001",
35770=>"000000000",
35771=>"100000000",
35772=>"111111111",
35773=>"011110110",
35774=>"001111011",
35775=>"111110111",
35776=>"001000001",
35777=>"011101111",
35778=>"000111111",
35779=>"011111011",
35780=>"000000000",
35781=>"111000000",
35782=>"010110101",
35783=>"011000001",
35784=>"000000001",
35785=>"101000001",
35786=>"000010110",
35787=>"111011111",
35788=>"111001000",
35789=>"010000000",
35790=>"011001101",
35791=>"000000000",
35792=>"010000010",
35793=>"010110110",
35794=>"001000001",
35795=>"110010010",
35796=>"101001101",
35797=>"110001110",
35798=>"100000100",
35799=>"110110000",
35800=>"111001001",
35801=>"000000110",
35802=>"110111011",
35803=>"101001001",
35804=>"001001111",
35805=>"111001010",
35806=>"000001101",
35807=>"111111111",
35808=>"101000000",
35809=>"001010011",
35810=>"001000000",
35811=>"000011001",
35812=>"000101101",
35813=>"110000000",
35814=>"000110110",
35815=>"000001011",
35816=>"110111111",
35817=>"111111101",
35818=>"111100101",
35819=>"000000111",
35820=>"000000000",
35821=>"010111111",
35822=>"111011000",
35823=>"000000000",
35824=>"010000001",
35825=>"111000011",
35826=>"001000000",
35827=>"110000111",
35828=>"000101100",
35829=>"101000000",
35830=>"011000101",
35831=>"111101000",
35832=>"000000000",
35833=>"110101100",
35834=>"111010000",
35835=>"000101100",
35836=>"111110101",
35837=>"000000000",
35838=>"110110110",
35839=>"111001101",
35840=>"100010000",
35841=>"000000001",
35842=>"011001111",
35843=>"011111000",
35844=>"000100000",
35845=>"000010001",
35846=>"000010010",
35847=>"101110011",
35848=>"000110100",
35849=>"111101110",
35850=>"011000001",
35851=>"000000000",
35852=>"000111010",
35853=>"111101001",
35854=>"101001000",
35855=>"000000011",
35856=>"110111001",
35857=>"111100111",
35858=>"111100000",
35859=>"111101101",
35860=>"010101111",
35861=>"111101111",
35862=>"101000101",
35863=>"011100101",
35864=>"110101010",
35865=>"000110110",
35866=>"000111111",
35867=>"000010000",
35868=>"111011001",
35869=>"101101111",
35870=>"011011000",
35871=>"101000000",
35872=>"011101001",
35873=>"010000100",
35874=>"111000000",
35875=>"000111010",
35876=>"110000011",
35877=>"000000000",
35878=>"000100111",
35879=>"110100010",
35880=>"000010110",
35881=>"010111011",
35882=>"111010100",
35883=>"010010011",
35884=>"000011000",
35885=>"000001000",
35886=>"101111111",
35887=>"100010000",
35888=>"010001001",
35889=>"111100110",
35890=>"111110100",
35891=>"101101000",
35892=>"000001101",
35893=>"100000000",
35894=>"110001111",
35895=>"001111000",
35896=>"111001100",
35897=>"000000000",
35898=>"000110111",
35899=>"100101001",
35900=>"011110110",
35901=>"111111111",
35902=>"100000111",
35903=>"111110111",
35904=>"111011110",
35905=>"000000001",
35906=>"101111010",
35907=>"111001000",
35908=>"000100111",
35909=>"000000000",
35910=>"111111111",
35911=>"010000101",
35912=>"101000000",
35913=>"110011001",
35914=>"101001101",
35915=>"111101001",
35916=>"111000100",
35917=>"011110000",
35918=>"111100101",
35919=>"110111010",
35920=>"101101101",
35921=>"111111111",
35922=>"101000001",
35923=>"000000000",
35924=>"011010000",
35925=>"111000001",
35926=>"110011001",
35927=>"000000011",
35928=>"101001001",
35929=>"111100110",
35930=>"111100100",
35931=>"000100010",
35932=>"000000000",
35933=>"000001111",
35934=>"111010110",
35935=>"100000001",
35936=>"111111111",
35937=>"000011111",
35938=>"100100111",
35939=>"110101111",
35940=>"000111000",
35941=>"001001000",
35942=>"110111000",
35943=>"000000000",
35944=>"101111011",
35945=>"100000111",
35946=>"101111111",
35947=>"111111001",
35948=>"000001111",
35949=>"110101000",
35950=>"000001000",
35951=>"000010000",
35952=>"001011001",
35953=>"010001001",
35954=>"111100100",
35955=>"000101000",
35956=>"101111000",
35957=>"001000000",
35958=>"000100000",
35959=>"011000000",
35960=>"010000100",
35961=>"001100000",
35962=>"101010011",
35963=>"100100101",
35964=>"101110110",
35965=>"010000000",
35966=>"100101111",
35967=>"000001101",
35968=>"101001011",
35969=>"010000000",
35970=>"000100100",
35971=>"001110111",
35972=>"100011010",
35973=>"111110001",
35974=>"000000000",
35975=>"101001001",
35976=>"000110110",
35977=>"001100000",
35978=>"010001000",
35979=>"010110111",
35980=>"101000101",
35981=>"111101000",
35982=>"111110110",
35983=>"001000110",
35984=>"000100000",
35985=>"101000000",
35986=>"101000000",
35987=>"011000011",
35988=>"100000000",
35989=>"000000001",
35990=>"110111000",
35991=>"110110000",
35992=>"110111010",
35993=>"011000011",
35994=>"100011101",
35995=>"000000011",
35996=>"011001011",
35997=>"111111111",
35998=>"010010010",
35999=>"101100001",
36000=>"101100110",
36001=>"110001111",
36002=>"110111010",
36003=>"001011000",
36004=>"110011010",
36005=>"100110100",
36006=>"011001001",
36007=>"000010010",
36008=>"110000011",
36009=>"110101111",
36010=>"101100111",
36011=>"010000101",
36012=>"111110100",
36013=>"000000010",
36014=>"000000000",
36015=>"101000000",
36016=>"111001101",
36017=>"101000100",
36018=>"000010010",
36019=>"010010000",
36020=>"111011101",
36021=>"100101110",
36022=>"111111000",
36023=>"111111001",
36024=>"101011000",
36025=>"101100000",
36026=>"010000100",
36027=>"010111100",
36028=>"010010000",
36029=>"111000111",
36030=>"000011011",
36031=>"111101111",
36032=>"001101011",
36033=>"000000000",
36034=>"111111000",
36035=>"110011100",
36036=>"000001011",
36037=>"110100001",
36038=>"000111011",
36039=>"000100000",
36040=>"111111111",
36041=>"100000010",
36042=>"001101111",
36043=>"001000101",
36044=>"111100100",
36045=>"101011011",
36046=>"111111011",
36047=>"111101101",
36048=>"111101111",
36049=>"011110000",
36050=>"000010111",
36051=>"010000000",
36052=>"001000000",
36053=>"011100010",
36054=>"000100100",
36055=>"100010001",
36056=>"000000000",
36057=>"000011111",
36058=>"110001011",
36059=>"111100111",
36060=>"000100100",
36061=>"001111011",
36062=>"010011010",
36063=>"111010000",
36064=>"000101111",
36065=>"011000000",
36066=>"111010111",
36067=>"000001011",
36068=>"001000101",
36069=>"010000011",
36070=>"101001000",
36071=>"000000000",
36072=>"000101011",
36073=>"000000101",
36074=>"110000110",
36075=>"000110111",
36076=>"101111111",
36077=>"111100111",
36078=>"000010100",
36079=>"000000000",
36080=>"000000100",
36081=>"110000000",
36082=>"101011010",
36083=>"001100011",
36084=>"000011011",
36085=>"111101111",
36086=>"000000000",
36087=>"110110111",
36088=>"111111111",
36089=>"110110001",
36090=>"101101101",
36091=>"000001001",
36092=>"000010011",
36093=>"111000000",
36094=>"000011001",
36095=>"111011000",
36096=>"110110110",
36097=>"000101110",
36098=>"101101000",
36099=>"000000110",
36100=>"011011010",
36101=>"010010010",
36102=>"100001111",
36103=>"011000000",
36104=>"010110111",
36105=>"001010000",
36106=>"011110110",
36107=>"111111010",
36108=>"000111111",
36109=>"101000000",
36110=>"000000001",
36111=>"100000111",
36112=>"000000000",
36113=>"110010111",
36114=>"000000000",
36115=>"000000000",
36116=>"111011000",
36117=>"011011000",
36118=>"110110110",
36119=>"111010010",
36120=>"101001110",
36121=>"100001000",
36122=>"110110000",
36123=>"000100110",
36124=>"100000101",
36125=>"111010000",
36126=>"111110000",
36127=>"111111111",
36128=>"111111000",
36129=>"010111000",
36130=>"000000111",
36131=>"110100000",
36132=>"001001001",
36133=>"111101001",
36134=>"000000101",
36135=>"000000000",
36136=>"101000100",
36137=>"010111000",
36138=>"001001000",
36139=>"010011110",
36140=>"000101001",
36141=>"111100000",
36142=>"110111111",
36143=>"010001001",
36144=>"111111111",
36145=>"001011001",
36146=>"110000101",
36147=>"001000001",
36148=>"000010111",
36149=>"111111010",
36150=>"010010000",
36151=>"100100101",
36152=>"010100100",
36153=>"001000100",
36154=>"111101111",
36155=>"110100010",
36156=>"011010000",
36157=>"111111111",
36158=>"000111101",
36159=>"011011011",
36160=>"100101100",
36161=>"010010010",
36162=>"000000000",
36163=>"010011110",
36164=>"101111010",
36165=>"000101111",
36166=>"101000000",
36167=>"101111000",
36168=>"000101001",
36169=>"111101111",
36170=>"101001101",
36171=>"100101100",
36172=>"101011111",
36173=>"110011011",
36174=>"000110110",
36175=>"111011010",
36176=>"111111010",
36177=>"010010000",
36178=>"001011000",
36179=>"111001000",
36180=>"111110010",
36181=>"000110110",
36182=>"110100110",
36183=>"000010010",
36184=>"110111110",
36185=>"001001000",
36186=>"000100000",
36187=>"000100110",
36188=>"100000101",
36189=>"001001001",
36190=>"001000000",
36191=>"010010001",
36192=>"000110011",
36193=>"011010010",
36194=>"000110100",
36195=>"101001001",
36196=>"110111111",
36197=>"000100100",
36198=>"111111011",
36199=>"011111011",
36200=>"111111101",
36201=>"011000000",
36202=>"010111111",
36203=>"000111111",
36204=>"101001001",
36205=>"000000010",
36206=>"000000000",
36207=>"011000110",
36208=>"101000001",
36209=>"000000010",
36210=>"010010000",
36211=>"000000000",
36212=>"111111000",
36213=>"100100111",
36214=>"110011000",
36215=>"111111110",
36216=>"100100010",
36217=>"111000110",
36218=>"100111100",
36219=>"010000000",
36220=>"000110010",
36221=>"111100100",
36222=>"010110001",
36223=>"010110010",
36224=>"000000000",
36225=>"010111000",
36226=>"111000000",
36227=>"101101111",
36228=>"010011101",
36229=>"101101111",
36230=>"110011011",
36231=>"000000000",
36232=>"100111101",
36233=>"110010000",
36234=>"001000000",
36235=>"011010000",
36236=>"010010010",
36237=>"111111010",
36238=>"101001001",
36239=>"111001001",
36240=>"110110100",
36241=>"000000000",
36242=>"000000010",
36243=>"111111000",
36244=>"100001111",
36245=>"000011000",
36246=>"000000000",
36247=>"010111111",
36248=>"011111011",
36249=>"010011011",
36250=>"101000100",
36251=>"101111101",
36252=>"001111111",
36253=>"100000001",
36254=>"111001000",
36255=>"111100001",
36256=>"000000011",
36257=>"000010010",
36258=>"000000100",
36259=>"000111101",
36260=>"111011000",
36261=>"100001100",
36262=>"111111101",
36263=>"100000000",
36264=>"010000111",
36265=>"000100010",
36266=>"000000000",
36267=>"000100100",
36268=>"101011101",
36269=>"101110111",
36270=>"110110100",
36271=>"000000010",
36272=>"000000101",
36273=>"001011000",
36274=>"111010110",
36275=>"100010010",
36276=>"111111011",
36277=>"010000000",
36278=>"000001111",
36279=>"000101010",
36280=>"000001000",
36281=>"000110101",
36282=>"100110000",
36283=>"111111111",
36284=>"010000111",
36285=>"111111111",
36286=>"110110110",
36287=>"011010010",
36288=>"001000101",
36289=>"000010010",
36290=>"101011111",
36291=>"110110100",
36292=>"001000000",
36293=>"110110100",
36294=>"000011111",
36295=>"000000101",
36296=>"000000000",
36297=>"100000001",
36298=>"000000111",
36299=>"110111010",
36300=>"011111001",
36301=>"000010000",
36302=>"010100100",
36303=>"111011101",
36304=>"111110110",
36305=>"010000011",
36306=>"000000000",
36307=>"111100000",
36308=>"101000100",
36309=>"111101110",
36310=>"000000011",
36311=>"000000000",
36312=>"000000000",
36313=>"000000000",
36314=>"000100101",
36315=>"101001000",
36316=>"011110110",
36317=>"011111110",
36318=>"111111111",
36319=>"111111000",
36320=>"110010011",
36321=>"111111100",
36322=>"011111000",
36323=>"111000000",
36324=>"000000111",
36325=>"110111010",
36326=>"000110010",
36327=>"001111100",
36328=>"111100000",
36329=>"011001000",
36330=>"011011011",
36331=>"000110010",
36332=>"010111111",
36333=>"000010111",
36334=>"100010000",
36335=>"100111111",
36336=>"110100100",
36337=>"011010001",
36338=>"000100111",
36339=>"100100100",
36340=>"010110010",
36341=>"111101000",
36342=>"000000000",
36343=>"111010000",
36344=>"100111011",
36345=>"000100000",
36346=>"011000000",
36347=>"111111100",
36348=>"101000101",
36349=>"010111010",
36350=>"110111000",
36351=>"000000000",
36352=>"110100111",
36353=>"110010111",
36354=>"101000100",
36355=>"001000001",
36356=>"010000000",
36357=>"110101111",
36358=>"001000111",
36359=>"000000111",
36360=>"110001001",
36361=>"010000000",
36362=>"100110111",
36363=>"111101100",
36364=>"000000110",
36365=>"010001100",
36366=>"111101100",
36367=>"111111000",
36368=>"010000000",
36369=>"000000111",
36370=>"111101111",
36371=>"000000011",
36372=>"011110111",
36373=>"001110100",
36374=>"010000011",
36375=>"010010101",
36376=>"101100000",
36377=>"000110000",
36378=>"000000001",
36379=>"100010111",
36380=>"110011011",
36381=>"000110100",
36382=>"010101111",
36383=>"000000000",
36384=>"000111000",
36385=>"010100111",
36386=>"101101100",
36387=>"010111000",
36388=>"100000001",
36389=>"111110010",
36390=>"000011010",
36391=>"000000001",
36392=>"111001011",
36393=>"000000111",
36394=>"010000111",
36395=>"000010010",
36396=>"111101100",
36397=>"100000001",
36398=>"110010000",
36399=>"010000000",
36400=>"110001000",
36401=>"110000100",
36402=>"000000011",
36403=>"000001001",
36404=>"010101111",
36405=>"100110110",
36406=>"000110010",
36407=>"111110000",
36408=>"011101110",
36409=>"101000011",
36410=>"111100010",
36411=>"000100100",
36412=>"011110110",
36413=>"111110110",
36414=>"101000000",
36415=>"111100101",
36416=>"011000000",
36417=>"011010111",
36418=>"101000101",
36419=>"111110010",
36420=>"111011010",
36421=>"001000000",
36422=>"010000101",
36423=>"000111011",
36424=>"000011110",
36425=>"111111010",
36426=>"101101001",
36427=>"111000110",
36428=>"000000100",
36429=>"101000011",
36430=>"010000000",
36431=>"111111101",
36432=>"000000111",
36433=>"010010000",
36434=>"000000110",
36435=>"110001010",
36436=>"000010010",
36437=>"111010010",
36438=>"111100110",
36439=>"001000000",
36440=>"000000011",
36441=>"001000000",
36442=>"101101011",
36443=>"110000110",
36444=>"101000110",
36445=>"100101110",
36446=>"111111111",
36447=>"001101010",
36448=>"010000111",
36449=>"000111111",
36450=>"111000010",
36451=>"000110111",
36452=>"111001011",
36453=>"010001011",
36454=>"010111100",
36455=>"110111000",
36456=>"001101100",
36457=>"011100011",
36458=>"000000010",
36459=>"010111000",
36460=>"000111111",
36461=>"101111101",
36462=>"000000101",
36463=>"110001111",
36464=>"000001011",
36465=>"000101101",
36466=>"000011001",
36467=>"000011000",
36468=>"011101001",
36469=>"010001000",
36470=>"101001101",
36471=>"000000000",
36472=>"111000001",
36473=>"000000110",
36474=>"101000001",
36475=>"101100100",
36476=>"100110011",
36477=>"111100010",
36478=>"000111011",
36479=>"101101111",
36480=>"111110000",
36481=>"111000000",
36482=>"000110000",
36483=>"000111111",
36484=>"100000111",
36485=>"110111100",
36486=>"110011001",
36487=>"100100100",
36488=>"000000100",
36489=>"101101101",
36490=>"100000000",
36491=>"000010000",
36492=>"111110000",
36493=>"000000100",
36494=>"101111001",
36495=>"000000001",
36496=>"011011100",
36497=>"000010111",
36498=>"100001000",
36499=>"010110000",
36500=>"101101000",
36501=>"000000100",
36502=>"011011001",
36503=>"110100100",
36504=>"000100101",
36505=>"001110000",
36506=>"000010000",
36507=>"100000111",
36508=>"111100100",
36509=>"000000111",
36510=>"000001000",
36511=>"000010010",
36512=>"011111110",
36513=>"001111010",
36514=>"010011000",
36515=>"000110010",
36516=>"101000111",
36517=>"111100001",
36518=>"000000000",
36519=>"100100111",
36520=>"010010101",
36521=>"101000101",
36522=>"111101011",
36523=>"100000111",
36524=>"010111111",
36525=>"001000000",
36526=>"001011011",
36527=>"000111011",
36528=>"111111000",
36529=>"100001100",
36530=>"111101101",
36531=>"000111011",
36532=>"111111110",
36533=>"000110110",
36534=>"000101000",
36535=>"111000000",
36536=>"100011011",
36537=>"001001001",
36538=>"000111111",
36539=>"111111100",
36540=>"010010110",
36541=>"010001101",
36542=>"000000111",
36543=>"000010010",
36544=>"000110010",
36545=>"000111111",
36546=>"111010000",
36547=>"111001100",
36548=>"001000101",
36549=>"011011000",
36550=>"100100000",
36551=>"010111011",
36552=>"000001001",
36553=>"111010110",
36554=>"011011000",
36555=>"001001101",
36556=>"000010000",
36557=>"101011010",
36558=>"000000000",
36559=>"000111111",
36560=>"111000000",
36561=>"110011010",
36562=>"010000001",
36563=>"000000100",
36564=>"110000101",
36565=>"001100111",
36566=>"101000011",
36567=>"010101010",
36568=>"010010000",
36569=>"000000100",
36570=>"110111001",
36571=>"101000101",
36572=>"000000110",
36573=>"100000000",
36574=>"000000000",
36575=>"111101111",
36576=>"010000101",
36577=>"001000001",
36578=>"011111000",
36579=>"010101011",
36580=>"000000001",
36581=>"000011010",
36582=>"000000001",
36583=>"000101111",
36584=>"111000010",
36585=>"000111101",
36586=>"000001111",
36587=>"001001000",
36588=>"000100111",
36589=>"000101100",
36590=>"001111111",
36591=>"010111011",
36592=>"011000000",
36593=>"111010000",
36594=>"000000001",
36595=>"001100100",
36596=>"001000011",
36597=>"111000111",
36598=>"010000000",
36599=>"110101101",
36600=>"110001000",
36601=>"001110010",
36602=>"011111001",
36603=>"111001110",
36604=>"110011100",
36605=>"000111010",
36606=>"000001010",
36607=>"110000111",
36608=>"000001100",
36609=>"000010000",
36610=>"000000100",
36611=>"000000100",
36612=>"111101100",
36613=>"010101001",
36614=>"100111111",
36615=>"001000011",
36616=>"101111011",
36617=>"000101111",
36618=>"000000001",
36619=>"010111000",
36620=>"000011111",
36621=>"111111110",
36622=>"100000011",
36623=>"011111000",
36624=>"101000001",
36625=>"000000001",
36626=>"000000101",
36627=>"101100111",
36628=>"101101011",
36629=>"111111000",
36630=>"111100100",
36631=>"000001001",
36632=>"000100001",
36633=>"111111111",
36634=>"000101000",
36635=>"100100011",
36636=>"101101011",
36637=>"111111111",
36638=>"110100000",
36639=>"101000000",
36640=>"111101000",
36641=>"111111010",
36642=>"000010100",
36643=>"000000011",
36644=>"100100110",
36645=>"011011011",
36646=>"111011000",
36647=>"000100111",
36648=>"010000000",
36649=>"111111111",
36650=>"110111011",
36651=>"001000010",
36652=>"011111000",
36653=>"100011111",
36654=>"011110000",
36655=>"000000000",
36656=>"101100000",
36657=>"000000100",
36658=>"000100010",
36659=>"001001000",
36660=>"100100001",
36661=>"111111111",
36662=>"110100001",
36663=>"000000000",
36664=>"001011010",
36665=>"100000000",
36666=>"000000000",
36667=>"000111101",
36668=>"010001101",
36669=>"100111101",
36670=>"101101000",
36671=>"011011010",
36672=>"101011111",
36673=>"111101111",
36674=>"000000001",
36675=>"111111101",
36676=>"111110110",
36677=>"100010111",
36678=>"101100100",
36679=>"011111111",
36680=>"011001110",
36681=>"101111111",
36682=>"100100111",
36683=>"111000000",
36684=>"111111010",
36685=>"011011011",
36686=>"010100100",
36687=>"111111011",
36688=>"111000100",
36689=>"010111111",
36690=>"000000000",
36691=>"001010110",
36692=>"000000000",
36693=>"110100000",
36694=>"011111111",
36695=>"000000101",
36696=>"010000000",
36697=>"000000011",
36698=>"110010001",
36699=>"111111010",
36700=>"100000101",
36701=>"000000000",
36702=>"010010000",
36703=>"111111001",
36704=>"111111010",
36705=>"110110010",
36706=>"111101111",
36707=>"110100000",
36708=>"000000110",
36709=>"001000111",
36710=>"000000100",
36711=>"100000111",
36712=>"011011000",
36713=>"111100000",
36714=>"010011010",
36715=>"110100000",
36716=>"000000000",
36717=>"000000000",
36718=>"000000000",
36719=>"000000111",
36720=>"111111100",
36721=>"000101111",
36722=>"011000100",
36723=>"000000110",
36724=>"101111111",
36725=>"100100000",
36726=>"110111100",
36727=>"111110100",
36728=>"011111001",
36729=>"011110100",
36730=>"111011011",
36731=>"000000011",
36732=>"001000010",
36733=>"100100000",
36734=>"100000000",
36735=>"111111111",
36736=>"111111010",
36737=>"110101000",
36738=>"111010011",
36739=>"111111000",
36740=>"111101011",
36741=>"111111110",
36742=>"111100111",
36743=>"011110110",
36744=>"101001000",
36745=>"001011110",
36746=>"100000111",
36747=>"000000000",
36748=>"010010000",
36749=>"011111111",
36750=>"000000001",
36751=>"000001101",
36752=>"100101101",
36753=>"111011011",
36754=>"101101000",
36755=>"101001001",
36756=>"101111101",
36757=>"000000111",
36758=>"010111011",
36759=>"000111010",
36760=>"111101101",
36761=>"111111111",
36762=>"111011111",
36763=>"000000001",
36764=>"000000000",
36765=>"011111111",
36766=>"101111111",
36767=>"000000000",
36768=>"111111110",
36769=>"011111000",
36770=>"101111100",
36771=>"000001100",
36772=>"000000000",
36773=>"110011011",
36774=>"011111011",
36775=>"000000000",
36776=>"000010111",
36777=>"101000000",
36778=>"111111010",
36779=>"100100111",
36780=>"110011100",
36781=>"100000101",
36782=>"000001001",
36783=>"010011111",
36784=>"011110001",
36785=>"001100110",
36786=>"011111011",
36787=>"001000100",
36788=>"100111010",
36789=>"011101000",
36790=>"011111100",
36791=>"111111000",
36792=>"011100111",
36793=>"111101000",
36794=>"000010111",
36795=>"000101111",
36796=>"111101000",
36797=>"111111111",
36798=>"111111111",
36799=>"100101011",
36800=>"000000100",
36801=>"000000000",
36802=>"000001011",
36803=>"100010110",
36804=>"000100010",
36805=>"000000110",
36806=>"111010111",
36807=>"111011010",
36808=>"000000111",
36809=>"010111100",
36810=>"100101101",
36811=>"011111111",
36812=>"000000000",
36813=>"110100000",
36814=>"100101101",
36815=>"000000000",
36816=>"110110110",
36817=>"111111111",
36818=>"111011010",
36819=>"111111111",
36820=>"000000000",
36821=>"000100100",
36822=>"100100011",
36823=>"011011010",
36824=>"101000011",
36825=>"000110000",
36826=>"111111111",
36827=>"000000011",
36828=>"001011001",
36829=>"011100000",
36830=>"011111010",
36831=>"100111010",
36832=>"000000000",
36833=>"000000100",
36834=>"000011111",
36835=>"001100110",
36836=>"000000000",
36837=>"101111000",
36838=>"111111011",
36839=>"011100100",
36840=>"000100111",
36841=>"100101001",
36842=>"000000000",
36843=>"011001100",
36844=>"000000110",
36845=>"010000000",
36846=>"111111000",
36847=>"001000000",
36848=>"110111011",
36849=>"000011111",
36850=>"000111100",
36851=>"101001100",
36852=>"110110000",
36853=>"101000011",
36854=>"000000000",
36855=>"001111011",
36856=>"000010111",
36857=>"100000000",
36858=>"111111111",
36859=>"011101111",
36860=>"111100000",
36861=>"001111011",
36862=>"111111001",
36863=>"000000000",
36864=>"111111100",
36865=>"111111000",
36866=>"000000100",
36867=>"010111000",
36868=>"111111111",
36869=>"000000001",
36870=>"110100011",
36871=>"000000000",
36872=>"000010000",
36873=>"000000000",
36874=>"011011111",
36875=>"001001000",
36876=>"000000000",
36877=>"111111001",
36878=>"100111100",
36879=>"100000001",
36880=>"000000100",
36881=>"000111111",
36882=>"110110001",
36883=>"000010010",
36884=>"010111110",
36885=>"111111111",
36886=>"111111111",
36887=>"111111010",
36888=>"100000000",
36889=>"000000000",
36890=>"000000000",
36891=>"111100111",
36892=>"000000000",
36893=>"110111111",
36894=>"011101111",
36895=>"010011101",
36896=>"000000000",
36897=>"111010111",
36898=>"010001111",
36899=>"011000000",
36900=>"011001011",
36901=>"000000001",
36902=>"110010000",
36903=>"011001001",
36904=>"111111000",
36905=>"110001100",
36906=>"000000001",
36907=>"000001000",
36908=>"001010111",
36909=>"111111111",
36910=>"111111111",
36911=>"000101100",
36912=>"000000000",
36913=>"001000010",
36914=>"001010111",
36915=>"100111111",
36916=>"111111101",
36917=>"111010001",
36918=>"111111000",
36919=>"011011111",
36920=>"010111110",
36921=>"000000110",
36922=>"010000011",
36923=>"001000000",
36924=>"000000000",
36925=>"111111111",
36926=>"000000001",
36927=>"110101001",
36928=>"000000110",
36929=>"000000000",
36930=>"011000000",
36931=>"011000100",
36932=>"111111111",
36933=>"001001001",
36934=>"100101111",
36935=>"111111101",
36936=>"011111111",
36937=>"111001000",
36938=>"000000000",
36939=>"000000000",
36940=>"000000011",
36941=>"000100100",
36942=>"000011111",
36943=>"000000111",
36944=>"010010110",
36945=>"111111111",
36946=>"000010111",
36947=>"001000000",
36948=>"010111100",
36949=>"111111111",
36950=>"000011000",
36951=>"000000000",
36952=>"010110110",
36953=>"111110110",
36954=>"000011111",
36955=>"111011000",
36956=>"111111111",
36957=>"000000000",
36958=>"111111111",
36959=>"000000110",
36960=>"000000000",
36961=>"010111011",
36962=>"000000001",
36963=>"000100011",
36964=>"010011111",
36965=>"011111101",
36966=>"011001010",
36967=>"110111101",
36968=>"111000010",
36969=>"001110010",
36970=>"011111110",
36971=>"111001000",
36972=>"110111001",
36973=>"111111111",
36974=>"011001000",
36975=>"000000000",
36976=>"100111101",
36977=>"111111010",
36978=>"111101100",
36979=>"000000000",
36980=>"001100000",
36981=>"000000000",
36982=>"111101000",
36983=>"000000010",
36984=>"000000101",
36985=>"111011111",
36986=>"111111011",
36987=>"111100100",
36988=>"111100100",
36989=>"110000000",
36990=>"111111111",
36991=>"001000000",
36992=>"000000000",
36993=>"000000000",
36994=>"111010100",
36995=>"110111111",
36996=>"000010111",
36997=>"100101001",
36998=>"000000000",
36999=>"000000000",
37000=>"100001001",
37001=>"000001001",
37002=>"010110010",
37003=>"000000000",
37004=>"101000001",
37005=>"000001011",
37006=>"000110111",
37007=>"000000000",
37008=>"100010111",
37009=>"000010111",
37010=>"111101111",
37011=>"000000000",
37012=>"000000010",
37013=>"000100111",
37014=>"010110000",
37015=>"000100111",
37016=>"000000010",
37017=>"000111111",
37018=>"000110010",
37019=>"000000000",
37020=>"100111110",
37021=>"001101000",
37022=>"000011111",
37023=>"101100101",
37024=>"100110111",
37025=>"111111111",
37026=>"111000000",
37027=>"111111000",
37028=>"011110001",
37029=>"000000000",
37030=>"000000101",
37031=>"100111011",
37032=>"000110100",
37033=>"000000001",
37034=>"000000000",
37035=>"000000000",
37036=>"000000101",
37037=>"110011001",
37038=>"110111111",
37039=>"011001011",
37040=>"000000000",
37041=>"000110010",
37042=>"111000001",
37043=>"111110000",
37044=>"111111110",
37045=>"110100000",
37046=>"000000000",
37047=>"000000000",
37048=>"000000000",
37049=>"000000000",
37050=>"000000000",
37051=>"000101010",
37052=>"000100010",
37053=>"100101101",
37054=>"001001000",
37055=>"111000011",
37056=>"011011001",
37057=>"000000000",
37058=>"000100010",
37059=>"011111110",
37060=>"000000111",
37061=>"111111111",
37062=>"111000000",
37063=>"101101111",
37064=>"100100100",
37065=>"000000011",
37066=>"000000000",
37067=>"011111010",
37068=>"111000000",
37069=>"000000001",
37070=>"000000000",
37071=>"000001000",
37072=>"010111111",
37073=>"000000100",
37074=>"000000000",
37075=>"111111110",
37076=>"000000000",
37077=>"000100000",
37078=>"010011110",
37079=>"111001001",
37080=>"111111111",
37081=>"011111010",
37082=>"010111011",
37083=>"000000000",
37084=>"111111111",
37085=>"000000000",
37086=>"000000000",
37087=>"111110110",
37088=>"000000111",
37089=>"011010010",
37090=>"110000100",
37091=>"000000000",
37092=>"000000000",
37093=>"010001100",
37094=>"000000001",
37095=>"011011111",
37096=>"000000010",
37097=>"000001000",
37098=>"110110110",
37099=>"000000100",
37100=>"000111111",
37101=>"101111000",
37102=>"000010000",
37103=>"001000100",
37104=>"001000111",
37105=>"111111111",
37106=>"000001000",
37107=>"111111000",
37108=>"111011000",
37109=>"010111111",
37110=>"011000000",
37111=>"000000000",
37112=>"001000000",
37113=>"111000010",
37114=>"000000111",
37115=>"100011101",
37116=>"000000010",
37117=>"011011000",
37118=>"101000011",
37119=>"011011000",
37120=>"100100111",
37121=>"101100001",
37122=>"101001001",
37123=>"111000111",
37124=>"100100110",
37125=>"001101011",
37126=>"111110111",
37127=>"011110011",
37128=>"011011001",
37129=>"001001101",
37130=>"101011111",
37131=>"001001101",
37132=>"111000000",
37133=>"111011001",
37134=>"000000001",
37135=>"111101001",
37136=>"000000000",
37137=>"000000110",
37138=>"000000000",
37139=>"111000000",
37140=>"101101111",
37141=>"101100111",
37142=>"000000000",
37143=>"000010010",
37144=>"101000010",
37145=>"111101111",
37146=>"000100101",
37147=>"000001001",
37148=>"100101010",
37149=>"111110100",
37150=>"000000000",
37151=>"110110010",
37152=>"000000000",
37153=>"000000101",
37154=>"000010010",
37155=>"101000000",
37156=>"111110011",
37157=>"001001111",
37158=>"001000010",
37159=>"000010011",
37160=>"000111111",
37161=>"111111111",
37162=>"111110111",
37163=>"001000011",
37164=>"111100010",
37165=>"010001010",
37166=>"000000011",
37167=>"111111100",
37168=>"111101001",
37169=>"000111111",
37170=>"001110000",
37171=>"101101101",
37172=>"001111111",
37173=>"100111111",
37174=>"001001001",
37175=>"111111011",
37176=>"100001110",
37177=>"111001000",
37178=>"111101000",
37179=>"000111111",
37180=>"111011011",
37181=>"011111111",
37182=>"000000001",
37183=>"000111010",
37184=>"011101000",
37185=>"000101111",
37186=>"001000011",
37187=>"100110100",
37188=>"011000000",
37189=>"000000100",
37190=>"001100110",
37191=>"011111101",
37192=>"111011111",
37193=>"000000001",
37194=>"111000001",
37195=>"111100101",
37196=>"101001111",
37197=>"010011101",
37198=>"110111011",
37199=>"001000111",
37200=>"001001000",
37201=>"111111111",
37202=>"000000000",
37203=>"001101100",
37204=>"100000000",
37205=>"110011011",
37206=>"111011111",
37207=>"100000000",
37208=>"001111111",
37209=>"011001001",
37210=>"011011011",
37211=>"000001100",
37212=>"000000000",
37213=>"110000101",
37214=>"111111000",
37215=>"001110000",
37216=>"000010011",
37217=>"001000011",
37218=>"000000000",
37219=>"101011111",
37220=>"011001010",
37221=>"111100100",
37222=>"010000110",
37223=>"111010110",
37224=>"111100001",
37225=>"000010110",
37226=>"001010111",
37227=>"011011111",
37228=>"010001011",
37229=>"001001001",
37230=>"011111000",
37231=>"101001101",
37232=>"010010011",
37233=>"101000010",
37234=>"100100100",
37235=>"010110110",
37236=>"100111111",
37237=>"000000111",
37238=>"111101111",
37239=>"000001111",
37240=>"000000000",
37241=>"000000000",
37242=>"001000101",
37243=>"111111010",
37244=>"001000001",
37245=>"101000001",
37246=>"101000000",
37247=>"001001101",
37248=>"010001100",
37249=>"010000011",
37250=>"101001110",
37251=>"111101110",
37252=>"111111111",
37253=>"011110100",
37254=>"100100111",
37255=>"010100101",
37256=>"110010110",
37257=>"010001001",
37258=>"000010000",
37259=>"011000000",
37260=>"000000011",
37261=>"111001001",
37262=>"011111100",
37263=>"000001000",
37264=>"111100100",
37265=>"001111111",
37266=>"000001110",
37267=>"111111000",
37268=>"111101000",
37269=>"001000000",
37270=>"110111000",
37271=>"010000101",
37272=>"111010000",
37273=>"000010001",
37274=>"111111111",
37275=>"000010000",
37276=>"111101101",
37277=>"001111100",
37278=>"000010111",
37279=>"011101111",
37280=>"011111110",
37281=>"000000100",
37282=>"011000001",
37283=>"001001111",
37284=>"000000101",
37285=>"101101011",
37286=>"000111110",
37287=>"000000000",
37288=>"101000000",
37289=>"000101000",
37290=>"001001000",
37291=>"000000000",
37292=>"000111111",
37293=>"000100101",
37294=>"100010000",
37295=>"000111000",
37296=>"000100001",
37297=>"010100000",
37298=>"111101111",
37299=>"100000111",
37300=>"111011010",
37301=>"010100000",
37302=>"001000110",
37303=>"111100111",
37304=>"111100110",
37305=>"111001101",
37306=>"101111111",
37307=>"111001101",
37308=>"100110110",
37309=>"000011011",
37310=>"000110000",
37311=>"000101111",
37312=>"000000101",
37313=>"000000010",
37314=>"100000010",
37315=>"011111000",
37316=>"010110010",
37317=>"001001000",
37318=>"110111100",
37319=>"001000100",
37320=>"111011011",
37321=>"111000111",
37322=>"000000101",
37323=>"000111111",
37324=>"110111111",
37325=>"000000100",
37326=>"011101101",
37327=>"101101010",
37328=>"000010000",
37329=>"001110011",
37330=>"111101101",
37331=>"111111000",
37332=>"100010000",
37333=>"011001100",
37334=>"100000000",
37335=>"110101010",
37336=>"010110010",
37337=>"000110000",
37338=>"001101000",
37339=>"000000001",
37340=>"110110010",
37341=>"100000010",
37342=>"110110111",
37343=>"100000000",
37344=>"000000000",
37345=>"000000100",
37346=>"110110110",
37347=>"000000000",
37348=>"101000001",
37349=>"000101111",
37350=>"101001000",
37351=>"111110001",
37352=>"111010110",
37353=>"101000111",
37354=>"110110110",
37355=>"101000101",
37356=>"000000000",
37357=>"000110001",
37358=>"111000110",
37359=>"010111010",
37360=>"111111110",
37361=>"101000110",
37362=>"000000001",
37363=>"111101001",
37364=>"010000110",
37365=>"000000011",
37366=>"101000110",
37367=>"100111111",
37368=>"000000111",
37369=>"110110111",
37370=>"101100111",
37371=>"011001000",
37372=>"111011000",
37373=>"000000100",
37374=>"101111001",
37375=>"000000010",
37376=>"001001100",
37377=>"000001010",
37378=>"110010000",
37379=>"111101101",
37380=>"111011111",
37381=>"001000111",
37382=>"111111010",
37383=>"010001111",
37384=>"101001010",
37385=>"000000000",
37386=>"011110010",
37387=>"000000001",
37388=>"000000101",
37389=>"100000101",
37390=>"000001011",
37391=>"110001101",
37392=>"000101111",
37393=>"100111111",
37394=>"101110000",
37395=>"110111011",
37396=>"111111110",
37397=>"000000000",
37398=>"110110001",
37399=>"001110110",
37400=>"100000101",
37401=>"000000001",
37402=>"000000100",
37403=>"001111111",
37404=>"101101000",
37405=>"011000000",
37406=>"000000101",
37407=>"010000000",
37408=>"111111101",
37409=>"000100111",
37410=>"111111010",
37411=>"000111110",
37412=>"111001011",
37413=>"100001000",
37414=>"110110111",
37415=>"000000000",
37416=>"111010000",
37417=>"101000001",
37418=>"100110111",
37419=>"000000000",
37420=>"111111110",
37421=>"001111000",
37422=>"000110100",
37423=>"110000000",
37424=>"111111001",
37425=>"001111111",
37426=>"111011001",
37427=>"000011010",
37428=>"000111011",
37429=>"000000000",
37430=>"000001111",
37431=>"011000110",
37432=>"110111111",
37433=>"000111010",
37434=>"001000000",
37435=>"100000000",
37436=>"000001001",
37437=>"010010010",
37438=>"000100100",
37439=>"110001100",
37440=>"011010101",
37441=>"101000000",
37442=>"000000110",
37443=>"011011001",
37444=>"111000111",
37445=>"111100000",
37446=>"111000000",
37447=>"111101100",
37448=>"101011011",
37449=>"101101111",
37450=>"101001011",
37451=>"000010111",
37452=>"000000001",
37453=>"101111111",
37454=>"000010111",
37455=>"111100111",
37456=>"000100000",
37457=>"111111010",
37458=>"000111101",
37459=>"011000110",
37460=>"000000111",
37461=>"100100000",
37462=>"111011000",
37463=>"000000111",
37464=>"000000111",
37465=>"001000001",
37466=>"011000001",
37467=>"001111100",
37468=>"111111010",
37469=>"110000001",
37470=>"010111111",
37471=>"110100000",
37472=>"011101111",
37473=>"001000100",
37474=>"001111111",
37475=>"100000000",
37476=>"000000001",
37477=>"000111000",
37478=>"111000000",
37479=>"111101100",
37480=>"010000100",
37481=>"111010000",
37482=>"111011111",
37483=>"111000111",
37484=>"111110110",
37485=>"111111110",
37486=>"111000000",
37487=>"000100010",
37488=>"101110111",
37489=>"111000111",
37490=>"001110111",
37491=>"111111100",
37492=>"111000000",
37493=>"000000101",
37494=>"001000111",
37495=>"000001100",
37496=>"111001000",
37497=>"010000110",
37498=>"111111010",
37499=>"110000000",
37500=>"011101110",
37501=>"110000001",
37502=>"111111000",
37503=>"000001101",
37504=>"100010000",
37505=>"000000000",
37506=>"101011000",
37507=>"011111000",
37508=>"010111111",
37509=>"011010000",
37510=>"001000000",
37511=>"000000000",
37512=>"000101111",
37513=>"000000000",
37514=>"011111101",
37515=>"110111001",
37516=>"000010000",
37517=>"010001000",
37518=>"111000000",
37519=>"000001101",
37520=>"101111011",
37521=>"000000110",
37522=>"101100001",
37523=>"100111111",
37524=>"011111101",
37525=>"100000111",
37526=>"000001000",
37527=>"100000000",
37528=>"010000000",
37529=>"110111111",
37530=>"110110101",
37531=>"011001000",
37532=>"110000110",
37533=>"000000111",
37534=>"000111010",
37535=>"000000000",
37536=>"111001000",
37537=>"000000010",
37538=>"010000001",
37539=>"100000011",
37540=>"111010011",
37541=>"100000000",
37542=>"111010000",
37543=>"000010010",
37544=>"001000111",
37545=>"000110000",
37546=>"000000000",
37547=>"000111111",
37548=>"111011100",
37549=>"001101001",
37550=>"000000001",
37551=>"111011011",
37552=>"010000000",
37553=>"000001010",
37554=>"111000000",
37555=>"101000100",
37556=>"111011110",
37557=>"111111100",
37558=>"010111111",
37559=>"001000000",
37560=>"000101010",
37561=>"100100101",
37562=>"000000111",
37563=>"111000000",
37564=>"001010000",
37565=>"111011111",
37566=>"000100001",
37567=>"101110011",
37568=>"100000010",
37569=>"000111010",
37570=>"101101111",
37571=>"011101100",
37572=>"111110000",
37573=>"100100110",
37574=>"111110110",
37575=>"000000000",
37576=>"111111001",
37577=>"101111101",
37578=>"111111110",
37579=>"111001000",
37580=>"111000100",
37581=>"100101011",
37582=>"000111011",
37583=>"011111110",
37584=>"000111111",
37585=>"000001111",
37586=>"000101111",
37587=>"010000000",
37588=>"000000111",
37589=>"101000010",
37590=>"000000111",
37591=>"110100111",
37592=>"111000000",
37593=>"011111111",
37594=>"010110000",
37595=>"111010000",
37596=>"011111100",
37597=>"110110000",
37598=>"001001100",
37599=>"000100111",
37600=>"101110111",
37601=>"111010011",
37602=>"010000101",
37603=>"000111110",
37604=>"110100101",
37605=>"110100111",
37606=>"000111111",
37607=>"010111100",
37608=>"001001100",
37609=>"110000001",
37610=>"100100100",
37611=>"000100111",
37612=>"000000110",
37613=>"000000001",
37614=>"000000010",
37615=>"111000000",
37616=>"000000001",
37617=>"001011001",
37618=>"010011000",
37619=>"110011011",
37620=>"100111111",
37621=>"010000011",
37622=>"000010111",
37623=>"111011000",
37624=>"001111000",
37625=>"111000000",
37626=>"111001001",
37627=>"000001111",
37628=>"111111000",
37629=>"111111111",
37630=>"000001100",
37631=>"101101110",
37632=>"001110100",
37633=>"100111010",
37634=>"111000101",
37635=>"001111111",
37636=>"000000100",
37637=>"000010000",
37638=>"000101110",
37639=>"010010100",
37640=>"100001111",
37641=>"111100000",
37642=>"011011000",
37643=>"011011001",
37644=>"010011001",
37645=>"000000111",
37646=>"011011000",
37647=>"001000000",
37648=>"000100100",
37649=>"100111010",
37650=>"001000010",
37651=>"000000000",
37652=>"111000011",
37653=>"001000000",
37654=>"101011100",
37655=>"001111110",
37656=>"100101100",
37657=>"001101101",
37658=>"000111111",
37659=>"011011000",
37660=>"101111011",
37661=>"100100000",
37662=>"111111100",
37663=>"000011111",
37664=>"010000110",
37665=>"000100111",
37666=>"111000100",
37667=>"111111001",
37668=>"111001110",
37669=>"010000000",
37670=>"100000000",
37671=>"111011001",
37672=>"011011000",
37673=>"101101111",
37674=>"000110111",
37675=>"000000000",
37676=>"100111110",
37677=>"000111011",
37678=>"011010000",
37679=>"110100001",
37680=>"111111110",
37681=>"011011011",
37682=>"100100111",
37683=>"110111111",
37684=>"011011000",
37685=>"000000000",
37686=>"001001010",
37687=>"000101111",
37688=>"110100001",
37689=>"000000111",
37690=>"000100100",
37691=>"111111010",
37692=>"111111001",
37693=>"111111001",
37694=>"011000000",
37695=>"111111100",
37696=>"000010101",
37697=>"001111111",
37698=>"000110110",
37699=>"111110100",
37700=>"000100101",
37701=>"100001101",
37702=>"010000100",
37703=>"100100111",
37704=>"001001111",
37705=>"011010000",
37706=>"101100101",
37707=>"100101111",
37708=>"100100111",
37709=>"010110110",
37710=>"111111000",
37711=>"000000100",
37712=>"111100000",
37713=>"101100111",
37714=>"000100101",
37715=>"011110000",
37716=>"011011000",
37717=>"101111000",
37718=>"111110000",
37719=>"111010000",
37720=>"110000100",
37721=>"101111001",
37722=>"111100011",
37723=>"011011011",
37724=>"000111101",
37725=>"001001011",
37726=>"101100111",
37727=>"111000100",
37728=>"001111111",
37729=>"111111000",
37730=>"010100100",
37731=>"111011110",
37732=>"000000000",
37733=>"001000011",
37734=>"001011000",
37735=>"000100110",
37736=>"101100000",
37737=>"010111111",
37738=>"000000111",
37739=>"000000101",
37740=>"100000111",
37741=>"110100010",
37742=>"111100110",
37743=>"111011011",
37744=>"110110010",
37745=>"000000000",
37746=>"100111011",
37747=>"110111110",
37748=>"001101000",
37749=>"000100111",
37750=>"111111000",
37751=>"000000001",
37752=>"111110111",
37753=>"000111111",
37754=>"000010010",
37755=>"000000100",
37756=>"110010010",
37757=>"110111100",
37758=>"000000100",
37759=>"111010000",
37760=>"101111010",
37761=>"100011100",
37762=>"100101000",
37763=>"100111111",
37764=>"011001000",
37765=>"110000111",
37766=>"010100101",
37767=>"010010000",
37768=>"111011000",
37769=>"000000000",
37770=>"111110011",
37771=>"000000000",
37772=>"111111000",
37773=>"110000000",
37774=>"011011111",
37775=>"110000010",
37776=>"110110100",
37777=>"000010111",
37778=>"100000000",
37779=>"011111001",
37780=>"011011000",
37781=>"010000101",
37782=>"000111111",
37783=>"100100111",
37784=>"100111011",
37785=>"101011111",
37786=>"000100111",
37787=>"100100101",
37788=>"000000111",
37789=>"000100010",
37790=>"110111111",
37791=>"100000100",
37792=>"100110111",
37793=>"000000000",
37794=>"000000111",
37795=>"100000101",
37796=>"000010001",
37797=>"010110100",
37798=>"100101011",
37799=>"000100111",
37800=>"000111111",
37801=>"110000010",
37802=>"111100000",
37803=>"010100000",
37804=>"100100111",
37805=>"011010000",
37806=>"111101000",
37807=>"010000001",
37808=>"100110101",
37809=>"001110111",
37810=>"100101010",
37811=>"000010100",
37812=>"001001000",
37813=>"101111010",
37814=>"100100100",
37815=>"000000000",
37816=>"111011011",
37817=>"110110100",
37818=>"010101000",
37819=>"100010111",
37820=>"000001101",
37821=>"110100000",
37822=>"101111011",
37823=>"000011100",
37824=>"000100100",
37825=>"000101010",
37826=>"111111111",
37827=>"110110000",
37828=>"011000000",
37829=>"101001011",
37830=>"000010111",
37831=>"011000110",
37832=>"000000100",
37833=>"100101110",
37834=>"000100101",
37835=>"111100000",
37836=>"000000110",
37837=>"011011100",
37838=>"011011011",
37839=>"111111111",
37840=>"100100111",
37841=>"001011110",
37842=>"010000111",
37843=>"100101110",
37844=>"011000000",
37845=>"111001110",
37846=>"100100111",
37847=>"000011110",
37848=>"000000011",
37849=>"100100100",
37850=>"001101101",
37851=>"110000000",
37852=>"110100100",
37853=>"100000011",
37854=>"000111010",
37855=>"111011111",
37856=>"000001111",
37857=>"011011100",
37858=>"011011010",
37859=>"110110000",
37860=>"101110000",
37861=>"100100000",
37862=>"000100101",
37863=>"110110111",
37864=>"111011010",
37865=>"010100111",
37866=>"111110000",
37867=>"111111100",
37868=>"010010000",
37869=>"011010000",
37870=>"010010000",
37871=>"000110011",
37872=>"101001000",
37873=>"001001101",
37874=>"100111100",
37875=>"100100110",
37876=>"100111011",
37877=>"010101110",
37878=>"011100000",
37879=>"110011110",
37880=>"000000100",
37881=>"110100100",
37882=>"000001001",
37883=>"100101010",
37884=>"101011010",
37885=>"011000000",
37886=>"001011000",
37887=>"011000000",
37888=>"010011001",
37889=>"001010000",
37890=>"111100100",
37891=>"011001010",
37892=>"100110110",
37893=>"010000011",
37894=>"000101111",
37895=>"100111110",
37896=>"101000100",
37897=>"000000111",
37898=>"000110010",
37899=>"100010011",
37900=>"111100100",
37901=>"000101011",
37902=>"101111001",
37903=>"001111111",
37904=>"000010010",
37905=>"000011010",
37906=>"011000000",
37907=>"000000011",
37908=>"111100101",
37909=>"001000000",
37910=>"111000000",
37911=>"110010111",
37912=>"010010100",
37913=>"001000111",
37914=>"111100000",
37915=>"000100000",
37916=>"000000000",
37917=>"100101011",
37918=>"000010011",
37919=>"111000011",
37920=>"011101100",
37921=>"111100000",
37922=>"011111100",
37923=>"101101001",
37924=>"010110110",
37925=>"000110100",
37926=>"110100100",
37927=>"001110111",
37928=>"000010100",
37929=>"010011011",
37930=>"000011111",
37931=>"101111110",
37932=>"011111100",
37933=>"111111111",
37934=>"010010111",
37935=>"111111011",
37936=>"111111101",
37937=>"111111111",
37938=>"111000001",
37939=>"111010011",
37940=>"000110111",
37941=>"011011001",
37942=>"000000010",
37943=>"000010000",
37944=>"000000011",
37945=>"001111011",
37946=>"000011010",
37947=>"000111000",
37948=>"000110110",
37949=>"011101110",
37950=>"010000000",
37951=>"110110101",
37952=>"010000000",
37953=>"111111000",
37954=>"111000100",
37955=>"111100111",
37956=>"111101101",
37957=>"000000101",
37958=>"000111101",
37959=>"000010000",
37960=>"110111001",
37961=>"000111011",
37962=>"111001111",
37963=>"000010010",
37964=>"111000001",
37965=>"111011011",
37966=>"010111111",
37967=>"111111000",
37968=>"011001011",
37969=>"011111111",
37970=>"111011000",
37971=>"011001000",
37972=>"000010010",
37973=>"000111011",
37974=>"011011001",
37975=>"000100101",
37976=>"100001011",
37977=>"011111011",
37978=>"101110111",
37979=>"000001111",
37980=>"111000000",
37981=>"101000000",
37982=>"101111011",
37983=>"001001001",
37984=>"111111001",
37985=>"110111011",
37986=>"110100101",
37987=>"010100000",
37988=>"000101111",
37989=>"100111111",
37990=>"111111111",
37991=>"101100101",
37992=>"111011110",
37993=>"000010110",
37994=>"000000000",
37995=>"011010001",
37996=>"111111001",
37997=>"100111111",
37998=>"011101100",
37999=>"100110111",
38000=>"001001101",
38001=>"101111111",
38002=>"000001011",
38003=>"101100100",
38004=>"000101111",
38005=>"000000101",
38006=>"011100111",
38007=>"111111111",
38008=>"010111000",
38009=>"000000100",
38010=>"001000100",
38011=>"111111101",
38012=>"000110010",
38013=>"111100000",
38014=>"111101101",
38015=>"101000111",
38016=>"110000000",
38017=>"010000000",
38018=>"000111010",
38019=>"000000110",
38020=>"100101000",
38021=>"000101000",
38022=>"100011111",
38023=>"100000011",
38024=>"111101111",
38025=>"101011101",
38026=>"000001001",
38027=>"100000111",
38028=>"111100101",
38029=>"000000000",
38030=>"000011111",
38031=>"100001001",
38032=>"011111111",
38033=>"111011011",
38034=>"000011100",
38035=>"000000000",
38036=>"000000000",
38037=>"000000100",
38038=>"000010011",
38039=>"110110100",
38040=>"101000010",
38041=>"111111000",
38042=>"000111011",
38043=>"000000100",
38044=>"101000000",
38045=>"001010010",
38046=>"001100011",
38047=>"111101000",
38048=>"110101011",
38049=>"111011011",
38050=>"010000101",
38051=>"111000000",
38052=>"011110100",
38053=>"100100111",
38054=>"001001001",
38055=>"000000000",
38056=>"000000000",
38057=>"111001000",
38058=>"011101101",
38059=>"000000010",
38060=>"000010000",
38061=>"110000000",
38062=>"011111100",
38063=>"111001000",
38064=>"011011000",
38065=>"001000110",
38066=>"100011111",
38067=>"001000000",
38068=>"000110111",
38069=>"010010111",
38070=>"111111110",
38071=>"001010010",
38072=>"000011111",
38073=>"000000011",
38074=>"000110111",
38075=>"111111010",
38076=>"000000111",
38077=>"110111111",
38078=>"001001000",
38079=>"111000000",
38080=>"000010010",
38081=>"000110111",
38082=>"111110101",
38083=>"001110110",
38084=>"000111101",
38085=>"010110101",
38086=>"111111100",
38087=>"000101100",
38088=>"101110111",
38089=>"111101000",
38090=>"111101000",
38091=>"111111111",
38092=>"000010010",
38093=>"000001010",
38094=>"010010010",
38095=>"111100100",
38096=>"000011111",
38097=>"011111001",
38098=>"101000000",
38099=>"000111011",
38100=>"101000100",
38101=>"100000000",
38102=>"111100000",
38103=>"000111111",
38104=>"010011000",
38105=>"101000000",
38106=>"000001000",
38107=>"111000111",
38108=>"011100100",
38109=>"111100000",
38110=>"000011111",
38111=>"000010110",
38112=>"111100000",
38113=>"011101101",
38114=>"000111111",
38115=>"110100101",
38116=>"101000000",
38117=>"000000000",
38118=>"010000000",
38119=>"110001000",
38120=>"111111100",
38121=>"011111110",
38122=>"000111011",
38123=>"010111101",
38124=>"111100000",
38125=>"101111110",
38126=>"010000000",
38127=>"000000011",
38128=>"000100111",
38129=>"100011001",
38130=>"010000000",
38131=>"110011001",
38132=>"000110011",
38133=>"110111111",
38134=>"000000010",
38135=>"011101100",
38136=>"000111000",
38137=>"111111111",
38138=>"010100101",
38139=>"010001101",
38140=>"000010010",
38141=>"000000000",
38142=>"011000101",
38143=>"111111000",
38144=>"011011100",
38145=>"111110010",
38146=>"000000010",
38147=>"000010111",
38148=>"010001001",
38149=>"000100000",
38150=>"000111111",
38151=>"111111011",
38152=>"000000101",
38153=>"111011111",
38154=>"100100100",
38155=>"100101000",
38156=>"111000000",
38157=>"000000111",
38158=>"100001100",
38159=>"000101010",
38160=>"000111011",
38161=>"000001000",
38162=>"101000010",
38163=>"011010000",
38164=>"000011111",
38165=>"000010010",
38166=>"011011111",
38167=>"000010111",
38168=>"101010010",
38169=>"101111111",
38170=>"000110100",
38171=>"111010110",
38172=>"101101000",
38173=>"110000000",
38174=>"001001010",
38175=>"001001000",
38176=>"000000010",
38177=>"101101110",
38178=>"010000000",
38179=>"111111011",
38180=>"001001000",
38181=>"001101000",
38182=>"010010100",
38183=>"010010101",
38184=>"111101101",
38185=>"010000001",
38186=>"101001111",
38187=>"010000010",
38188=>"110100000",
38189=>"011010000",
38190=>"000000110",
38191=>"110110001",
38192=>"000101111",
38193=>"101101100",
38194=>"100100001",
38195=>"000110111",
38196=>"111000000",
38197=>"011010111",
38198=>"111110010",
38199=>"010000101",
38200=>"111001001",
38201=>"000111000",
38202=>"000000010",
38203=>"001110010",
38204=>"110111010",
38205=>"011101000",
38206=>"000001100",
38207=>"011011011",
38208=>"111011000",
38209=>"001101100",
38210=>"001111001",
38211=>"011001000",
38212=>"000001000",
38213=>"000001000",
38214=>"010110000",
38215=>"010000100",
38216=>"111110001",
38217=>"111111111",
38218=>"000000000",
38219=>"101110111",
38220=>"000010111",
38221=>"100100100",
38222=>"011001001",
38223=>"000000001",
38224=>"111100000",
38225=>"000000111",
38226=>"101101010",
38227=>"001000010",
38228=>"111111101",
38229=>"011111110",
38230=>"100101100",
38231=>"000010000",
38232=>"111111111",
38233=>"011100100",
38234=>"111100000",
38235=>"110101111",
38236=>"000011011",
38237=>"000000010",
38238=>"000011111",
38239=>"110100100",
38240=>"111100000",
38241=>"101000000",
38242=>"000000111",
38243=>"001001100",
38244=>"100100000",
38245=>"111001001",
38246=>"100111000",
38247=>"000001101",
38248=>"111010011",
38249=>"111000111",
38250=>"000000111",
38251=>"000111111",
38252=>"110000000",
38253=>"000000111",
38254=>"100110111",
38255=>"101000100",
38256=>"111101010",
38257=>"000111111",
38258=>"111011010",
38259=>"101000000",
38260=>"100000000",
38261=>"000100100",
38262=>"000011111",
38263=>"000000100",
38264=>"000010111",
38265=>"111011111",
38266=>"100100101",
38267=>"011001101",
38268=>"001001011",
38269=>"110100010",
38270=>"111100001",
38271=>"101101101",
38272=>"010111111",
38273=>"100000000",
38274=>"000000011",
38275=>"000000011",
38276=>"100111010",
38277=>"111101111",
38278=>"100100000",
38279=>"000001001",
38280=>"111100100",
38281=>"000000000",
38282=>"100110011",
38283=>"110010010",
38284=>"010110101",
38285=>"000101100",
38286=>"011101000",
38287=>"100100100",
38288=>"101101100",
38289=>"011111000",
38290=>"101111111",
38291=>"110000101",
38292=>"000001101",
38293=>"000010111",
38294=>"010111011",
38295=>"010011110",
38296=>"111111100",
38297=>"010111111",
38298=>"111101111",
38299=>"001000000",
38300=>"000000000",
38301=>"111111000",
38302=>"111111111",
38303=>"111111100",
38304=>"111001001",
38305=>"111111111",
38306=>"000000000",
38307=>"011101101",
38308=>"001110111",
38309=>"011001000",
38310=>"101000101",
38311=>"011111100",
38312=>"100000111",
38313=>"011000000",
38314=>"101101111",
38315=>"101010010",
38316=>"111000010",
38317=>"111001100",
38318=>"110100000",
38319=>"111111101",
38320=>"111110000",
38321=>"001101100",
38322=>"010000111",
38323=>"011000000",
38324=>"011111110",
38325=>"100100000",
38326=>"111011111",
38327=>"101110010",
38328=>"001011010",
38329=>"000000111",
38330=>"011010000",
38331=>"100100111",
38332=>"111100000",
38333=>"100111111",
38334=>"010010110",
38335=>"111000000",
38336=>"101111111",
38337=>"000010010",
38338=>"000110010",
38339=>"011001000",
38340=>"000011111",
38341=>"011001001",
38342=>"111011011",
38343=>"000000110",
38344=>"000111111",
38345=>"010010110",
38346=>"010011011",
38347=>"100100000",
38348=>"001100000",
38349=>"000100110",
38350=>"101000000",
38351=>"010010000",
38352=>"001000000",
38353=>"111101001",
38354=>"000000101",
38355=>"001000000",
38356=>"110101101",
38357=>"110100000",
38358=>"000010010",
38359=>"010011010",
38360=>"011111000",
38361=>"010000000",
38362=>"110101100",
38363=>"100000110",
38364=>"111110111",
38365=>"111111111",
38366=>"111111101",
38367=>"000000001",
38368=>"000000111",
38369=>"000000111",
38370=>"111111001",
38371=>"001001001",
38372=>"000010110",
38373=>"010100000",
38374=>"101000000",
38375=>"111011001",
38376=>"110000000",
38377=>"111001010",
38378=>"001001000",
38379=>"101110111",
38380=>"000000000",
38381=>"000111111",
38382=>"000000000",
38383=>"100010000",
38384=>"111000000",
38385=>"000100000",
38386=>"001000111",
38387=>"111001011",
38388=>"110110000",
38389=>"101000000",
38390=>"000000010",
38391=>"101111101",
38392=>"000110101",
38393=>"000001010",
38394=>"111001110",
38395=>"010000100",
38396=>"010000000",
38397=>"000111111",
38398=>"110100000",
38399=>"010010000",
38400=>"001000100",
38401=>"000011000",
38402=>"000000101",
38403=>"101110100",
38404=>"111111011",
38405=>"001000011",
38406=>"000000110",
38407=>"000101000",
38408=>"111111010",
38409=>"111110100",
38410=>"111110111",
38411=>"000000100",
38412=>"000000000",
38413=>"101111111",
38414=>"011011000",
38415=>"001001101",
38416=>"111101011",
38417=>"110000000",
38418=>"000000000",
38419=>"010000001",
38420=>"111111010",
38421=>"111110000",
38422=>"111001000",
38423=>"000111000",
38424=>"000000111",
38425=>"000000000",
38426=>"100100000",
38427=>"110111111",
38428=>"100000000",
38429=>"000000101",
38430=>"000000111",
38431=>"010000001",
38432=>"000000010",
38433=>"111111010",
38434=>"111101010",
38435=>"011111111",
38436=>"010110111",
38437=>"011011011",
38438=>"110000000",
38439=>"111111001",
38440=>"110111100",
38441=>"111111111",
38442=>"100000001",
38443=>"101111111",
38444=>"000000001",
38445=>"111100000",
38446=>"000100100",
38447=>"101111010",
38448=>"000111000",
38449=>"000100100",
38450=>"000111110",
38451=>"010110100",
38452=>"010000000",
38453=>"000000000",
38454=>"111111000",
38455=>"000000101",
38456=>"111111111",
38457=>"000000000",
38458=>"000000111",
38459=>"110000010",
38460=>"000000000",
38461=>"111111011",
38462=>"100001111",
38463=>"111111100",
38464=>"001111111",
38465=>"000011000",
38466=>"000100000",
38467=>"011111011",
38468=>"111001111",
38469=>"000000000",
38470=>"111111110",
38471=>"111111111",
38472=>"110110010",
38473=>"000000001",
38474=>"000000000",
38475=>"101100000",
38476=>"000000011",
38477=>"111111110",
38478=>"000011001",
38479=>"000000000",
38480=>"111111000",
38481=>"111111111",
38482=>"111011111",
38483=>"001100111",
38484=>"000000000",
38485=>"111110000",
38486=>"111011000",
38487=>"001000011",
38488=>"011100000",
38489=>"000100100",
38490=>"011011000",
38491=>"111111111",
38492=>"010111111",
38493=>"011001100",
38494=>"111111000",
38495=>"111110110",
38496=>"111111111",
38497=>"111111100",
38498=>"101000111",
38499=>"100000001",
38500=>"101101000",
38501=>"010000101",
38502=>"000000111",
38503=>"111001111",
38504=>"101010101",
38505=>"111111111",
38506=>"100000010",
38507=>"001111000",
38508=>"111111111",
38509=>"110000110",
38510=>"101101111",
38511=>"000000111",
38512=>"011001011",
38513=>"111111111",
38514=>"111111000",
38515=>"111000001",
38516=>"000000110",
38517=>"000001111",
38518=>"101000111",
38519=>"111111111",
38520=>"000000101",
38521=>"111001101",
38522=>"101100001",
38523=>"111111000",
38524=>"111010100",
38525=>"100001110",
38526=>"110111111",
38527=>"001001001",
38528=>"000111111",
38529=>"000000101",
38530=>"111111111",
38531=>"101101111",
38532=>"000000000",
38533=>"111111010",
38534=>"100110000",
38535=>"110110110",
38536=>"110110000",
38537=>"110111100",
38538=>"111111110",
38539=>"001110001",
38540=>"000000010",
38541=>"000101000",
38542=>"001001000",
38543=>"011110000",
38544=>"001001111",
38545=>"101111111",
38546=>"000000000",
38547=>"000000000",
38548=>"111011000",
38549=>"010110000",
38550=>"111111111",
38551=>"001011011",
38552=>"000000000",
38553=>"011010001",
38554=>"101111011",
38555=>"000000000",
38556=>"101110011",
38557=>"010111111",
38558=>"111111000",
38559=>"000000000",
38560=>"001101011",
38561=>"000000111",
38562=>"000101011",
38563=>"000010000",
38564=>"111111011",
38565=>"001011011",
38566=>"110100000",
38567=>"001001111",
38568=>"111001010",
38569=>"111111111",
38570=>"111111110",
38571=>"000001000",
38572=>"101101110",
38573=>"000000111",
38574=>"100100111",
38575=>"111111110",
38576=>"000000100",
38577=>"011010011",
38578=>"000000000",
38579=>"100010001",
38580=>"001000000",
38581=>"111111111",
38582=>"000000111",
38583=>"100000000",
38584=>"100000100",
38585=>"011101000",
38586=>"001111111",
38587=>"001000000",
38588=>"000000000",
38589=>"000000000",
38590=>"110110010",
38591=>"010000101",
38592=>"000010000",
38593=>"000000000",
38594=>"011111110",
38595=>"000000000",
38596=>"000000111",
38597=>"111001000",
38598=>"000001111",
38599=>"111110000",
38600=>"000101001",
38601=>"000000000",
38602=>"100110111",
38603=>"000000010",
38604=>"000000000",
38605=>"111100000",
38606=>"000100101",
38607=>"111111000",
38608=>"110011010",
38609=>"110111111",
38610=>"000000001",
38611=>"000000000",
38612=>"000000100",
38613=>"100000000",
38614=>"111111111",
38615=>"001111111",
38616=>"000000001",
38617=>"111000000",
38618=>"000001110",
38619=>"000000111",
38620=>"111110010",
38621=>"111111000",
38622=>"000001101",
38623=>"111111000",
38624=>"010010001",
38625=>"100110000",
38626=>"010000000",
38627=>"111111000",
38628=>"001000001",
38629=>"100111111",
38630=>"101101010",
38631=>"000010010",
38632=>"001000101",
38633=>"100101000",
38634=>"111111110",
38635=>"001111100",
38636=>"010010000",
38637=>"000000101",
38638=>"111111000",
38639=>"111101000",
38640=>"000000001",
38641=>"111000100",
38642=>"111111110",
38643=>"000001000",
38644=>"001011011",
38645=>"111110000",
38646=>"100101111",
38647=>"000000000",
38648=>"000111111",
38649=>"000100000",
38650=>"110000000",
38651=>"110000000",
38652=>"000001000",
38653=>"000000011",
38654=>"111111110",
38655=>"000000100",
38656=>"000000100",
38657=>"000011111",
38658=>"000000110",
38659=>"111111011",
38660=>"100001001",
38661=>"111100111",
38662=>"101101111",
38663=>"000111111",
38664=>"001001001",
38665=>"000001010",
38666=>"100100000",
38667=>"110110111",
38668=>"111110010",
38669=>"000000001",
38670=>"000010000",
38671=>"000100110",
38672=>"000110111",
38673=>"100011100",
38674=>"111101011",
38675=>"010000001",
38676=>"000000110",
38677=>"000101111",
38678=>"000000000",
38679=>"111111111",
38680=>"111010010",
38681=>"010000101",
38682=>"111001000",
38683=>"100111000",
38684=>"100111110",
38685=>"101100000",
38686=>"000000111",
38687=>"000000000",
38688=>"000010010",
38689=>"000001111",
38690=>"111000110",
38691=>"001111111",
38692=>"010000110",
38693=>"001000000",
38694=>"011111111",
38695=>"101000111",
38696=>"001001000",
38697=>"000111111",
38698=>"000000000",
38699=>"110111110",
38700=>"000011000",
38701=>"100111001",
38702=>"111110111",
38703=>"000000011",
38704=>"000000000",
38705=>"000000000",
38706=>"000000110",
38707=>"000000011",
38708=>"011000001",
38709=>"010111111",
38710=>"011011000",
38711=>"000000001",
38712=>"111100010",
38713=>"000101000",
38714=>"010010010",
38715=>"111010001",
38716=>"010000000",
38717=>"111000111",
38718=>"010000001",
38719=>"011001000",
38720=>"111110111",
38721=>"001111010",
38722=>"000001010",
38723=>"111011000",
38724=>"000000001",
38725=>"000000000",
38726=>"010011011",
38727=>"101100111",
38728=>"001110110",
38729=>"010101011",
38730=>"000000000",
38731=>"001001101",
38732=>"110111100",
38733=>"100100100",
38734=>"001001001",
38735=>"011001011",
38736=>"000001001",
38737=>"111111111",
38738=>"111111111",
38739=>"000010011",
38740=>"001001101",
38741=>"011000000",
38742=>"010001000",
38743=>"000000111",
38744=>"010001001",
38745=>"110110011",
38746=>"000100100",
38747=>"111010110",
38748=>"101001001",
38749=>"000000100",
38750=>"111111111",
38751=>"000000010",
38752=>"010111001",
38753=>"000001000",
38754=>"111110000",
38755=>"110111111",
38756=>"010001000",
38757=>"110000000",
38758=>"000001100",
38759=>"101111111",
38760=>"000000000",
38761=>"000000111",
38762=>"000000000",
38763=>"001101111",
38764=>"000000000",
38765=>"000001111",
38766=>"011001001",
38767=>"000000010",
38768=>"111011000",
38769=>"000010010",
38770=>"110100000",
38771=>"000110011",
38772=>"111110000",
38773=>"010010000",
38774=>"000000001",
38775=>"001010000",
38776=>"111111100",
38777=>"110111111",
38778=>"000000000",
38779=>"111111111",
38780=>"000001000",
38781=>"000010010",
38782=>"111010110",
38783=>"111111010",
38784=>"000000000",
38785=>"000110000",
38786=>"000101011",
38787=>"001101111",
38788=>"111111111",
38789=>"000000000",
38790=>"000000000",
38791=>"000000000",
38792=>"111110000",
38793=>"000000000",
38794=>"000111111",
38795=>"000101111",
38796=>"000000010",
38797=>"111111111",
38798=>"111111111",
38799=>"011010011",
38800=>"110100000",
38801=>"111101000",
38802=>"011001110",
38803=>"000000000",
38804=>"110101100",
38805=>"110010010",
38806=>"111111111",
38807=>"110010101",
38808=>"111111101",
38809=>"000000101",
38810=>"111000000",
38811=>"111010010",
38812=>"110110000",
38813=>"100101111",
38814=>"010100010",
38815=>"000000000",
38816=>"110110011",
38817=>"011000111",
38818=>"011000000",
38819=>"000001111",
38820=>"000110110",
38821=>"110110110",
38822=>"011001011",
38823=>"101001101",
38824=>"000000001",
38825=>"111101111",
38826=>"111000000",
38827=>"001001101",
38828=>"111000000",
38829=>"000000110",
38830=>"111111111",
38831=>"100110111",
38832=>"111000010",
38833=>"000100010",
38834=>"010010000",
38835=>"010010000",
38836=>"111010100",
38837=>"101000011",
38838=>"000010001",
38839=>"001101110",
38840=>"100000000",
38841=>"110000000",
38842=>"010101100",
38843=>"000001000",
38844=>"010000010",
38845=>"110000000",
38846=>"100100100",
38847=>"000010000",
38848=>"001001011",
38849=>"000000000",
38850=>"001011111",
38851=>"101110110",
38852=>"000000000",
38853=>"111011111",
38854=>"000000101",
38855=>"111111010",
38856=>"111101101",
38857=>"111010000",
38858=>"011001110",
38859=>"000001001",
38860=>"110111111",
38861=>"010000001",
38862=>"111111110",
38863=>"111111110",
38864=>"111000111",
38865=>"111111110",
38866=>"000000001",
38867=>"000000010",
38868=>"111111001",
38869=>"000000001",
38870=>"111101101",
38871=>"100000000",
38872=>"001001000",
38873=>"000000010",
38874=>"111011111",
38875=>"000111111",
38876=>"000111010",
38877=>"000000111",
38878=>"000000101",
38879=>"110111100",
38880=>"111001101",
38881=>"101001111",
38882=>"110110110",
38883=>"001000001",
38884=>"111001110",
38885=>"000000111",
38886=>"110100001",
38887=>"000101101",
38888=>"111000100",
38889=>"000111000",
38890=>"011001000",
38891=>"111111111",
38892=>"000001001",
38893=>"110111100",
38894=>"110010010",
38895=>"000010000",
38896=>"000000000",
38897=>"100100011",
38898=>"111110111",
38899=>"110111101",
38900=>"011111111",
38901=>"000101111",
38902=>"110101000",
38903=>"111111111",
38904=>"110111000",
38905=>"000111111",
38906=>"111101101",
38907=>"001000000",
38908=>"111111110",
38909=>"111011111",
38910=>"001011000",
38911=>"111111011",
38912=>"011011001",
38913=>"000100111",
38914=>"101101001",
38915=>"000010111",
38916=>"100000110",
38917=>"111110000",
38918=>"001000000",
38919=>"101101111",
38920=>"111111111",
38921=>"111111001",
38922=>"001100000",
38923=>"011111111",
38924=>"000010011",
38925=>"000000001",
38926=>"100100101",
38927=>"000110000",
38928=>"000001111",
38929=>"000111100",
38930=>"110011010",
38931=>"111111111",
38932=>"111000000",
38933=>"000000011",
38934=>"100000100",
38935=>"010010010",
38936=>"000000011",
38937=>"001010011",
38938=>"111111101",
38939=>"110000000",
38940=>"111111000",
38941=>"000000101",
38942=>"110110000",
38943=>"000000100",
38944=>"111111000",
38945=>"111011001",
38946=>"111000000",
38947=>"000011111",
38948=>"011011001",
38949=>"111110101",
38950=>"111101000",
38951=>"000010000",
38952=>"000000000",
38953=>"001111111",
38954=>"011111101",
38955=>"011000000",
38956=>"001011011",
38957=>"000000010",
38958=>"111011111",
38959=>"000111001",
38960=>"000010010",
38961=>"001111111",
38962=>"111111011",
38963=>"000001000",
38964=>"111000000",
38965=>"000010011",
38966=>"101001000",
38967=>"000010010",
38968=>"000000001",
38969=>"000000000",
38970=>"001010111",
38971=>"000100111",
38972=>"000110110",
38973=>"011001010",
38974=>"000000100",
38975=>"011011001",
38976=>"101111011",
38977=>"111111000",
38978=>"011111111",
38979=>"101001011",
38980=>"010010000",
38981=>"100110011",
38982=>"111111011",
38983=>"111000110",
38984=>"000000100",
38985=>"010010011",
38986=>"000000111",
38987=>"110100010",
38988=>"001111111",
38989=>"110100111",
38990=>"000111011",
38991=>"000111110",
38992=>"010000101",
38993=>"000000000",
38994=>"010111101",
38995=>"011011001",
38996=>"101111111",
38997=>"000000001",
38998=>"011111001",
38999=>"111111101",
39000=>"000001000",
39001=>"100111111",
39002=>"010111110",
39003=>"111010111",
39004=>"111111001",
39005=>"001011000",
39006=>"101000110",
39007=>"110111111",
39008=>"110111111",
39009=>"110110000",
39010=>"111101100",
39011=>"100100101",
39012=>"010110010",
39013=>"101111100",
39014=>"111111101",
39015=>"000010001",
39016=>"111010010",
39017=>"111111010",
39018=>"101111111",
39019=>"000010000",
39020=>"000010000",
39021=>"000100100",
39022=>"000010010",
39023=>"101111100",
39024=>"111110010",
39025=>"000000010",
39026=>"101000100",
39027=>"101111011",
39028=>"111011011",
39029=>"101000101",
39030=>"000001111",
39031=>"111111111",
39032=>"110111101",
39033=>"011110000",
39034=>"010010000",
39035=>"000000000",
39036=>"100110110",
39037=>"110110100",
39038=>"000000000",
39039=>"111000100",
39040=>"010110101",
39041=>"111111000",
39042=>"111111111",
39043=>"000000100",
39044=>"000111111",
39045=>"000000111",
39046=>"111111001",
39047=>"100101111",
39048=>"011111100",
39049=>"111100010",
39050=>"011111110",
39051=>"010011000",
39052=>"110010100",
39053=>"100111111",
39054=>"111111000",
39055=>"111001001",
39056=>"010111011",
39057=>"100000000",
39058=>"010010111",
39059=>"111000011",
39060=>"001011111",
39061=>"101111111",
39062=>"010011000",
39063=>"001011011",
39064=>"100111111",
39065=>"100111111",
39066=>"111000101",
39067=>"011111101",
39068=>"100101100",
39069=>"010011000",
39070=>"111111101",
39071=>"000000000",
39072=>"101001000",
39073=>"000101000",
39074=>"000000000",
39075=>"001011100",
39076=>"111111110",
39077=>"001000110",
39078=>"111110110",
39079=>"010010000",
39080=>"000000101",
39081=>"000011111",
39082=>"000111111",
39083=>"111100000",
39084=>"111011110",
39085=>"111111111",
39086=>"111100000",
39087=>"101101111",
39088=>"111000111",
39089=>"001101001",
39090=>"111111111",
39091=>"101010000",
39092=>"000000100",
39093=>"000110011",
39094=>"111011001",
39095=>"010010111",
39096=>"010111011",
39097=>"000100111",
39098=>"111111100",
39099=>"000110111",
39100=>"010011001",
39101=>"011111111",
39102=>"111111111",
39103=>"001000000",
39104=>"111001111",
39105=>"110111111",
39106=>"011101101",
39107=>"000010011",
39108=>"101000000",
39109=>"000000001",
39110=>"000011010",
39111=>"111100111",
39112=>"000111111",
39113=>"010000111",
39114=>"111000000",
39115=>"000000011",
39116=>"100000100",
39117=>"000011011",
39118=>"111010110",
39119=>"000111011",
39120=>"010000010",
39121=>"101110011",
39122=>"111011111",
39123=>"111111011",
39124=>"001000101",
39125=>"110000110",
39126=>"000000100",
39127=>"000011111",
39128=>"100101101",
39129=>"010000000",
39130=>"010100000",
39131=>"000111000",
39132=>"001001101",
39133=>"010111111",
39134=>"011101111",
39135=>"000000111",
39136=>"000000110",
39137=>"111000100",
39138=>"000000111",
39139=>"001111000",
39140=>"111111100",
39141=>"000011010",
39142=>"111111111",
39143=>"000001000",
39144=>"110010010",
39145=>"101000101",
39146=>"100000000",
39147=>"011010010",
39148=>"000000101",
39149=>"011111111",
39150=>"010010010",
39151=>"010110000",
39152=>"010111100",
39153=>"000000000",
39154=>"011011111",
39155=>"000111011",
39156=>"110110100",
39157=>"111010010",
39158=>"000000000",
39159=>"000000011",
39160=>"001000111",
39161=>"111100110",
39162=>"000010101",
39163=>"100100111",
39164=>"000000000",
39165=>"000000000",
39166=>"000111101",
39167=>"110110111",
39168=>"011011001",
39169=>"110100110",
39170=>"111000100",
39171=>"011000000",
39172=>"000000110",
39173=>"101101000",
39174=>"010110000",
39175=>"000101101",
39176=>"000000000",
39177=>"100000000",
39178=>"001001101",
39179=>"111111010",
39180=>"111101101",
39181=>"110111001",
39182=>"010101011",
39183=>"011110000",
39184=>"000000010",
39185=>"000000000",
39186=>"010111000",
39187=>"000000111",
39188=>"000000100",
39189=>"111100100",
39190=>"100010011",
39191=>"111000000",
39192=>"000000000",
39193=>"000110110",
39194=>"010111000",
39195=>"111000111",
39196=>"110010111",
39197=>"111000000",
39198=>"110010000",
39199=>"111111011",
39200=>"001000000",
39201=>"001010010",
39202=>"001001000",
39203=>"101101000",
39204=>"110110110",
39205=>"000100100",
39206=>"101000111",
39207=>"000010010",
39208=>"010010000",
39209=>"000011011",
39210=>"000001000",
39211=>"000110111",
39212=>"100111101",
39213=>"111111110",
39214=>"010001101",
39215=>"000110000",
39216=>"101000001",
39217=>"110000110",
39218=>"000000000",
39219=>"000111111",
39220=>"100000100",
39221=>"000000000",
39222=>"110111111",
39223=>"111111101",
39224=>"010111010",
39225=>"111011011",
39226=>"000000000",
39227=>"000010000",
39228=>"110100100",
39229=>"001010001",
39230=>"010101001",
39231=>"001001101",
39232=>"000011111",
39233=>"101000000",
39234=>"111111000",
39235=>"101001001",
39236=>"110000000",
39237=>"001000000",
39238=>"010111111",
39239=>"010110000",
39240=>"011101001",
39241=>"111101000",
39242=>"111000000",
39243=>"001001000",
39244=>"000000000",
39245=>"110110111",
39246=>"001001111",
39247=>"100000000",
39248=>"001010010",
39249=>"111111111",
39250=>"000011010",
39251=>"010010000",
39252=>"000000000",
39253=>"101101111",
39254=>"000001010",
39255=>"111000111",
39256=>"010000100",
39257=>"011010111",
39258=>"000101111",
39259=>"001011000",
39260=>"000010000",
39261=>"001001000",
39262=>"111111101",
39263=>"100000110",
39264=>"000010000",
39265=>"010000001",
39266=>"111101000",
39267=>"000000100",
39268=>"011101010",
39269=>"000011000",
39270=>"000000101",
39271=>"011000000",
39272=>"000010110",
39273=>"111011001",
39274=>"000010011",
39275=>"111101100",
39276=>"010010001",
39277=>"111000110",
39278=>"111101000",
39279=>"101000100",
39280=>"000111101",
39281=>"010000000",
39282=>"001011011",
39283=>"000000000",
39284=>"100010111",
39285=>"101100010",
39286=>"011111110",
39287=>"101000000",
39288=>"000000001",
39289=>"110011010",
39290=>"111111111",
39291=>"011101101",
39292=>"000100100",
39293=>"000010000",
39294=>"110000001",
39295=>"000001001",
39296=>"010110000",
39297=>"010101100",
39298=>"111010000",
39299=>"000001101",
39300=>"111100000",
39301=>"110110000",
39302=>"010011001",
39303=>"000001011",
39304=>"000111000",
39305=>"111011000",
39306=>"111000111",
39307=>"101001010",
39308=>"111000000",
39309=>"000111111",
39310=>"111111000",
39311=>"000000000",
39312=>"111101011",
39313=>"010000111",
39314=>"000010000",
39315=>"101000000",
39316=>"000000111",
39317=>"000000010",
39318=>"101001000",
39319=>"100100110",
39320=>"110010100",
39321=>"011000000",
39322=>"110111000",
39323=>"100100100",
39324=>"010100000",
39325=>"001000000",
39326=>"010010010",
39327=>"111000010",
39328=>"110101111",
39329=>"000000110",
39330=>"110101111",
39331=>"000100001",
39332=>"110110110",
39333=>"100110110",
39334=>"000000110",
39335=>"000110000",
39336=>"010110011",
39337=>"011111110",
39338=>"101110110",
39339=>"000000000",
39340=>"000001101",
39341=>"110000010",
39342=>"001110100",
39343=>"110011000",
39344=>"100101101",
39345=>"100101101",
39346=>"111101000",
39347=>"011000000",
39348=>"001011110",
39349=>"010011000",
39350=>"000011011",
39351=>"010011001",
39352=>"011001001",
39353=>"000100110",
39354=>"110110010",
39355=>"111111000",
39356=>"010010000",
39357=>"111111111",
39358=>"001000100",
39359=>"110000011",
39360=>"000000000",
39361=>"010000001",
39362=>"111101001",
39363=>"001010110",
39364=>"011000000",
39365=>"110101111",
39366=>"110110110",
39367=>"001000001",
39368=>"000000101",
39369=>"101000000",
39370=>"010110000",
39371=>"101001111",
39372=>"000000001",
39373=>"100011001",
39374=>"000000000",
39375=>"001111101",
39376=>"111000000",
39377=>"010111011",
39378=>"000100011",
39379=>"111000000",
39380=>"101000000",
39381=>"111111001",
39382=>"110101000",
39383=>"110010000",
39384=>"000000000",
39385=>"101000000",
39386=>"111001111",
39387=>"011001111",
39388=>"001100010",
39389=>"001111000",
39390=>"010110000",
39391=>"100110011",
39392=>"111000101",
39393=>"101101100",
39394=>"111111111",
39395=>"001001000",
39396=>"111000010",
39397=>"011011010",
39398=>"000111111",
39399=>"010000011",
39400=>"100101000",
39401=>"000000101",
39402=>"110000001",
39403=>"001111111",
39404=>"101001000",
39405=>"000000011",
39406=>"010000000",
39407=>"000001010",
39408=>"111001000",
39409=>"011001100",
39410=>"101101101",
39411=>"010110001",
39412=>"010110111",
39413=>"011000011",
39414=>"010000000",
39415=>"000010110",
39416=>"010010011",
39417=>"111000000",
39418=>"010010011",
39419=>"001011000",
39420=>"111100101",
39421=>"111111111",
39422=>"000011011",
39423=>"010001111",
39424=>"011001000",
39425=>"000000100",
39426=>"101001101",
39427=>"011101001",
39428=>"011011010",
39429=>"100000001",
39430=>"010000000",
39431=>"000011010",
39432=>"000100010",
39433=>"111101111",
39434=>"101001011",
39435=>"011011000",
39436=>"010000000",
39437=>"100000101",
39438=>"000011001",
39439=>"010110111",
39440=>"000110010",
39441=>"111101000",
39442=>"000001001",
39443=>"000010000",
39444=>"000111101",
39445=>"110000000",
39446=>"001100101",
39447=>"101101111",
39448=>"101000011",
39449=>"111010110",
39450=>"000000000",
39451=>"101101000",
39452=>"000000000",
39453=>"000001111",
39454=>"111000000",
39455=>"111111101",
39456=>"000110111",
39457=>"010011111",
39458=>"000011000",
39459=>"000011010",
39460=>"000001011",
39461=>"000000000",
39462=>"011110000",
39463=>"011000100",
39464=>"000000001",
39465=>"111110111",
39466=>"001011000",
39467=>"111011000",
39468=>"000000001",
39469=>"100000011",
39470=>"011111111",
39471=>"111101110",
39472=>"000010111",
39473=>"001011110",
39474=>"000000010",
39475=>"000110111",
39476=>"010010000",
39477=>"010110100",
39478=>"100001001",
39479=>"000000110",
39480=>"100111111",
39481=>"000000100",
39482=>"000000000",
39483=>"101100100",
39484=>"110110100",
39485=>"010111001",
39486=>"000000000",
39487=>"111011111",
39488=>"111011111",
39489=>"010010110",
39490=>"000000111",
39491=>"001000000",
39492=>"010111101",
39493=>"010010000",
39494=>"000000111",
39495=>"010010111",
39496=>"011001100",
39497=>"010000000",
39498=>"000000001",
39499=>"111101001",
39500=>"111111110",
39501=>"001110110",
39502=>"100110010",
39503=>"100101001",
39504=>"100000100",
39505=>"000000010",
39506=>"000100111",
39507=>"011000000",
39508=>"001000001",
39509=>"111100100",
39510=>"001001011",
39511=>"000110000",
39512=>"111111000",
39513=>"000000111",
39514=>"111111000",
39515=>"000100000",
39516=>"111011010",
39517=>"000000000",
39518=>"000000110",
39519=>"000001000",
39520=>"110111111",
39521=>"010111101",
39522=>"010001100",
39523=>"111011001",
39524=>"000000000",
39525=>"000100111",
39526=>"111010111",
39527=>"000010111",
39528=>"000001111",
39529=>"000000111",
39530=>"000000000",
39531=>"011010011",
39532=>"100111111",
39533=>"101101111",
39534=>"000000000",
39535=>"000000110",
39536=>"001001010",
39537=>"000000010",
39538=>"001100010",
39539=>"111111111",
39540=>"000000000",
39541=>"000100000",
39542=>"010010011",
39543=>"111101000",
39544=>"111000000",
39545=>"111111000",
39546=>"000000100",
39547=>"000001001",
39548=>"100111011",
39549=>"110000100",
39550=>"010001001",
39551=>"100011000",
39552=>"000000000",
39553=>"000010010",
39554=>"110000100",
39555=>"010100000",
39556=>"001000110",
39557=>"000000000",
39558=>"011000000",
39559=>"000111000",
39560=>"110110110",
39561=>"101010011",
39562=>"111101111",
39563=>"111011001",
39564=>"111000111",
39565=>"011111101",
39566=>"100111010",
39567=>"001001110",
39568=>"100111011",
39569=>"101010000",
39570=>"111000010",
39571=>"011101111",
39572=>"000011011",
39573=>"010110111",
39574=>"000111111",
39575=>"000011001",
39576=>"000000101",
39577=>"000000000",
39578=>"000000111",
39579=>"000101111",
39580=>"110010100",
39581=>"000000010",
39582=>"000000110",
39583=>"111111000",
39584=>"111100000",
39585=>"111000000",
39586=>"010111101",
39587=>"000110101",
39588=>"111000000",
39589=>"110010000",
39590=>"000110000",
39591=>"000000010",
39592=>"000000010",
39593=>"000010111",
39594=>"111111100",
39595=>"111000000",
39596=>"111111000",
39597=>"100110110",
39598=>"111101111",
39599=>"101101110",
39600=>"000001000",
39601=>"100000101",
39602=>"000000000",
39603=>"000000000",
39604=>"111000100",
39605=>"001011111",
39606=>"011011111",
39607=>"011011001",
39608=>"011110000",
39609=>"000110111",
39610=>"110000001",
39611=>"111011000",
39612=>"011001101",
39613=>"000100111",
39614=>"011010010",
39615=>"011001000",
39616=>"100000000",
39617=>"101000000",
39618=>"001001101",
39619=>"111110111",
39620=>"000111000",
39621=>"101011111",
39622=>"000010010",
39623=>"100000101",
39624=>"000111111",
39625=>"110000000",
39626=>"011011111",
39627=>"000001111",
39628=>"000000000",
39629=>"001011110",
39630=>"111110110",
39631=>"110111111",
39632=>"111101000",
39633=>"110110110",
39634=>"100010111",
39635=>"111011111",
39636=>"000000011",
39637=>"001100100",
39638=>"010011111",
39639=>"000011110",
39640=>"111101101",
39641=>"000000111",
39642=>"111011001",
39643=>"000001101",
39644=>"111100101",
39645=>"000111011",
39646=>"111010000",
39647=>"000001101",
39648=>"101000100",
39649=>"011001101",
39650=>"111111101",
39651=>"101111110",
39652=>"101000011",
39653=>"110110000",
39654=>"111011111",
39655=>"011111111",
39656=>"001000000",
39657=>"010000100",
39658=>"100100111",
39659=>"110111111",
39660=>"111110000",
39661=>"111010000",
39662=>"000000000",
39663=>"011111100",
39664=>"111111100",
39665=>"111111101",
39666=>"011010000",
39667=>"000001001",
39668=>"110110000",
39669=>"110100111",
39670=>"000000000",
39671=>"000000000",
39672=>"010000000",
39673=>"000000001",
39674=>"111100000",
39675=>"100111111",
39676=>"000000011",
39677=>"000010111",
39678=>"100011001",
39679=>"000000101",
39680=>"111111111",
39681=>"010000101",
39682=>"000000000",
39683=>"000001111",
39684=>"000111111",
39685=>"001001000",
39686=>"000101101",
39687=>"101001111",
39688=>"111001010",
39689=>"001001111",
39690=>"001000000",
39691=>"001000111",
39692=>"000000000",
39693=>"011001001",
39694=>"111101101",
39695=>"111011111",
39696=>"110000111",
39697=>"000000000",
39698=>"110000100",
39699=>"000000000",
39700=>"111111111",
39701=>"010000110",
39702=>"001011001",
39703=>"101010000",
39704=>"000000000",
39705=>"111111111",
39706=>"111011011",
39707=>"111111000",
39708=>"000000000",
39709=>"111001001",
39710=>"001011111",
39711=>"001000000",
39712=>"111111110",
39713=>"101111111",
39714=>"000000000",
39715=>"000011011",
39716=>"000100000",
39717=>"011011011",
39718=>"001011110",
39719=>"000001000",
39720=>"111111010",
39721=>"011111111",
39722=>"000000011",
39723=>"100000111",
39724=>"010111100",
39725=>"111111100",
39726=>"000001000",
39727=>"010111011",
39728=>"101111000",
39729=>"100100001",
39730=>"001010001",
39731=>"010111101",
39732=>"000000000",
39733=>"101111111",
39734=>"000000001",
39735=>"111101101",
39736=>"100011111",
39737=>"111001000",
39738=>"111000111",
39739=>"000011111",
39740=>"011011010",
39741=>"001111111",
39742=>"000000000",
39743=>"001101110",
39744=>"010100111",
39745=>"001111110",
39746=>"000000000",
39747=>"100000100",
39748=>"111100000",
39749=>"000000000",
39750=>"100110111",
39751=>"001001011",
39752=>"011110001",
39753=>"011111001",
39754=>"101001000",
39755=>"111100000",
39756=>"111000000",
39757=>"000010001",
39758=>"110001111",
39759=>"001001011",
39760=>"000000000",
39761=>"101111111",
39762=>"111111010",
39763=>"101111010",
39764=>"000001111",
39765=>"000010011",
39766=>"000111110",
39767=>"101001111",
39768=>"111000010",
39769=>"110000001",
39770=>"101011011",
39771=>"010101000",
39772=>"000111111",
39773=>"100000101",
39774=>"111111100",
39775=>"001000001",
39776=>"001000000",
39777=>"010000101",
39778=>"000001000",
39779=>"011000000",
39780=>"111110111",
39781=>"101111000",
39782=>"110110001",
39783=>"111010010",
39784=>"011101000",
39785=>"110010101",
39786=>"000111100",
39787=>"001000111",
39788=>"010001111",
39789=>"000000001",
39790=>"000000111",
39791=>"111101000",
39792=>"001011010",
39793=>"111111111",
39794=>"000000001",
39795=>"000000000",
39796=>"001000000",
39797=>"011000110",
39798=>"001111001",
39799=>"000000111",
39800=>"111011001",
39801=>"100101111",
39802=>"111111110",
39803=>"100000000",
39804=>"001011011",
39805=>"011000000",
39806=>"000000001",
39807=>"001000000",
39808=>"010100000",
39809=>"001001000",
39810=>"000011011",
39811=>"111000111",
39812=>"000110000",
39813=>"010110110",
39814=>"100111100",
39815=>"111100101",
39816=>"001101000",
39817=>"110111010",
39818=>"001111111",
39819=>"001000101",
39820=>"111000000",
39821=>"001001001",
39822=>"001111111",
39823=>"110000000",
39824=>"111110010",
39825=>"011111000",
39826=>"111111001",
39827=>"111111111",
39828=>"111101001",
39829=>"000000001",
39830=>"000000000",
39831=>"101100111",
39832=>"001000010",
39833=>"000100111",
39834=>"001111111",
39835=>"001001011",
39836=>"111101100",
39837=>"000100000",
39838=>"011111110",
39839=>"111000000",
39840=>"000010011",
39841=>"000000000",
39842=>"001000000",
39843=>"000000000",
39844=>"000111111",
39845=>"101000010",
39846=>"011111111",
39847=>"000111011",
39848=>"000000100",
39849=>"101001111",
39850=>"000000001",
39851=>"100000000",
39852=>"000101111",
39853=>"000000000",
39854=>"000000000",
39855=>"000000110",
39856=>"000001000",
39857=>"000100101",
39858=>"111111101",
39859=>"011010011",
39860=>"111010000",
39861=>"110111011",
39862=>"010000001",
39863=>"111111111",
39864=>"100100100",
39865=>"011110011",
39866=>"110110110",
39867=>"000000011",
39868=>"111111111",
39869=>"110000010",
39870=>"010001000",
39871=>"000001011",
39872=>"010000000",
39873=>"000000111",
39874=>"111010011",
39875=>"000000000",
39876=>"111111111",
39877=>"011010111",
39878=>"000001001",
39879=>"001001111",
39880=>"000000111",
39881=>"000000000",
39882=>"000000000",
39883=>"000001111",
39884=>"000000000",
39885=>"100100100",
39886=>"111111111",
39887=>"110001111",
39888=>"000000000",
39889=>"001001100",
39890=>"110100111",
39891=>"111001001",
39892=>"000001001",
39893=>"000001000",
39894=>"011000000",
39895=>"001001011",
39896=>"011111000",
39897=>"111111000",
39898=>"111101111",
39899=>"000000000",
39900=>"111101100",
39901=>"000000111",
39902=>"000000110",
39903=>"111110000",
39904=>"111001001",
39905=>"101001001",
39906=>"110000001",
39907=>"111010011",
39908=>"011000001",
39909=>"111001100",
39910=>"000100111",
39911=>"001000000",
39912=>"000110000",
39913=>"111001001",
39914=>"000001000",
39915=>"001011111",
39916=>"101011000",
39917=>"000000000",
39918=>"100000101",
39919=>"000000111",
39920=>"000110110",
39921=>"101111111",
39922=>"001001110",
39923=>"010101000",
39924=>"110111000",
39925=>"110000001",
39926=>"000000000",
39927=>"111111110",
39928=>"111000000",
39929=>"001010110",
39930=>"111111111",
39931=>"111110111",
39932=>"111010011",
39933=>"110111111",
39934=>"000111111",
39935=>"010000000",
39936=>"011001100",
39937=>"000001000",
39938=>"101100111",
39939=>"101101011",
39940=>"111101110",
39941=>"011000111",
39942=>"101100000",
39943=>"001010010",
39944=>"000000000",
39945=>"000000010",
39946=>"001001101",
39947=>"101000000",
39948=>"111000000",
39949=>"010010000",
39950=>"001011000",
39951=>"100100101",
39952=>"000000000",
39953=>"111000010",
39954=>"001011000",
39955=>"111011000",
39956=>"111011101",
39957=>"100100111",
39958=>"100101100",
39959=>"111101000",
39960=>"001000010",
39961=>"011011111",
39962=>"011111111",
39963=>"111111100",
39964=>"100000000",
39965=>"000000011",
39966=>"101010010",
39967=>"000001111",
39968=>"000001101",
39969=>"111111111",
39970=>"111100000",
39971=>"111000000",
39972=>"011011011",
39973=>"011000111",
39974=>"111011111",
39975=>"000101111",
39976=>"111110000",
39977=>"010010000",
39978=>"000100000",
39979=>"011000000",
39980=>"001011111",
39981=>"001010011",
39982=>"111111111",
39983=>"000101100",
39984=>"001000111",
39985=>"111110100",
39986=>"010111011",
39987=>"100000111",
39988=>"011010001",
39989=>"000111000",
39990=>"000000001",
39991=>"000000010",
39992=>"101000000",
39993=>"001000100",
39994=>"000100000",
39995=>"101101111",
39996=>"111111111",
39997=>"001101101",
39998=>"010000000",
39999=>"011011110",
40000=>"111000000",
40001=>"111010000",
40002=>"010111111",
40003=>"111110000",
40004=>"000000111",
40005=>"000000000",
40006=>"010001111",
40007=>"111111000",
40008=>"010111111",
40009=>"100100000",
40010=>"001000000",
40011=>"000100111",
40012=>"000000000",
40013=>"101010000",
40014=>"111111111",
40015=>"100000001",
40016=>"000111111",
40017=>"011000000",
40018=>"011101111",
40019=>"011000100",
40020=>"111001111",
40021=>"011011111",
40022=>"111011000",
40023=>"100111110",
40024=>"111000000",
40025=>"100100100",
40026=>"100000011",
40027=>"111100000",
40028=>"000010000",
40029=>"000001111",
40030=>"010010010",
40031=>"011011000",
40032=>"111111010",
40033=>"000000111",
40034=>"010000101",
40035=>"000000100",
40036=>"000000000",
40037=>"111111100",
40038=>"110111100",
40039=>"100111100",
40040=>"000001011",
40041=>"111001111",
40042=>"011111010",
40043=>"011111000",
40044=>"000110111",
40045=>"001001000",
40046=>"000000111",
40047=>"011000011",
40048=>"001011110",
40049=>"010010110",
40050=>"010100100",
40051=>"111111111",
40052=>"100111100",
40053=>"001000000",
40054=>"100000000",
40055=>"111000000",
40056=>"111111000",
40057=>"111111000",
40058=>"000000101",
40059=>"101001011",
40060=>"000010011",
40061=>"110100001",
40062=>"110000001",
40063=>"000000000",
40064=>"101010000",
40065=>"000000011",
40066=>"110000001",
40067=>"000000000",
40068=>"111011100",
40069=>"011100000",
40070=>"011101111",
40071=>"010000110",
40072=>"100000011",
40073=>"000000111",
40074=>"111101100",
40075=>"111111000",
40076=>"000000111",
40077=>"000001111",
40078=>"000000010",
40079=>"000000000",
40080=>"000000001",
40081=>"001001010",
40082=>"101101111",
40083=>"111101100",
40084=>"100100100",
40085=>"111000000",
40086=>"000101111",
40087=>"011001000",
40088=>"101100000",
40089=>"000111011",
40090=>"111010010",
40091=>"100100011",
40092=>"000000000",
40093=>"111111111",
40094=>"111000110",
40095=>"000000000",
40096=>"000010011",
40097=>"100100111",
40098=>"111000000",
40099=>"111111111",
40100=>"000101000",
40101=>"010001001",
40102=>"111111000",
40103=>"001111110",
40104=>"000010111",
40105=>"000111011",
40106=>"101100000",
40107=>"101000010",
40108=>"111011000",
40109=>"111000100",
40110=>"101001010",
40111=>"110010000",
40112=>"000000000",
40113=>"100001001",
40114=>"000101111",
40115=>"000100000",
40116=>"100101000",
40117=>"100100011",
40118=>"000000000",
40119=>"110111111",
40120=>"001111110",
40121=>"011001001",
40122=>"101110111",
40123=>"111110011",
40124=>"001010001",
40125=>"000011110",
40126=>"001001100",
40127=>"001000011",
40128=>"000000111",
40129=>"101000101",
40130=>"101111111",
40131=>"000010000",
40132=>"000101000",
40133=>"001011111",
40134=>"000010000",
40135=>"000100111",
40136=>"000011000",
40137=>"000000000",
40138=>"111101110",
40139=>"101100010",
40140=>"101100101",
40141=>"010000111",
40142=>"000000111",
40143=>"111111000",
40144=>"111001101",
40145=>"110110110",
40146=>"111100000",
40147=>"101100000",
40148=>"000000111",
40149=>"000100111",
40150=>"111111111",
40151=>"111000000",
40152=>"111011100",
40153=>"001011000",
40154=>"000100100",
40155=>"001000001",
40156=>"010010111",
40157=>"100011010",
40158=>"110100011",
40159=>"110010010",
40160=>"010000000",
40161=>"100000111",
40162=>"111100000",
40163=>"101111000",
40164=>"111000111",
40165=>"000111111",
40166=>"011000000",
40167=>"000100111",
40168=>"111000101",
40169=>"000010111",
40170=>"001001111",
40171=>"000000110",
40172=>"011010000",
40173=>"111000001",
40174=>"000000000",
40175=>"000000110",
40176=>"000110000",
40177=>"100011010",
40178=>"001110000",
40179=>"101101011",
40180=>"110001000",
40181=>"111100110",
40182=>"001111011",
40183=>"101000000",
40184=>"000000111",
40185=>"100001000",
40186=>"111001111",
40187=>"100101000",
40188=>"000010000",
40189=>"001101000",
40190=>"110101000",
40191=>"101011000",
40192=>"000111111",
40193=>"111000111",
40194=>"000100011",
40195=>"111010000",
40196=>"110111111",
40197=>"001000000",
40198=>"000110111",
40199=>"100111010",
40200=>"000110111",
40201=>"100010111",
40202=>"000000000",
40203=>"100001111",
40204=>"000000101",
40205=>"000010101",
40206=>"011101001",
40207=>"011100111",
40208=>"111000010",
40209=>"000000011",
40210=>"110101101",
40211=>"001011111",
40212=>"111101001",
40213=>"001001001",
40214=>"101100100",
40215=>"000100100",
40216=>"000000111",
40217=>"010111111",
40218=>"000000000",
40219=>"000011011",
40220=>"001001100",
40221=>"110010000",
40222=>"101101000",
40223=>"111000000",
40224=>"001000001",
40225=>"101111111",
40226=>"100111111",
40227=>"000100000",
40228=>"000100101",
40229=>"100000100",
40230=>"000000000",
40231=>"000001111",
40232=>"111111110",
40233=>"000101111",
40234=>"111000000",
40235=>"110000001",
40236=>"110000001",
40237=>"111101101",
40238=>"000101111",
40239=>"000111010",
40240=>"001010011",
40241=>"001011101",
40242=>"000000110",
40243=>"001111110",
40244=>"010000101",
40245=>"111010110",
40246=>"000000000",
40247=>"100000000",
40248=>"101101010",
40249=>"001101000",
40250=>"010000000",
40251=>"101111110",
40252=>"000000000",
40253=>"000010101",
40254=>"001000000",
40255=>"100000000",
40256=>"000111111",
40257=>"100101000",
40258=>"111010010",
40259=>"100101000",
40260=>"011000111",
40261=>"010001111",
40262=>"010010000",
40263=>"010010111",
40264=>"101100100",
40265=>"011111101",
40266=>"101001000",
40267=>"000111011",
40268=>"000000000",
40269=>"001101000",
40270=>"100100101",
40271=>"001100111",
40272=>"111000000",
40273=>"000011111",
40274=>"000010111",
40275=>"000001000",
40276=>"100000001",
40277=>"100100100",
40278=>"101101100",
40279=>"100000100",
40280=>"110110000",
40281=>"110000011",
40282=>"111001000",
40283=>"100100100",
40284=>"000101100",
40285=>"011101100",
40286=>"011101101",
40287=>"011100000",
40288=>"110101100",
40289=>"000101111",
40290=>"101000100",
40291=>"111110000",
40292=>"111110000",
40293=>"001100000",
40294=>"000110001",
40295=>"111010010",
40296=>"110111110",
40297=>"111111011",
40298=>"101101110",
40299=>"010000000",
40300=>"000100001",
40301=>"110010110",
40302=>"011111011",
40303=>"000101001",
40304=>"101101101",
40305=>"111100010",
40306=>"000000000",
40307=>"000000100",
40308=>"101011010",
40309=>"001000000",
40310=>"111011010",
40311=>"000101101",
40312=>"111100010",
40313=>"111101101",
40314=>"110110111",
40315=>"101111101",
40316=>"111000111",
40317=>"000110000",
40318=>"111110110",
40319=>"000000000",
40320=>"101101011",
40321=>"100101111",
40322=>"000101100",
40323=>"010000010",
40324=>"111111000",
40325=>"010111011",
40326=>"001001001",
40327=>"001001111",
40328=>"001101101",
40329=>"001010010",
40330=>"101010011",
40331=>"000000010",
40332=>"011010000",
40333=>"000010011",
40334=>"110011011",
40335=>"100000010",
40336=>"101101100",
40337=>"111001010",
40338=>"100000000",
40339=>"000001101",
40340=>"011010011",
40341=>"101000010",
40342=>"011011100",
40343=>"011000000",
40344=>"010010011",
40345=>"111110000",
40346=>"000010111",
40347=>"000000011",
40348=>"011000010",
40349=>"000000100",
40350=>"111000100",
40351=>"010010111",
40352=>"101101001",
40353=>"111010000",
40354=>"110000100",
40355=>"101001010",
40356=>"110101000",
40357=>"001100100",
40358=>"010010011",
40359=>"001010110",
40360=>"110000110",
40361=>"010010110",
40362=>"010100000",
40363=>"101000000",
40364=>"111100101",
40365=>"010000000",
40366=>"000011000",
40367=>"000000000",
40368=>"011011011",
40369=>"010001111",
40370=>"010110101",
40371=>"111001110",
40372=>"010011001",
40373=>"000000011",
40374=>"011100100",
40375=>"011101000",
40376=>"000001101",
40377=>"110010110",
40378=>"010010010",
40379=>"001111101",
40380=>"111111111",
40381=>"010001110",
40382=>"000001101",
40383=>"000010010",
40384=>"101101101",
40385=>"000000000",
40386=>"110111000",
40387=>"001001001",
40388=>"110111111",
40389=>"100011001",
40390=>"111110000",
40391=>"000010111",
40392=>"111010111",
40393=>"000101000",
40394=>"011111111",
40395=>"110101110",
40396=>"100111111",
40397=>"111000011",
40398=>"010000101",
40399=>"010111010",
40400=>"011011000",
40401=>"111101100",
40402=>"010111111",
40403=>"011110000",
40404=>"100101101",
40405=>"110000101",
40406=>"101101000",
40407=>"111100000",
40408=>"101101000",
40409=>"000010101",
40410=>"101110111",
40411=>"000010010",
40412=>"101001001",
40413=>"010000000",
40414=>"010000010",
40415=>"001001111",
40416=>"001000100",
40417=>"011010111",
40418=>"010010010",
40419=>"111001000",
40420=>"000000000",
40421=>"111111011",
40422=>"011011111",
40423=>"010110000",
40424=>"100101101",
40425=>"010000000",
40426=>"000000000",
40427=>"010000001",
40428=>"000000000",
40429=>"000000011",
40430=>"000000110",
40431=>"101101101",
40432=>"000010011",
40433=>"001100100",
40434=>"000101011",
40435=>"110100000",
40436=>"100110110",
40437=>"111010000",
40438=>"000000111",
40439=>"111111111",
40440=>"100101101",
40441=>"111110111",
40442=>"010111101",
40443=>"101011011",
40444=>"001100100",
40445=>"110111100",
40446=>"100001101",
40447=>"101011000",
40448=>"000000000",
40449=>"000001000",
40450=>"101101101",
40451=>"000001000",
40452=>"111100000",
40453=>"111001000",
40454=>"011011000",
40455=>"010111111",
40456=>"001110110",
40457=>"000010110",
40458=>"011001100",
40459=>"000010101",
40460=>"111000101",
40461=>"111010000",
40462=>"011000000",
40463=>"010000000",
40464=>"010000000",
40465=>"010000111",
40466=>"010101100",
40467=>"011000000",
40468=>"000111011",
40469=>"000101111",
40470=>"011101001",
40471=>"011010100",
40472=>"000000000",
40473=>"100000101",
40474=>"101101001",
40475=>"001001010",
40476=>"000000110",
40477=>"111110010",
40478=>"001101000",
40479=>"101111011",
40480=>"000101000",
40481=>"110110000",
40482=>"101101100",
40483=>"110100000",
40484=>"100111000",
40485=>"100100100",
40486=>"000000000",
40487=>"110110000",
40488=>"001111111",
40489=>"000000100",
40490=>"000000111",
40491=>"000110000",
40492=>"011110110",
40493=>"010000011",
40494=>"100000000",
40495=>"000111010",
40496=>"101100100",
40497=>"010100000",
40498=>"101101100",
40499=>"101101000",
40500=>"001000101",
40501=>"101101111",
40502=>"010111110",
40503=>"000001011",
40504=>"000000000",
40505=>"000000000",
40506=>"000101100",
40507=>"110111101",
40508=>"110101011",
40509=>"111111111",
40510=>"100001000",
40511=>"011110100",
40512=>"111111101",
40513=>"010100100",
40514=>"111010011",
40515=>"011100100",
40516=>"010000001",
40517=>"000100000",
40518=>"111000011",
40519=>"000101010",
40520=>"011111101",
40521=>"001001010",
40522=>"101101000",
40523=>"010110000",
40524=>"110000011",
40525=>"110110000",
40526=>"001000100",
40527=>"010101000",
40528=>"000101000",
40529=>"111111011",
40530=>"101101111",
40531=>"011011000",
40532=>"000000101",
40533=>"111111111",
40534=>"000100111",
40535=>"101010010",
40536=>"001101101",
40537=>"001000001",
40538=>"100011011",
40539=>"001011000",
40540=>"000010000",
40541=>"001001001",
40542=>"111011001",
40543=>"000001001",
40544=>"000000100",
40545=>"000100110",
40546=>"111100101",
40547=>"000111110",
40548=>"111110000",
40549=>"001001111",
40550=>"010000001",
40551=>"000010010",
40552=>"100100000",
40553=>"111101000",
40554=>"000010111",
40555=>"111111101",
40556=>"000110111",
40557=>"011000000",
40558=>"000001010",
40559=>"010000111",
40560=>"100001001",
40561=>"001000110",
40562=>"010011011",
40563=>"001000000",
40564=>"111010000",
40565=>"000001000",
40566=>"111001000",
40567=>"000010110",
40568=>"000100100",
40569=>"101111110",
40570=>"111100101",
40571=>"111101101",
40572=>"111110011",
40573=>"010100000",
40574=>"010110011",
40575=>"000101101",
40576=>"010000000",
40577=>"000101000",
40578=>"010111101",
40579=>"111101000",
40580=>"011000000",
40581=>"111111111",
40582=>"000011000",
40583=>"000010000",
40584=>"110001111",
40585=>"111000000",
40586=>"010000110",
40587=>"010010111",
40588=>"000111110",
40589=>"100101000",
40590=>"011100110",
40591=>"000000000",
40592=>"101100000",
40593=>"101101101",
40594=>"010111111",
40595=>"000000000",
40596=>"000000000",
40597=>"001010110",
40598=>"100101101",
40599=>"001000000",
40600=>"111000000",
40601=>"101111011",
40602=>"100000111",
40603=>"111010000",
40604=>"000010001",
40605=>"011001101",
40606=>"000000111",
40607=>"110000000",
40608=>"010110111",
40609=>"000101111",
40610=>"101101001",
40611=>"111101000",
40612=>"001000001",
40613=>"100110000",
40614=>"111111000",
40615=>"000000010",
40616=>"001001001",
40617=>"000000001",
40618=>"101101111",
40619=>"111000000",
40620=>"111110000",
40621=>"101110111",
40622=>"001001100",
40623=>"101001111",
40624=>"000000000",
40625=>"100100001",
40626=>"001101011",
40627=>"000110110",
40628=>"110111101",
40629=>"010001011",
40630=>"111111001",
40631=>"110000111",
40632=>"001101010",
40633=>"000000000",
40634=>"010001111",
40635=>"000111011",
40636=>"000010000",
40637=>"111001111",
40638=>"111011001",
40639=>"000000001",
40640=>"001000110",
40641=>"000000000",
40642=>"101000011",
40643=>"110111001",
40644=>"011000000",
40645=>"110011001",
40646=>"010001111",
40647=>"000111111",
40648=>"111100111",
40649=>"011011000",
40650=>"101101010",
40651=>"100100101",
40652=>"000011000",
40653=>"101110110",
40654=>"000010111",
40655=>"111111111",
40656=>"001101111",
40657=>"101011011",
40658=>"000000000",
40659=>"101101001",
40660=>"111011001",
40661=>"001000100",
40662=>"111001101",
40663=>"000010101",
40664=>"001000000",
40665=>"000000111",
40666=>"101000100",
40667=>"111000101",
40668=>"111100000",
40669=>"111011111",
40670=>"111101000",
40671=>"010111011",
40672=>"110000000",
40673=>"001000000",
40674=>"011011011",
40675=>"111100001",
40676=>"001011011",
40677=>"101111110",
40678=>"111000000",
40679=>"000001010",
40680=>"110110000",
40681=>"000110110",
40682=>"100000001",
40683=>"101001000",
40684=>"000010100",
40685=>"110110110",
40686=>"100000101",
40687=>"110111111",
40688=>"110010010",
40689=>"111111110",
40690=>"000001100",
40691=>"111110000",
40692=>"100100001",
40693=>"000011000",
40694=>"000010011",
40695=>"100010111",
40696=>"111001110",
40697=>"101001111",
40698=>"111101000",
40699=>"001010000",
40700=>"100101101",
40701=>"011010111",
40702=>"011001001",
40703=>"110000000",
40704=>"000000000",
40705=>"000001010",
40706=>"000000001",
40707=>"111111101",
40708=>"111111111",
40709=>"111011011",
40710=>"000000010",
40711=>"000000000",
40712=>"110000000",
40713=>"000001101",
40714=>"111110000",
40715=>"010110111",
40716=>"000000001",
40717=>"111111111",
40718=>"110000000",
40719=>"000000000",
40720=>"010010010",
40721=>"110110111",
40722=>"001111000",
40723=>"000101111",
40724=>"000100000",
40725=>"111111111",
40726=>"000000001",
40727=>"000000000",
40728=>"100111000",
40729=>"111110000",
40730=>"110000110",
40731=>"000000010",
40732=>"001001111",
40733=>"000101101",
40734=>"000001000",
40735=>"000000100",
40736=>"000000000",
40737=>"111111000",
40738=>"000000101",
40739=>"100001111",
40740=>"100100101",
40741=>"111111111",
40742=>"111111001",
40743=>"000000111",
40744=>"110110010",
40745=>"000010000",
40746=>"000000000",
40747=>"010110100",
40748=>"000000010",
40749=>"111000000",
40750=>"111110000",
40751=>"001000001",
40752=>"000000000",
40753=>"100111110",
40754=>"100001000",
40755=>"110111111",
40756=>"110010110",
40757=>"000000011",
40758=>"100000110",
40759=>"000000101",
40760=>"111011000",
40761=>"000000000",
40762=>"000000000",
40763=>"110111111",
40764=>"111011011",
40765=>"111111011",
40766=>"000000100",
40767=>"111011011",
40768=>"110111110",
40769=>"111111100",
40770=>"110111111",
40771=>"001010110",
40772=>"000000011",
40773=>"000110111",
40774=>"000000000",
40775=>"000000111",
40776=>"001101100",
40777=>"111111000",
40778=>"000000000",
40779=>"111111111",
40780=>"010011010",
40781=>"111111110",
40782=>"001111111",
40783=>"000000001",
40784=>"111001111",
40785=>"110110010",
40786=>"000100111",
40787=>"001000001",
40788=>"010000000",
40789=>"001101101",
40790=>"001000000",
40791=>"111110100",
40792=>"000000001",
40793=>"000000011",
40794=>"111111110",
40795=>"010110000",
40796=>"111111000",
40797=>"001001000",
40798=>"111111110",
40799=>"001011111",
40800=>"111111000",
40801=>"000000000",
40802=>"001001101",
40803=>"111111000",
40804=>"110110000",
40805=>"110010000",
40806=>"000110000",
40807=>"000010001",
40808=>"000000111",
40809=>"000111010",
40810=>"110111111",
40811=>"111111010",
40812=>"000000001",
40813=>"110010000",
40814=>"000000001",
40815=>"110010010",
40816=>"001110110",
40817=>"111111000",
40818=>"010100110",
40819=>"000110111",
40820=>"001111111",
40821=>"000000001",
40822=>"111110100",
40823=>"111111000",
40824=>"111111010",
40825=>"000110010",
40826=>"001001001",
40827=>"111111111",
40828=>"110000100",
40829=>"100100000",
40830=>"000000010",
40831=>"101000100",
40832=>"001001000",
40833=>"101000000",
40834=>"010011000",
40835=>"011100101",
40836=>"111001010",
40837=>"000001000",
40838=>"110110110",
40839=>"110110111",
40840=>"011011011",
40841=>"000000000",
40842=>"010111011",
40843=>"110111111",
40844=>"110111010",
40845=>"000001001",
40846=>"000000000",
40847=>"001000000",
40848=>"111111111",
40849=>"110010011",
40850=>"111000010",
40851=>"000010000",
40852=>"110110110",
40853=>"001000000",
40854=>"010110001",
40855=>"110010110",
40856=>"011111000",
40857=>"000000001",
40858=>"111111110",
40859=>"000001110",
40860=>"000000000",
40861=>"110110000",
40862=>"100101000",
40863=>"000000000",
40864=>"001001001",
40865=>"010110010",
40866=>"110111010",
40867=>"000000001",
40868=>"110000001",
40869=>"000000000",
40870=>"111011111",
40871=>"000111110",
40872=>"110110001",
40873=>"000111111",
40874=>"001001100",
40875=>"100101110",
40876=>"000000000",
40877=>"111110110",
40878=>"000000000",
40879=>"111001111",
40880=>"111111010",
40881=>"010110100",
40882=>"111111011",
40883=>"000100101",
40884=>"110101111",
40885=>"000000000",
40886=>"111010101",
40887=>"111111111",
40888=>"111100101",
40889=>"111111101",
40890=>"111111011",
40891=>"110111110",
40892=>"000111110",
40893=>"011111111",
40894=>"101100100",
40895=>"110110000",
40896=>"111010000",
40897=>"001001000",
40898=>"110000100",
40899=>"100100110",
40900=>"110000000",
40901=>"100100000",
40902=>"000000000",
40903=>"111111000",
40904=>"110001111",
40905=>"111111000",
40906=>"101001000",
40907=>"000000101",
40908=>"010111110",
40909=>"011010111",
40910=>"010111110",
40911=>"101101011",
40912=>"000000010",
40913=>"101110110",
40914=>"111110010",
40915=>"000000010",
40916=>"111010000",
40917=>"001101001",
40918=>"000000101",
40919=>"000001000",
40920=>"000000000",
40921=>"111101111",
40922=>"000001100",
40923=>"001001111",
40924=>"101111100",
40925=>"101111111",
40926=>"010110000",
40927=>"111111111",
40928=>"111000111",
40929=>"110000000",
40930=>"011110111",
40931=>"000000010",
40932=>"110110010",
40933=>"101111111",
40934=>"100100111",
40935=>"010000000",
40936=>"111111011",
40937=>"010000110",
40938=>"111011000",
40939=>"001000000",
40940=>"110110110",
40941=>"111111111",
40942=>"110010001",
40943=>"001001000",
40944=>"000001111",
40945=>"011010100",
40946=>"000000111",
40947=>"001001111",
40948=>"000001001",
40949=>"110111110",
40950=>"110110100",
40951=>"000001011",
40952=>"011011000",
40953=>"000110110",
40954=>"000000000",
40955=>"010010010",
40956=>"111010000",
40957=>"101101100",
40958=>"100110110",
40959=>"000000000",
40960=>"100101111",
40961=>"101101000",
40962=>"000000000",
40963=>"011000000",
40964=>"010010011",
40965=>"111100100",
40966=>"010011111",
40967=>"011111000",
40968=>"010000101",
40969=>"000101000",
40970=>"010111000",
40971=>"101000000",
40972=>"101000000",
40973=>"000000110",
40974=>"100000111",
40975=>"111110010",
40976=>"100111011",
40977=>"100111111",
40978=>"000000101",
40979=>"000000000",
40980=>"001000000",
40981=>"111100000",
40982=>"110101000",
40983=>"010111111",
40984=>"111001000",
40985=>"111111111",
40986=>"110100101",
40987=>"011101101",
40988=>"110000000",
40989=>"011111110",
40990=>"111111100",
40991=>"000000110",
40992=>"111001001",
40993=>"010000000",
40994=>"000010010",
40995=>"111001101",
40996=>"000000011",
40997=>"001111001",
40998=>"111010000",
40999=>"000101101",
41000=>"000000000",
41001=>"111111111",
41002=>"100111000",
41003=>"000000101",
41004=>"011111000",
41005=>"000101000",
41006=>"111101000",
41007=>"111111111",
41008=>"111010001",
41009=>"010000111",
41010=>"101101001",
41011=>"010011010",
41012=>"000000000",
41013=>"000111111",
41014=>"111110111",
41015=>"010111111",
41016=>"101000000",
41017=>"000000010",
41018=>"000000000",
41019=>"000010111",
41020=>"100110001",
41021=>"010111010",
41022=>"010000011",
41023=>"100000111",
41024=>"111101100",
41025=>"111010001",
41026=>"101101111",
41027=>"001100111",
41028=>"100111010",
41029=>"000101111",
41030=>"011011011",
41031=>"000001111",
41032=>"010000001",
41033=>"000000111",
41034=>"001000000",
41035=>"101000000",
41036=>"000111000",
41037=>"110011000",
41038=>"111111111",
41039=>"000010011",
41040=>"111000000",
41041=>"010111000",
41042=>"011010000",
41043=>"111000111",
41044=>"111111000",
41045=>"001000001",
41046=>"000000110",
41047=>"000111100",
41048=>"100011010",
41049=>"010010010",
41050=>"000110010",
41051=>"100000110",
41052=>"111110000",
41053=>"100100000",
41054=>"000111111",
41055=>"100001111",
41056=>"111101111",
41057=>"111000000",
41058=>"000010000",
41059=>"000010110",
41060=>"110000000",
41061=>"011011111",
41062=>"100000111",
41063=>"001111111",
41064=>"000100101",
41065=>"101111111",
41066=>"111001101",
41067=>"010010111",
41068=>"010000000",
41069=>"000111011",
41070=>"101000000",
41071=>"100000010",
41072=>"000000011",
41073=>"010000111",
41074=>"111111011",
41075=>"000111000",
41076=>"111010011",
41077=>"101000101",
41078=>"000000000",
41079=>"000000000",
41080=>"000100000",
41081=>"111111000",
41082=>"000111111",
41083=>"111000000",
41084=>"000100001",
41085=>"111101111",
41086=>"000100111",
41087=>"101000000",
41088=>"011001000",
41089=>"000000000",
41090=>"111111010",
41091=>"011010111",
41092=>"111111000",
41093=>"010001000",
41094=>"110111100",
41095=>"110011110",
41096=>"110010000",
41097=>"000000111",
41098=>"111111100",
41099=>"000100111",
41100=>"000101010",
41101=>"001100101",
41102=>"101000100",
41103=>"001000010",
41104=>"111001111",
41105=>"100100000",
41106=>"110000001",
41107=>"011000010",
41108=>"100000110",
41109=>"000000010",
41110=>"000110010",
41111=>"011011111",
41112=>"111111111",
41113=>"100111001",
41114=>"101011000",
41115=>"110101111",
41116=>"010000010",
41117=>"001111111",
41118=>"010000111",
41119=>"001000000",
41120=>"000000100",
41121=>"000100111",
41122=>"111000101",
41123=>"111010000",
41124=>"000000101",
41125=>"111000011",
41126=>"011000000",
41127=>"000000000",
41128=>"011111110",
41129=>"000000000",
41130=>"111100100",
41131=>"101000000",
41132=>"001000001",
41133=>"000000001",
41134=>"010010110",
41135=>"000001011",
41136=>"011000100",
41137=>"001110111",
41138=>"111101100",
41139=>"000100100",
41140=>"100100101",
41141=>"010001110",
41142=>"111000000",
41143=>"000010101",
41144=>"000010110",
41145=>"001000011",
41146=>"111111000",
41147=>"110110111",
41148=>"000000011",
41149=>"000111111",
41150=>"101111011",
41151=>"000100000",
41152=>"000000010",
41153=>"000010011",
41154=>"000000111",
41155=>"010001101",
41156=>"000000101",
41157=>"000011101",
41158=>"111010000",
41159=>"000000111",
41160=>"111000010",
41161=>"111101101",
41162=>"111011011",
41163=>"001000101",
41164=>"011100111",
41165=>"000011000",
41166=>"010111111",
41167=>"111111111",
41168=>"001111111",
41169=>"111011011",
41170=>"000010111",
41171=>"111100000",
41172=>"000000111",
41173=>"000111000",
41174=>"000000000",
41175=>"111110111",
41176=>"000000010",
41177=>"000000001",
41178=>"011100001",
41179=>"101000011",
41180=>"101100000",
41181=>"000101111",
41182=>"101000101",
41183=>"000000111",
41184=>"111000101",
41185=>"000000101",
41186=>"000101101",
41187=>"111100111",
41188=>"000000101",
41189=>"010000111",
41190=>"111000000",
41191=>"100001001",
41192=>"111000000",
41193=>"111111000",
41194=>"011111100",
41195=>"111111111",
41196=>"000000100",
41197=>"000111000",
41198=>"000000001",
41199=>"111000000",
41200=>"000111001",
41201=>"010110000",
41202=>"000000100",
41203=>"010011001",
41204=>"111110111",
41205=>"101111010",
41206=>"100011010",
41207=>"111001101",
41208=>"000000010",
41209=>"000001000",
41210=>"111111111",
41211=>"010111111",
41212=>"111111100",
41213=>"000001111",
41214=>"100000011",
41215=>"111000000",
41216=>"101100100",
41217=>"001110010",
41218=>"000001111",
41219=>"111000110",
41220=>"111101101",
41221=>"100001110",
41222=>"000100111",
41223=>"000010000",
41224=>"111010010",
41225=>"100101111",
41226=>"101100101",
41227=>"000100000",
41228=>"000101110",
41229=>"110010000",
41230=>"000000000",
41231=>"000111111",
41232=>"111000111",
41233=>"100100111",
41234=>"111111011",
41235=>"000000000",
41236=>"101101111",
41237=>"011011100",
41238=>"011111011",
41239=>"110110000",
41240=>"101111000",
41241=>"000000100",
41242=>"110001000",
41243=>"000101111",
41244=>"110000010",
41245=>"000000000",
41246=>"111000000",
41247=>"000000000",
41248=>"100001111",
41249=>"011111000",
41250=>"110000100",
41251=>"010010000",
41252=>"001001001",
41253=>"111011111",
41254=>"010110000",
41255=>"100001000",
41256=>"111001000",
41257=>"000000000",
41258=>"000101111",
41259=>"010011000",
41260=>"101111001",
41261=>"011000000",
41262=>"111010000",
41263=>"000010101",
41264=>"100101010",
41265=>"111011101",
41266=>"101010001",
41267=>"101000000",
41268=>"110101111",
41269=>"010110111",
41270=>"111001101",
41271=>"100000000",
41272=>"101100111",
41273=>"000000111",
41274=>"101001000",
41275=>"101100000",
41276=>"111111001",
41277=>"111010111",
41278=>"001000101",
41279=>"101000000",
41280=>"100010111",
41281=>"101101011",
41282=>"101101001",
41283=>"111101100",
41284=>"100101111",
41285=>"111000100",
41286=>"001001000",
41287=>"011100100",
41288=>"111110010",
41289=>"111101100",
41290=>"001000111",
41291=>"011010111",
41292=>"000000000",
41293=>"111100010",
41294=>"111100110",
41295=>"101010111",
41296=>"111101101",
41297=>"011111111",
41298=>"111101110",
41299=>"010001000",
41300=>"000010001",
41301=>"010010000",
41302=>"111100000",
41303=>"101000111",
41304=>"001010000",
41305=>"000001001",
41306=>"000000000",
41307=>"101011100",
41308=>"000000001",
41309=>"011001000",
41310=>"011111111",
41311=>"100101001",
41312=>"010010000",
41313=>"010010101",
41314=>"001101111",
41315=>"110010000",
41316=>"101001000",
41317=>"100101101",
41318=>"111110000",
41319=>"000000111",
41320=>"010010000",
41321=>"111111000",
41322=>"101111110",
41323=>"110000110",
41324=>"100010000",
41325=>"001101001",
41326=>"011010010",
41327=>"101111000",
41328=>"101100000",
41329=>"001101000",
41330=>"111100000",
41331=>"000000101",
41332=>"101010000",
41333=>"000000110",
41334=>"001101110",
41335=>"000000000",
41336=>"000010000",
41337=>"000000001",
41338=>"101100111",
41339=>"000101001",
41340=>"100001100",
41341=>"010010000",
41342=>"010111100",
41343=>"100101101",
41344=>"111101001",
41345=>"101100000",
41346=>"100000001",
41347=>"100010111",
41348=>"111000100",
41349=>"000000101",
41350=>"100100010",
41351=>"000000100",
41352=>"101100011",
41353=>"001100111",
41354=>"101000101",
41355=>"000100111",
41356=>"011111101",
41357=>"111111101",
41358=>"000111101",
41359=>"000000000",
41360=>"111001000",
41361=>"000000000",
41362=>"010000000",
41363=>"010110000",
41364=>"111100000",
41365=>"101001111",
41366=>"111000101",
41367=>"111001000",
41368=>"011000011",
41369=>"011010011",
41370=>"101100101",
41371=>"000000001",
41372=>"001100010",
41373=>"000000111",
41374=>"100100011",
41375=>"000101100",
41376=>"011011001",
41377=>"100010011",
41378=>"011111000",
41379=>"000011111",
41380=>"001011000",
41381=>"101100001",
41382=>"111001101",
41383=>"011011000",
41384=>"011101100",
41385=>"010100000",
41386=>"000101111",
41387=>"101000111",
41388=>"011111000",
41389=>"101101111",
41390=>"011011001",
41391=>"000000111",
41392=>"010010111",
41393=>"110000000",
41394=>"100101000",
41395=>"100001000",
41396=>"111011000",
41397=>"010010100",
41398=>"111100100",
41399=>"110100000",
41400=>"011111110",
41401=>"110001000",
41402=>"111010110",
41403=>"011000101",
41404=>"111110101",
41405=>"101111101",
41406=>"111000000",
41407=>"010000000",
41408=>"001100000",
41409=>"000000111",
41410=>"111111000",
41411=>"100101100",
41412=>"000000100",
41413=>"111111100",
41414=>"100011011",
41415=>"101101111",
41416=>"010010101",
41417=>"001010100",
41418=>"000000000",
41419=>"111010110",
41420=>"100101111",
41421=>"111110001",
41422=>"000101110",
41423=>"001010011",
41424=>"000000111",
41425=>"111100000",
41426=>"000000000",
41427=>"001010000",
41428=>"000000111",
41429=>"110110000",
41430=>"111000000",
41431=>"001000101",
41432=>"010011100",
41433=>"111111110",
41434=>"100110100",
41435=>"000100111",
41436=>"110100000",
41437=>"011011001",
41438=>"111101101",
41439=>"101101001",
41440=>"100101100",
41441=>"000000011",
41442=>"110010101",
41443=>"111101001",
41444=>"101000001",
41445=>"111111000",
41446=>"100101110",
41447=>"000110000",
41448=>"101101111",
41449=>"000010000",
41450=>"101100110",
41451=>"111000101",
41452=>"000010110",
41453=>"101100111",
41454=>"100111010",
41455=>"101111000",
41456=>"100000000",
41457=>"111011000",
41458=>"101101010",
41459=>"110110000",
41460=>"111000100",
41461=>"000001101",
41462=>"010000111",
41463=>"000111000",
41464=>"100111011",
41465=>"100010000",
41466=>"111011001",
41467=>"101111000",
41468=>"000101111",
41469=>"000010110",
41470=>"100000101",
41471=>"000101111",
41472=>"011001100",
41473=>"111111101",
41474=>"000000000",
41475=>"001000000",
41476=>"100011011",
41477=>"111000111",
41478=>"111111111",
41479=>"011111111",
41480=>"111111111",
41481=>"001000111",
41482=>"001000001",
41483=>"011101001",
41484=>"000010000",
41485=>"101001001",
41486=>"000000100",
41487=>"001011011",
41488=>"101000111",
41489=>"001000111",
41490=>"111001111",
41491=>"111100000",
41492=>"111111000",
41493=>"001101111",
41494=>"100011001",
41495=>"111111010",
41496=>"101101111",
41497=>"100111110",
41498=>"110010111",
41499=>"000000101",
41500=>"000000001",
41501=>"111101000",
41502=>"110101111",
41503=>"000000000",
41504=>"000000000",
41505=>"011111011",
41506=>"000011110",
41507=>"001011010",
41508=>"111111001",
41509=>"011001001",
41510=>"000111111",
41511=>"101010011",
41512=>"010010000",
41513=>"110111111",
41514=>"101100111",
41515=>"010010000",
41516=>"111111111",
41517=>"001111011",
41518=>"110000010",
41519=>"111000111",
41520=>"111111010",
41521=>"111111000",
41522=>"000010111",
41523=>"111101101",
41524=>"000000000",
41525=>"100110001",
41526=>"111011000",
41527=>"100001000",
41528=>"011010000",
41529=>"000000111",
41530=>"001000111",
41531=>"101111110",
41532=>"001000000",
41533=>"111010000",
41534=>"000000001",
41535=>"110011011",
41536=>"111111111",
41537=>"001101101",
41538=>"111000000",
41539=>"011000000",
41540=>"111111010",
41541=>"001000000",
41542=>"100100000",
41543=>"111011111",
41544=>"111011111",
41545=>"001101111",
41546=>"101000101",
41547=>"101110000",
41548=>"000000000",
41549=>"000110110",
41550=>"101110010",
41551=>"100011000",
41552=>"000100100",
41553=>"111111111",
41554=>"111000111",
41555=>"011000000",
41556=>"000000111",
41557=>"100110110",
41558=>"001010000",
41559=>"000000000",
41560=>"000100101",
41561=>"110001001",
41562=>"000110110",
41563=>"000011011",
41564=>"111110111",
41565=>"100000110",
41566=>"111111110",
41567=>"100000000",
41568=>"000000000",
41569=>"010000101",
41570=>"000000000",
41571=>"001001001",
41572=>"001000001",
41573=>"011001000",
41574=>"000001101",
41575=>"000000101",
41576=>"111111000",
41577=>"111000100",
41578=>"010110111",
41579=>"111010111",
41580=>"001001011",
41581=>"000000101",
41582=>"101101110",
41583=>"000101011",
41584=>"111111100",
41585=>"111000011",
41586=>"011011000",
41587=>"000000000",
41588=>"000011000",
41589=>"111000100",
41590=>"111001011",
41591=>"111111110",
41592=>"000000000",
41593=>"100001001",
41594=>"000010111",
41595=>"000111110",
41596=>"000011001",
41597=>"110000011",
41598=>"011010000",
41599=>"000000000",
41600=>"111011100",
41601=>"000010001",
41602=>"101101101",
41603=>"100111001",
41604=>"101000011",
41605=>"111111000",
41606=>"110100100",
41607=>"100001110",
41608=>"100111001",
41609=>"000000000",
41610=>"100000000",
41611=>"111010111",
41612=>"011000000",
41613=>"100011111",
41614=>"111000000",
41615=>"000000000",
41616=>"010110101",
41617=>"000000000",
41618=>"111000010",
41619=>"111111110",
41620=>"010110100",
41621=>"111000111",
41622=>"111001110",
41623=>"100111111",
41624=>"101011000",
41625=>"111101001",
41626=>"010011010",
41627=>"010000101",
41628=>"000000110",
41629=>"111100001",
41630=>"111000100",
41631=>"011000111",
41632=>"001011111",
41633=>"010000111",
41634=>"000111010",
41635=>"000000000",
41636=>"111111111",
41637=>"000100110",
41638=>"101110100",
41639=>"000000111",
41640=>"110101000",
41641=>"000000001",
41642=>"010000000",
41643=>"000000111",
41644=>"101111010",
41645=>"000000111",
41646=>"000000001",
41647=>"010000001",
41648=>"001011001",
41649=>"111111111",
41650=>"010000000",
41651=>"001000011",
41652=>"101001011",
41653=>"101011000",
41654=>"111001101",
41655=>"001111000",
41656=>"000000000",
41657=>"111011001",
41658=>"000000000",
41659=>"111000000",
41660=>"000000001",
41661=>"110111110",
41662=>"110111000",
41663=>"000000000",
41664=>"000000111",
41665=>"101000000",
41666=>"110111001",
41667=>"110001000",
41668=>"010111101",
41669=>"101111111",
41670=>"001000000",
41671=>"110010000",
41672=>"111111100",
41673=>"000011000",
41674=>"010011000",
41675=>"101111000",
41676=>"011101101",
41677=>"000010110",
41678=>"101101101",
41679=>"111010011",
41680=>"111000000",
41681=>"000111011",
41682=>"001000000",
41683=>"001111011",
41684=>"000000000",
41685=>"011001001",
41686=>"000000000",
41687=>"011000100",
41688=>"111111000",
41689=>"000110000",
41690=>"100110010",
41691=>"110000101",
41692=>"000000110",
41693=>"111000101",
41694=>"010100000",
41695=>"111111000",
41696=>"100000000",
41697=>"000000011",
41698=>"111010010",
41699=>"001111111",
41700=>"000000001",
41701=>"000111000",
41702=>"010111101",
41703=>"000001100",
41704=>"011000111",
41705=>"000001000",
41706=>"100000100",
41707=>"000110000",
41708=>"111111001",
41709=>"010000110",
41710=>"010000000",
41711=>"000011010",
41712=>"001111000",
41713=>"111011111",
41714=>"111111111",
41715=>"111110110",
41716=>"110011111",
41717=>"101101101",
41718=>"000000101",
41719=>"001000000",
41720=>"001111010",
41721=>"000110111",
41722=>"110011000",
41723=>"000011111",
41724=>"010010000",
41725=>"111011111",
41726=>"001011111",
41727=>"110110111",
41728=>"111010000",
41729=>"000000111",
41730=>"101000001",
41731=>"111000101",
41732=>"011101111",
41733=>"101000000",
41734=>"010011011",
41735=>"001000101",
41736=>"011110111",
41737=>"111011001",
41738=>"010000111",
41739=>"101001101",
41740=>"000010000",
41741=>"101100000",
41742=>"100011011",
41743=>"011111001",
41744=>"000010110",
41745=>"010000000",
41746=>"000001000",
41747=>"000000110",
41748=>"111111101",
41749=>"011000000",
41750=>"100100111",
41751=>"000000110",
41752=>"000001101",
41753=>"101011101",
41754=>"111111010",
41755=>"111111000",
41756=>"110110101",
41757=>"000000000",
41758=>"110010000",
41759=>"011000000",
41760=>"000110000",
41761=>"000111011",
41762=>"000111011",
41763=>"111000000",
41764=>"110111000",
41765=>"110110000",
41766=>"000000000",
41767=>"111111111",
41768=>"110110111",
41769=>"110111111",
41770=>"000100111",
41771=>"011000000",
41772=>"000011011",
41773=>"101010011",
41774=>"111111111",
41775=>"000000000",
41776=>"111000000",
41777=>"000100000",
41778=>"000000110",
41779=>"001110111",
41780=>"110000000",
41781=>"111111000",
41782=>"100011011",
41783=>"000000101",
41784=>"010000000",
41785=>"101000001",
41786=>"011000101",
41787=>"000000010",
41788=>"110110110",
41789=>"010111110",
41790=>"000010000",
41791=>"110011010",
41792=>"001101111",
41793=>"111010001",
41794=>"000000101",
41795=>"000110110",
41796=>"000111111",
41797=>"101000110",
41798=>"011111000",
41799=>"111000000",
41800=>"000001000",
41801=>"011000111",
41802=>"101000001",
41803=>"111111100",
41804=>"010010110",
41805=>"001001000",
41806=>"000101100",
41807=>"010111110",
41808=>"101000000",
41809=>"000000001",
41810=>"111101111",
41811=>"011100100",
41812=>"111111111",
41813=>"000110110",
41814=>"111011001",
41815=>"111010000",
41816=>"111100011",
41817=>"100110110",
41818=>"001110000",
41819=>"111111000",
41820=>"000110111",
41821=>"111001000",
41822=>"011111011",
41823=>"000011011",
41824=>"000111111",
41825=>"001010000",
41826=>"111110101",
41827=>"000111111",
41828=>"111111000",
41829=>"011001000",
41830=>"101111111",
41831=>"011001001",
41832=>"000000001",
41833=>"011010001",
41834=>"110010111",
41835=>"000101101",
41836=>"011000110",
41837=>"101000111",
41838=>"011001000",
41839=>"111010111",
41840=>"000101000",
41841=>"010010111",
41842=>"001100100",
41843=>"110000000",
41844=>"000100111",
41845=>"000000101",
41846=>"000000000",
41847=>"111111111",
41848=>"000111111",
41849=>"111001001",
41850=>"000101111",
41851=>"100000000",
41852=>"000110110",
41853=>"110100000",
41854=>"011101000",
41855=>"011000000",
41856=>"001000000",
41857=>"010000000",
41858=>"111111000",
41859=>"111110101",
41860=>"011111111",
41861=>"110111000",
41862=>"110011000",
41863=>"001010000",
41864=>"100101100",
41865=>"010000000",
41866=>"000000000",
41867=>"101000000",
41868=>"000111001",
41869=>"011111110",
41870=>"010010010",
41871=>"000001000",
41872=>"001001000",
41873=>"010010000",
41874=>"011001101",
41875=>"011001111",
41876=>"000011111",
41877=>"000010111",
41878=>"111101111",
41879=>"000011011",
41880=>"000000000",
41881=>"001010111",
41882=>"000111111",
41883=>"000000101",
41884=>"000010000",
41885=>"010111110",
41886=>"000000110",
41887=>"000000100",
41888=>"000000000",
41889=>"000010000",
41890=>"000000000",
41891=>"111111101",
41892=>"111010000",
41893=>"000000000",
41894=>"101111111",
41895=>"110111000",
41896=>"001000010",
41897=>"000111000",
41898=>"111110101",
41899=>"000000000",
41900=>"101001111",
41901=>"101001000",
41902=>"110000000",
41903=>"101110011",
41904=>"000101000",
41905=>"101011100",
41906=>"000000010",
41907=>"001100100",
41908=>"111101000",
41909=>"101010010",
41910=>"111101100",
41911=>"111111010",
41912=>"001011010",
41913=>"000100111",
41914=>"000100101",
41915=>"111010011",
41916=>"111111000",
41917=>"000111111",
41918=>"011111100",
41919=>"111000000",
41920=>"111010000",
41921=>"111001000",
41922=>"010101111",
41923=>"000100100",
41924=>"010000000",
41925=>"000001001",
41926=>"010001010",
41927=>"000000000",
41928=>"111101000",
41929=>"000000000",
41930=>"011001101",
41931=>"000000001",
41932=>"000000000",
41933=>"000011011",
41934=>"001101101",
41935=>"000111100",
41936=>"111001000",
41937=>"111110100",
41938=>"111000111",
41939=>"000001001",
41940=>"100010010",
41941=>"111100000",
41942=>"000000110",
41943=>"010010110",
41944=>"000001011",
41945=>"000000111",
41946=>"001000101",
41947=>"001000101",
41948=>"001011111",
41949=>"100011000",
41950=>"111111010",
41951=>"100000110",
41952=>"000010001",
41953=>"111000111",
41954=>"111101000",
41955=>"111111100",
41956=>"000010000",
41957=>"000000111",
41958=>"111000000",
41959=>"011000000",
41960=>"000000101",
41961=>"001111111",
41962=>"010000111",
41963=>"001111110",
41964=>"000000101",
41965=>"000000000",
41966=>"000010000",
41967=>"000000000",
41968=>"000000011",
41969=>"000000110",
41970=>"110000000",
41971=>"011011001",
41972=>"100111001",
41973=>"000101000",
41974=>"000000000",
41975=>"000101111",
41976=>"000010110",
41977=>"101101111",
41978=>"010111100",
41979=>"000101011",
41980=>"000010110",
41981=>"000000001",
41982=>"000100011",
41983=>"000000000",
41984=>"000001100",
41985=>"000100101",
41986=>"100100010",
41987=>"111101111",
41988=>"001101010",
41989=>"100101100",
41990=>"100010111",
41991=>"011011111",
41992=>"001001101",
41993=>"100111111",
41994=>"100100101",
41995=>"000000011",
41996=>"011011011",
41997=>"011011001",
41998=>"101101001",
41999=>"000000001",
42000=>"010011000",
42001=>"110100000",
42002=>"101000101",
42003=>"100000010",
42004=>"111000000",
42005=>"111111111",
42006=>"000011111",
42007=>"100100000",
42008=>"100100100",
42009=>"000000001",
42010=>"000011100",
42011=>"100111011",
42012=>"100110011",
42013=>"000001111",
42014=>"111001111",
42015=>"011001000",
42016=>"110010110",
42017=>"000111110",
42018=>"000011011",
42019=>"000101111",
42020=>"100100110",
42021=>"110101011",
42022=>"000100011",
42023=>"100110110",
42024=>"111111011",
42025=>"011001010",
42026=>"100100110",
42027=>"000100101",
42028=>"111011011",
42029=>"101011111",
42030=>"111000001",
42031=>"000000100",
42032=>"111101111",
42033=>"111110110",
42034=>"000001000",
42035=>"000011001",
42036=>"000000000",
42037=>"011010011",
42038=>"000101101",
42039=>"011110000",
42040=>"111101011",
42041=>"000100100",
42042=>"000000000",
42043=>"100011011",
42044=>"011011101",
42045=>"011011001",
42046=>"000000011",
42047=>"101001011",
42048=>"011011001",
42049=>"000011001",
42050=>"100110000",
42051=>"000000101",
42052=>"000000000",
42053=>"011000000",
42054=>"100100111",
42055=>"110111011",
42056=>"111110110",
42057=>"001111000",
42058=>"000110100",
42059=>"011011001",
42060=>"000000000",
42061=>"011111111",
42062=>"111001101",
42063=>"111011001",
42064=>"100100100",
42065=>"000111111",
42066=>"011000000",
42067=>"000000000",
42068=>"100010011",
42069=>"110111111",
42070=>"100100000",
42071=>"100100100",
42072=>"111011000",
42073=>"010010011",
42074=>"110000110",
42075=>"011111100",
42076=>"110111110",
42077=>"000000000",
42078=>"111100000",
42079=>"110101100",
42080=>"000110110",
42081=>"010110100",
42082=>"100110111",
42083=>"100000101",
42084=>"010000010",
42085=>"000100100",
42086=>"111111000",
42087=>"111010011",
42088=>"000111111",
42089=>"110100001",
42090=>"111010011",
42091=>"011101000",
42092=>"101111001",
42093=>"111000000",
42094=>"100110111",
42095=>"011111000",
42096=>"000111010",
42097=>"100101000",
42098=>"000110100",
42099=>"011000100",
42100=>"101100000",
42101=>"100100000",
42102=>"011011011",
42103=>"011111101",
42104=>"100100110",
42105=>"000100000",
42106=>"011110000",
42107=>"110001111",
42108=>"110010111",
42109=>"110110111",
42110=>"000011111",
42111=>"100110011",
42112=>"000100000",
42113=>"100111111",
42114=>"110110000",
42115=>"011101000",
42116=>"111011011",
42117=>"000011111",
42118=>"000100010",
42119=>"000110001",
42120=>"110101001",
42121=>"001000100",
42122=>"110110011",
42123=>"000110000",
42124=>"111011010",
42125=>"111110111",
42126=>"000000010",
42127=>"000001010",
42128=>"010000100",
42129=>"000000011",
42130=>"100110011",
42131=>"010111101",
42132=>"001001101",
42133=>"100000111",
42134=>"000001111",
42135=>"001001000",
42136=>"010100011",
42137=>"000000011",
42138=>"100100111",
42139=>"100010010",
42140=>"101100100",
42141=>"000110111",
42142=>"100110111",
42143=>"000011000",
42144=>"000011101",
42145=>"000000000",
42146=>"011000111",
42147=>"000000010",
42148=>"100000110",
42149=>"011011000",
42150=>"011101110",
42151=>"000100100",
42152=>"100000111",
42153=>"011011101",
42154=>"111101111",
42155=>"000100111",
42156=>"011001000",
42157=>"100100100",
42158=>"100101111",
42159=>"000010111",
42160=>"000111101",
42161=>"000001101",
42162=>"011001000",
42163=>"100000000",
42164=>"011011010",
42165=>"011010111",
42166=>"001000001",
42167=>"001100110",
42168=>"101010110",
42169=>"011011111",
42170=>"000011000",
42171=>"110110000",
42172=>"011001101",
42173=>"111110111",
42174=>"000000011",
42175=>"001111101",
42176=>"100111011",
42177=>"100000111",
42178=>"000111110",
42179=>"100101100",
42180=>"011000100",
42181=>"110110000",
42182=>"011001011",
42183=>"100011011",
42184=>"100000101",
42185=>"011011011",
42186=>"000000010",
42187=>"011111011",
42188=>"000010100",
42189=>"001000111",
42190=>"011011000",
42191=>"011011000",
42192=>"000101001",
42193=>"011101001",
42194=>"011011000",
42195=>"011001110",
42196=>"100110011",
42197=>"010111100",
42198=>"100111101",
42199=>"100000111",
42200=>"011100100",
42201=>"011001000",
42202=>"010001000",
42203=>"100100100",
42204=>"111110000",
42205=>"001011101",
42206=>"111000000",
42207=>"111101011",
42208=>"001111001",
42209=>"100110101",
42210=>"101001101",
42211=>"100010110",
42212=>"100100100",
42213=>"110011010",
42214=>"000111111",
42215=>"100000000",
42216=>"100011011",
42217=>"110110000",
42218=>"000000000",
42219=>"000000100",
42220=>"001011011",
42221=>"100111000",
42222=>"101001001",
42223=>"000000011",
42224=>"011011000",
42225=>"111101101",
42226=>"111011101",
42227=>"111000100",
42228=>"011111111",
42229=>"100100100",
42230=>"100000001",
42231=>"110110000",
42232=>"000000110",
42233=>"111001000",
42234=>"011001000",
42235=>"011000001",
42236=>"100100101",
42237=>"000100001",
42238=>"111011011",
42239=>"100110111",
42240=>"011010110",
42241=>"010011101",
42242=>"101000111",
42243=>"110111011",
42244=>"001001110",
42245=>"110000111",
42246=>"010111111",
42247=>"001111111",
42248=>"001101111",
42249=>"000000111",
42250=>"000100000",
42251=>"110101000",
42252=>"010000110",
42253=>"000000110",
42254=>"000000100",
42255=>"001011000",
42256=>"000110111",
42257=>"000000011",
42258=>"000000110",
42259=>"011010000",
42260=>"111011001",
42261=>"111101101",
42262=>"001011001",
42263=>"111111101",
42264=>"100000100",
42265=>"101101101",
42266=>"110101111",
42267=>"101101101",
42268=>"111010000",
42269=>"000000000",
42270=>"110010100",
42271=>"000000000",
42272=>"001101000",
42273=>"011111011",
42274=>"010101100",
42275=>"010110000",
42276=>"001110110",
42277=>"111010001",
42278=>"101000000",
42279=>"000001110",
42280=>"010011111",
42281=>"000001001",
42282=>"000000010",
42283=>"000111000",
42284=>"100111000",
42285=>"101001101",
42286=>"111011000",
42287=>"001011000",
42288=>"110010101",
42289=>"000110010",
42290=>"000100000",
42291=>"111101000",
42292=>"011000001",
42293=>"010001001",
42294=>"110110010",
42295=>"010011001",
42296=>"110010011",
42297=>"000000000",
42298=>"000000000",
42299=>"111101000",
42300=>"100000001",
42301=>"111000000",
42302=>"000000011",
42303=>"000000000",
42304=>"111101101",
42305=>"111011000",
42306=>"001100101",
42307=>"011010000",
42308=>"100010010",
42309=>"000010000",
42310=>"000101101",
42311=>"000000111",
42312=>"110111110",
42313=>"010010000",
42314=>"000001001",
42315=>"111100111",
42316=>"011000100",
42317=>"110111011",
42318=>"100101011",
42319=>"111111100",
42320=>"000111011",
42321=>"000111111",
42322=>"010010100",
42323=>"011001010",
42324=>"110001100",
42325=>"100000100",
42326=>"001011010",
42327=>"100000110",
42328=>"100110011",
42329=>"000011011",
42330=>"000000001",
42331=>"011011111",
42332=>"011000000",
42333=>"000100110",
42334=>"111010111",
42335=>"100110101",
42336=>"000000000",
42337=>"100010010",
42338=>"001000111",
42339=>"000010100",
42340=>"000001011",
42341=>"011000000",
42342=>"000011010",
42343=>"000010111",
42344=>"000000000",
42345=>"111000100",
42346=>"111010111",
42347=>"111110110",
42348=>"100111110",
42349=>"001011111",
42350=>"100101000",
42351=>"110111111",
42352=>"000101100",
42353=>"010100101",
42354=>"011011101",
42355=>"000000101",
42356=>"111100000",
42357=>"100000101",
42358=>"100111111",
42359=>"001001001",
42360=>"011000111",
42361=>"010000000",
42362=>"100101101",
42363=>"000100010",
42364=>"101001001",
42365=>"100100010",
42366=>"000000101",
42367=>"000000111",
42368=>"010111001",
42369=>"011001000",
42370=>"101011101",
42371=>"000101111",
42372=>"011000000",
42373=>"101100101",
42374=>"111010100",
42375=>"101100110",
42376=>"100110011",
42377=>"010011101",
42378=>"111111111",
42379=>"010111100",
42380=>"100101111",
42381=>"100000001",
42382=>"010010101",
42383=>"000100111",
42384=>"101011111",
42385=>"001010000",
42386=>"101101101",
42387=>"001111000",
42388=>"001100110",
42389=>"010101110",
42390=>"111111111",
42391=>"000110110",
42392=>"111110000",
42393=>"101111000",
42394=>"101011000",
42395=>"101000111",
42396=>"111100100",
42397=>"111111010",
42398=>"010010101",
42399=>"001111010",
42400=>"000001001",
42401=>"000010011",
42402=>"000001110",
42403=>"111111100",
42404=>"100001000",
42405=>"100001011",
42406=>"110110000",
42407=>"010111110",
42408=>"101011000",
42409=>"010111101",
42410=>"111001110",
42411=>"000100010",
42412=>"101111100",
42413=>"000011111",
42414=>"100110011",
42415=>"110101111",
42416=>"110000101",
42417=>"111001001",
42418=>"000010011",
42419=>"001001011",
42420=>"101111100",
42421=>"111011011",
42422=>"011101111",
42423=>"000000010",
42424=>"001000100",
42425=>"101101001",
42426=>"000010010",
42427=>"010000111",
42428=>"010000000",
42429=>"111001011",
42430=>"101100010",
42431=>"000000000",
42432=>"000010001",
42433=>"100000000",
42434=>"110010000",
42435=>"000011000",
42436=>"000001100",
42437=>"000100110",
42438=>"011010110",
42439=>"000110111",
42440=>"000000101",
42441=>"010000001",
42442=>"111111000",
42443=>"000001111",
42444=>"000100100",
42445=>"000100100",
42446=>"000001011",
42447=>"000100000",
42448=>"101010010",
42449=>"001011011",
42450=>"011111001",
42451=>"000101111",
42452=>"100000001",
42453=>"101111001",
42454=>"000000010",
42455=>"111111111",
42456=>"000000000",
42457=>"001010000",
42458=>"010110100",
42459=>"101000101",
42460=>"001101001",
42461=>"111010100",
42462=>"111101000",
42463=>"010000001",
42464=>"100000101",
42465=>"111000011",
42466=>"010000101",
42467=>"000010010",
42468=>"000000001",
42469=>"111111000",
42470=>"111001000",
42471=>"000110110",
42472=>"000000101",
42473=>"000011000",
42474=>"100111010",
42475=>"010101010",
42476=>"000000111",
42477=>"111010100",
42478=>"001000000",
42479=>"011100110",
42480=>"101100000",
42481=>"001001011",
42482=>"111011001",
42483=>"001110110",
42484=>"100110110",
42485=>"000000100",
42486=>"100000111",
42487=>"000000100",
42488=>"000111111",
42489=>"000110111",
42490=>"000111111",
42491=>"100001000",
42492=>"010100000",
42493=>"000000000",
42494=>"101011111",
42495=>"001010000",
42496=>"111111111",
42497=>"000010010",
42498=>"000000101",
42499=>"000110101",
42500=>"000001000",
42501=>"001000100",
42502=>"011111011",
42503=>"111111000",
42504=>"101000000",
42505=>"000000001",
42506=>"011011010",
42507=>"111010101",
42508=>"000000000",
42509=>"000000100",
42510=>"110100000",
42511=>"111111111",
42512=>"001000000",
42513=>"011111110",
42514=>"000111000",
42515=>"010010010",
42516=>"111111010",
42517=>"100100111",
42518=>"000011010",
42519=>"000111011",
42520=>"101100000",
42521=>"111011011",
42522=>"000101100",
42523=>"000000000",
42524=>"001111001",
42525=>"000011111",
42526=>"111101000",
42527=>"000000000",
42528=>"000100100",
42529=>"000000000",
42530=>"000000111",
42531=>"010001001",
42532=>"101111111",
42533=>"100101000",
42534=>"000010010",
42535=>"100010000",
42536=>"101111110",
42537=>"111111000",
42538=>"000000110",
42539=>"001100000",
42540=>"001111111",
42541=>"011110000",
42542=>"010000000",
42543=>"101000100",
42544=>"000011010",
42545=>"010101000",
42546=>"001101100",
42547=>"011111001",
42548=>"000111011",
42549=>"111111011",
42550=>"000011011",
42551=>"100111010",
42552=>"111100000",
42553=>"000111111",
42554=>"000000101",
42555=>"011011011",
42556=>"110010000",
42557=>"111111011",
42558=>"000000100",
42559=>"000111111",
42560=>"001011010",
42561=>"101010100",
42562=>"111000000",
42563=>"111101111",
42564=>"000000000",
42565=>"101101111",
42566=>"001111011",
42567=>"011011111",
42568=>"000000000",
42569=>"000101100",
42570=>"111111101",
42571=>"110111111",
42572=>"101111110",
42573=>"001111101",
42574=>"101001001",
42575=>"111000000",
42576=>"000000010",
42577=>"111111111",
42578=>"111011111",
42579=>"001111000",
42580=>"000000111",
42581=>"100111100",
42582=>"001111011",
42583=>"011000000",
42584=>"010011111",
42585=>"010111010",
42586=>"000111000",
42587=>"000111010",
42588=>"101101000",
42589=>"110000000",
42590=>"101111000",
42591=>"111101001",
42592=>"101000001",
42593=>"000000000",
42594=>"000000101",
42595=>"011111100",
42596=>"010000101",
42597=>"010010010",
42598=>"000000000",
42599=>"110111010",
42600=>"111111111",
42601=>"011011110",
42602=>"000000000",
42603=>"100111011",
42604=>"000001000",
42605=>"000111000",
42606=>"100000000",
42607=>"101100000",
42608=>"110110100",
42609=>"010111110",
42610=>"010010010",
42611=>"111100000",
42612=>"101111000",
42613=>"000000111",
42614=>"001011000",
42615=>"000000011",
42616=>"000111111",
42617=>"000000000",
42618=>"101011110",
42619=>"111100000",
42620=>"101101100",
42621=>"101001000",
42622=>"100000000",
42623=>"111100101",
42624=>"101100000",
42625=>"111111111",
42626=>"000000010",
42627=>"000000011",
42628=>"111101010",
42629=>"010010111",
42630=>"011111000",
42631=>"000000000",
42632=>"001011011",
42633=>"111111000",
42634=>"111100000",
42635=>"111110000",
42636=>"111100100",
42637=>"111111111",
42638=>"000111111",
42639=>"100000000",
42640=>"000110110",
42641=>"000011010",
42642=>"000000010",
42643=>"100011010",
42644=>"000011011",
42645=>"101000000",
42646=>"011011000",
42647=>"111111100",
42648=>"000000011",
42649=>"011111111",
42650=>"000011010",
42651=>"101000110",
42652=>"100111111",
42653=>"000001000",
42654=>"111010001",
42655=>"010111111",
42656=>"111000110",
42657=>"101111001",
42658=>"010101001",
42659=>"000011011",
42660=>"000111011",
42661=>"010010011",
42662=>"011101100",
42663=>"000111110",
42664=>"010000010",
42665=>"011000001",
42666=>"000000000",
42667=>"000000111",
42668=>"110000101",
42669=>"000000101",
42670=>"110111101",
42671=>"111000000",
42672=>"100100101",
42673=>"010010000",
42674=>"111111111",
42675=>"011110110",
42676=>"100111011",
42677=>"000011010",
42678=>"000000000",
42679=>"000000000",
42680=>"000011100",
42681=>"000000010",
42682=>"000000011",
42683=>"000111001",
42684=>"100011010",
42685=>"111111111",
42686=>"110100100",
42687=>"000111011",
42688=>"000000000",
42689=>"000111000",
42690=>"011111010",
42691=>"010001001",
42692=>"000111010",
42693=>"111101011",
42694=>"100010010",
42695=>"000101111",
42696=>"000010111",
42697=>"100111111",
42698=>"000010011",
42699=>"000011000",
42700=>"100101110",
42701=>"111111010",
42702=>"000011110",
42703=>"110100100",
42704=>"000111010",
42705=>"111111101",
42706=>"010000000",
42707=>"111111000",
42708=>"101000101",
42709=>"000001000",
42710=>"100000000",
42711=>"000111000",
42712=>"000011000",
42713=>"000000100",
42714=>"010111000",
42715=>"010000000",
42716=>"000111010",
42717=>"000100100",
42718=>"100000010",
42719=>"000000000",
42720=>"101000100",
42721=>"001000000",
42722=>"111111101",
42723=>"000010000",
42724=>"100000000",
42725=>"111011000",
42726=>"100111001",
42727=>"001110110",
42728=>"000001010",
42729=>"010111000",
42730=>"000111010",
42731=>"010000011",
42732=>"000000000",
42733=>"100011000",
42734=>"101101111",
42735=>"011000101",
42736=>"010111011",
42737=>"011101111",
42738=>"010000000",
42739=>"100111100",
42740=>"100101011",
42741=>"011010000",
42742=>"111000000",
42743=>"110000111",
42744=>"000111000",
42745=>"011110010",
42746=>"000011000",
42747=>"101110100",
42748=>"000111010",
42749=>"111111000",
42750=>"100111001",
42751=>"010111000",
42752=>"100001111",
42753=>"110100110",
42754=>"001011001",
42755=>"000011101",
42756=>"110111000",
42757=>"001011000",
42758=>"001000000",
42759=>"100000000",
42760=>"100110111",
42761=>"011011001",
42762=>"110100000",
42763=>"100010100",
42764=>"011011000",
42765=>"000001111",
42766=>"111000000",
42767=>"100111010",
42768=>"100010011",
42769=>"011011011",
42770=>"010010100",
42771=>"100100000",
42772=>"100100100",
42773=>"001011001",
42774=>"101100100",
42775=>"001001010",
42776=>"010011011",
42777=>"001101100",
42778=>"001011011",
42779=>"001101100",
42780=>"000110110",
42781=>"110100100",
42782=>"010011011",
42783=>"100100100",
42784=>"011010011",
42785=>"010011111",
42786=>"011001000",
42787=>"010110110",
42788=>"111000100",
42789=>"100101000",
42790=>"010011000",
42791=>"111011000",
42792=>"010100100",
42793=>"010110000",
42794=>"110010110",
42795=>"100100100",
42796=>"100100100",
42797=>"000011111",
42798=>"110111001",
42799=>"111100110",
42800=>"110110110",
42801=>"110110110",
42802=>"011011001",
42803=>"001011011",
42804=>"100100111",
42805=>"110100100",
42806=>"110100000",
42807=>"100100111",
42808=>"101011011",
42809=>"100000100",
42810=>"100100000",
42811=>"010000111",
42812=>"010000000",
42813=>"100100100",
42814=>"001011001",
42815=>"010011011",
42816=>"111011011",
42817=>"100010111",
42818=>"101001001",
42819=>"000011011",
42820=>"011001001",
42821=>"001011001",
42822=>"000010000",
42823=>"000000000",
42824=>"110100000",
42825=>"000110110",
42826=>"110011110",
42827=>"001001111",
42828=>"001001001",
42829=>"000000001",
42830=>"100001101",
42831=>"011100111",
42832=>"110000100",
42833=>"100100111",
42834=>"001011001",
42835=>"100100111",
42836=>"110100100",
42837=>"100100100",
42838=>"010000000",
42839=>"001011001",
42840=>"111011001",
42841=>"111110100",
42842=>"100100110",
42843=>"011010010",
42844=>"001001011",
42845=>"110100100",
42846=>"011011011",
42847=>"010110100",
42848=>"011011011",
42849=>"001010101",
42850=>"001011001",
42851=>"110000000",
42852=>"000000101",
42853=>"110100010",
42854=>"110100100",
42855=>"100100111",
42856=>"000101101",
42857=>"001011011",
42858=>"111011000",
42859=>"101111111",
42860=>"011011111",
42861=>"111011001",
42862=>"001001000",
42863=>"110100000",
42864=>"110101101",
42865=>"010011011",
42866=>"100100110",
42867=>"000011000",
42868=>"101111111",
42869=>"000011011",
42870=>"001111001",
42871=>"001001001",
42872=>"100010110",
42873=>"110000100",
42874=>"000001101",
42875=>"011011001",
42876=>"100101110",
42877=>"100000000",
42878=>"100100100",
42879=>"111111100",
42880=>"001011001",
42881=>"110010110",
42882=>"000011000",
42883=>"111011101",
42884=>"011001101",
42885=>"000101101",
42886=>"000100011",
42887=>"011011000",
42888=>"100100100",
42889=>"110111101",
42890=>"000100111",
42891=>"101011110",
42892=>"011100000",
42893=>"101111110",
42894=>"000011101",
42895=>"011001001",
42896=>"111101101",
42897=>"010010110",
42898=>"000010010",
42899=>"100100100",
42900=>"000000000",
42901=>"011011001",
42902=>"111101101",
42903=>"000001000",
42904=>"000100100",
42905=>"101101111",
42906=>"001001001",
42907=>"001001011",
42908=>"100111001",
42909=>"000001111",
42910=>"000011111",
42911=>"110110100",
42912=>"010110111",
42913=>"101111111",
42914=>"110101111",
42915=>"001001001",
42916=>"100001000",
42917=>"001001001",
42918=>"001111000",
42919=>"110101001",
42920=>"111001011",
42921=>"001000110",
42922=>"011011011",
42923=>"100010001",
42924=>"011100011",
42925=>"000010110",
42926=>"110100100",
42927=>"011111101",
42928=>"011011011",
42929=>"000100010",
42930=>"110000100",
42931=>"000011110",
42932=>"110000110",
42933=>"100100000",
42934=>"011011010",
42935=>"000110110",
42936=>"000100110",
42937=>"101101100",
42938=>"100110110",
42939=>"000000100",
42940=>"000110110",
42941=>"000001001",
42942=>"000010010",
42943=>"000111110",
42944=>"001111011",
42945=>"100001001",
42946=>"000011111",
42947=>"100100110",
42948=>"001011001",
42949=>"110111110",
42950=>"111011001",
42951=>"000010000",
42952=>"110101000",
42953=>"011000110",
42954=>"001111110",
42955=>"001011000",
42956=>"110100100",
42957=>"110100000",
42958=>"100000000",
42959=>"011011011",
42960=>"100100111",
42961=>"100100100",
42962=>"001101100",
42963=>"001100111",
42964=>"111011011",
42965=>"100100100",
42966=>"101111111",
42967=>"111011111",
42968=>"100100100",
42969=>"011110010",
42970=>"010000000",
42971=>"011011011",
42972=>"000000100",
42973=>"001011001",
42974=>"100000000",
42975=>"111011011",
42976=>"000010011",
42977=>"001011001",
42978=>"111101100",
42979=>"011111101",
42980=>"110110000",
42981=>"100100110",
42982=>"100110000",
42983=>"000100100",
42984=>"000011001",
42985=>"110110110",
42986=>"100100101",
42987=>"011011000",
42988=>"001011011",
42989=>"011010100",
42990=>"000000000",
42991=>"111011110",
42992=>"000110110",
42993=>"100001011",
42994=>"010011011",
42995=>"100000000",
42996=>"111110100",
42997=>"011011011",
42998=>"011011011",
42999=>"111000110",
43000=>"100001000",
43001=>"100111110",
43002=>"111111101",
43003=>"111011111",
43004=>"111110110",
43005=>"110011011",
43006=>"111110001",
43007=>"000010100",
43008=>"011001100",
43009=>"111101000",
43010=>"000010010",
43011=>"000001011",
43012=>"001011010",
43013=>"100001111",
43014=>"110111111",
43015=>"100010010",
43016=>"001101001",
43017=>"110000111",
43018=>"111111110",
43019=>"001111111",
43020=>"000110110",
43021=>"000000000",
43022=>"101011011",
43023=>"000000001",
43024=>"000010010",
43025=>"001001000",
43026=>"101001000",
43027=>"110001111",
43028=>"111000000",
43029=>"000010011",
43030=>"011101100",
43031=>"111001111",
43032=>"010000001",
43033=>"011001101",
43034=>"000000000",
43035=>"000110110",
43036=>"111101111",
43037=>"000000000",
43038=>"110100000",
43039=>"001111101",
43040=>"000111111",
43041=>"111000101",
43042=>"000000100",
43043=>"000000111",
43044=>"111111011",
43045=>"110000100",
43046=>"010111011",
43047=>"000000000",
43048=>"111111000",
43049=>"011000000",
43050=>"111011001",
43051=>"111101001",
43052=>"100000001",
43053=>"110000000",
43054=>"101100110",
43055=>"101000000",
43056=>"111010010",
43057=>"111101101",
43058=>"000000000",
43059=>"111001000",
43060=>"111111101",
43061=>"111111111",
43062=>"010110110",
43063=>"000000000",
43064=>"111010110",
43065=>"000111011",
43066=>"010000000",
43067=>"111100000",
43068=>"000001000",
43069=>"111101111",
43070=>"000010000",
43071=>"000011001",
43072=>"111001000",
43073=>"000100110",
43074=>"101101111",
43075=>"001111110",
43076=>"111101000",
43077=>"000010010",
43078=>"101011110",
43079=>"101000000",
43080=>"000000000",
43081=>"111101100",
43082=>"010010010",
43083=>"000100100",
43084=>"110000101",
43085=>"011111111",
43086=>"100111110",
43087=>"000010111",
43088=>"001111101",
43089=>"111111111",
43090=>"111111111",
43091=>"011001110",
43092=>"000111110",
43093=>"001001000",
43094=>"111011010",
43095=>"100010010",
43096=>"001111001",
43097=>"011111111",
43098=>"000111100",
43099=>"101101000",
43100=>"011101101",
43101=>"000111001",
43102=>"010111111",
43103=>"100110011",
43104=>"001101101",
43105=>"010010000",
43106=>"010111000",
43107=>"000010001",
43108=>"001101101",
43109=>"111001001",
43110=>"001000111",
43111=>"111001111",
43112=>"111000010",
43113=>"111000000",
43114=>"110011000",
43115=>"000000101",
43116=>"011011011",
43117=>"100001011",
43118=>"111111001",
43119=>"010100101",
43120=>"110100000",
43121=>"111000000",
43122=>"111011101",
43123=>"000000111",
43124=>"011111000",
43125=>"000000111",
43126=>"000000110",
43127=>"111111111",
43128=>"000011110",
43129=>"001101111",
43130=>"000000000",
43131=>"101010010",
43132=>"011101110",
43133=>"110100000",
43134=>"111101000",
43135=>"000111100",
43136=>"111101010",
43137=>"111010010",
43138=>"111111100",
43139=>"000001100",
43140=>"111110000",
43141=>"101110111",
43142=>"110000001",
43143=>"011111000",
43144=>"011101101",
43145=>"010001011",
43146=>"000000001",
43147=>"000000000",
43148=>"010111111",
43149=>"000110111",
43150=>"000111111",
43151=>"001000001",
43152=>"111101011",
43153=>"101101001",
43154=>"111101001",
43155=>"001011010",
43156=>"000001101",
43157=>"111010110",
43158=>"001111111",
43159=>"000001001",
43160=>"000110100",
43161=>"001000000",
43162=>"011111111",
43163=>"001010000",
43164=>"000001011",
43165=>"000111100",
43166=>"111000101",
43167=>"111001111",
43168=>"000000000",
43169=>"010010000",
43170=>"001111111",
43171=>"011011000",
43172=>"111111010",
43173=>"110100100",
43174=>"001110000",
43175=>"101101101",
43176=>"111011000",
43177=>"000010001",
43178=>"111111100",
43179=>"111111101",
43180=>"111000010",
43181=>"010111000",
43182=>"101101000",
43183=>"001111111",
43184=>"101000100",
43185=>"100000000",
43186=>"101101000",
43187=>"001100100",
43188=>"000011011",
43189=>"001100111",
43190=>"000110111",
43191=>"000111010",
43192=>"011001000",
43193=>"000100000",
43194=>"001101101",
43195=>"110111111",
43196=>"100000000",
43197=>"111110000",
43198=>"000100100",
43199=>"000000000",
43200=>"010000000",
43201=>"000001111",
43202=>"111000101",
43203=>"111101001",
43204=>"001111010",
43205=>"101000000",
43206=>"000100001",
43207=>"111000000",
43208=>"000000101",
43209=>"000101111",
43210=>"010100111",
43211=>"010111110",
43212=>"011001001",
43213=>"110000011",
43214=>"111101000",
43215=>"000111111",
43216=>"111111001",
43217=>"011010000",
43218=>"111111011",
43219=>"000000100",
43220=>"111111110",
43221=>"101110000",
43222=>"101111111",
43223=>"110000000",
43224=>"000111111",
43225=>"110111001",
43226=>"101001001",
43227=>"111000000",
43228=>"111011111",
43229=>"000001101",
43230=>"110011110",
43231=>"111000000",
43232=>"111110111",
43233=>"001010010",
43234=>"000111111",
43235=>"001101011",
43236=>"000000000",
43237=>"100111110",
43238=>"000000000",
43239=>"011011101",
43240=>"111100000",
43241=>"111000101",
43242=>"010110111",
43243=>"000010010",
43244=>"010111111",
43245=>"000111111",
43246=>"001011000",
43247=>"010001000",
43248=>"111111111",
43249=>"011000000",
43250=>"111110111",
43251=>"000111110",
43252=>"110100001",
43253=>"001101101",
43254=>"000001101",
43255=>"101001001",
43256=>"010111111",
43257=>"111110000",
43258=>"111111101",
43259=>"001001010",
43260=>"011111011",
43261=>"111111111",
43262=>"110101101",
43263=>"000000000",
43264=>"011100001",
43265=>"010110111",
43266=>"000000111",
43267=>"100001111",
43268=>"000001111",
43269=>"000000000",
43270=>"110111111",
43271=>"111111111",
43272=>"111000000",
43273=>"111000111",
43274=>"011011100",
43275=>"010111111",
43276=>"000000001",
43277=>"000000000",
43278=>"101001001",
43279=>"000000111",
43280=>"101100110",
43281=>"000000000",
43282=>"100100011",
43283=>"111111000",
43284=>"101101110",
43285=>"111111100",
43286=>"011011011",
43287=>"111111000",
43288=>"111111000",
43289=>"101101111",
43290=>"100101100",
43291=>"111111111",
43292=>"011111111",
43293=>"111110000",
43294=>"100000111",
43295=>"110000000",
43296=>"101111001",
43297=>"000000111",
43298=>"010010000",
43299=>"000000000",
43300=>"111110100",
43301=>"000000010",
43302=>"010011000",
43303=>"000000001",
43304=>"101000111",
43305=>"111111110",
43306=>"111001111",
43307=>"011000000",
43308=>"011110110",
43309=>"111101111",
43310=>"100000111",
43311=>"001000000",
43312=>"010000000",
43313=>"001001000",
43314=>"010010110",
43315=>"111111010",
43316=>"111111011",
43317=>"111111010",
43318=>"100000000",
43319=>"100111100",
43320=>"000011111",
43321=>"110100111",
43322=>"111111110",
43323=>"011110011",
43324=>"011001000",
43325=>"011111011",
43326=>"001000101",
43327=>"111011011",
43328=>"111000101",
43329=>"000111000",
43330=>"101001000",
43331=>"100100111",
43332=>"010111110",
43333=>"001000000",
43334=>"000000111",
43335=>"111000110",
43336=>"101111111",
43337=>"000101111",
43338=>"111111101",
43339=>"100100111",
43340=>"111110000",
43341=>"001111000",
43342=>"000100111",
43343=>"010111110",
43344=>"011000000",
43345=>"010010011",
43346=>"010111111",
43347=>"111111001",
43348=>"000000000",
43349=>"111100110",
43350=>"000000000",
43351=>"100100111",
43352=>"110111111",
43353=>"111011001",
43354=>"100001100",
43355=>"000000000",
43356=>"100101101",
43357=>"001011111",
43358=>"000000100",
43359=>"000000001",
43360=>"111111111",
43361=>"000010000",
43362=>"001001111",
43363=>"001111011",
43364=>"110011011",
43365=>"011000000",
43366=>"110111101",
43367=>"111111000",
43368=>"010111110",
43369=>"000111111",
43370=>"001111111",
43371=>"000101101",
43372=>"111111110",
43373=>"101111100",
43374=>"110100000",
43375=>"000000110",
43376=>"111001000",
43377=>"001111111",
43378=>"000000000",
43379=>"000000000",
43380=>"111011000",
43381=>"001101111",
43382=>"000000000",
43383=>"000010000",
43384=>"000000111",
43385=>"111111111",
43386=>"011001001",
43387=>"000000000",
43388=>"110000010",
43389=>"111001100",
43390=>"000000001",
43391=>"000000111",
43392=>"111111110",
43393=>"111111111",
43394=>"111111111",
43395=>"010110111",
43396=>"110110000",
43397=>"111111111",
43398=>"110011001",
43399=>"011010011",
43400=>"110100000",
43401=>"011011000",
43402=>"111010111",
43403=>"001000100",
43404=>"000000000",
43405=>"011111111",
43406=>"111100110",
43407=>"000001000",
43408=>"001001000",
43409=>"111111101",
43410=>"110111101",
43411=>"000000000",
43412=>"111100100",
43413=>"000000101",
43414=>"001101111",
43415=>"000110000",
43416=>"010010000",
43417=>"111111111",
43418=>"000010111",
43419=>"000000111",
43420=>"111111000",
43421=>"000101011",
43422=>"111101111",
43423=>"010011111",
43424=>"111111011",
43425=>"111111111",
43426=>"000000000",
43427=>"111111111",
43428=>"000111000",
43429=>"110110110",
43430=>"000000000",
43431=>"111101011",
43432=>"101000000",
43433=>"010110111",
43434=>"000000111",
43435=>"010000001",
43436=>"100110001",
43437=>"000010101",
43438=>"011001100",
43439=>"111000111",
43440=>"100100001",
43441=>"100010100",
43442=>"000000000",
43443=>"000100100",
43444=>"100010011",
43445=>"010000000",
43446=>"111111001",
43447=>"101000111",
43448=>"111010000",
43449=>"101001000",
43450=>"010000111",
43451=>"111110010",
43452=>"111111101",
43453=>"100000100",
43454=>"111001111",
43455=>"000011000",
43456=>"000000000",
43457=>"110111001",
43458=>"111111111",
43459=>"100100100",
43460=>"011011000",
43461=>"111001111",
43462=>"111111111",
43463=>"000000000",
43464=>"111111111",
43465=>"111110010",
43466=>"111111000",
43467=>"000111111",
43468=>"111111111",
43469=>"100000110",
43470=>"010111101",
43471=>"001100111",
43472=>"010011000",
43473=>"111011000",
43474=>"111111010",
43475=>"001101101",
43476=>"101111111",
43477=>"000000001",
43478=>"111101111",
43479=>"000000010",
43480=>"111011000",
43481=>"010110010",
43482=>"111111111",
43483=>"010011000",
43484=>"111000110",
43485=>"000000110",
43486=>"100010000",
43487=>"000001101",
43488=>"000000000",
43489=>"101000111",
43490=>"000000000",
43491=>"001111111",
43492=>"000011001",
43493=>"000000000",
43494=>"111111111",
43495=>"101100100",
43496=>"111111001",
43497=>"000111001",
43498=>"100010000",
43499=>"000000000",
43500=>"000011000",
43501=>"100111000",
43502=>"010010110",
43503=>"010000101",
43504=>"110111001",
43505=>"111101111",
43506=>"010000111",
43507=>"111111000",
43508=>"111111010",
43509=>"111111000",
43510=>"000000000",
43511=>"110011000",
43512=>"000000010",
43513=>"110010000",
43514=>"111111111",
43515=>"000100101",
43516=>"101100011",
43517=>"100000000",
43518=>"011111110",
43519=>"010000000",
43520=>"110100000",
43521=>"000001000",
43522=>"000000000",
43523=>"000010010",
43524=>"011011011",
43525=>"111111001",
43526=>"000010001",
43527=>"111111100",
43528=>"010111111",
43529=>"010111111",
43530=>"000011111",
43531=>"000000010",
43532=>"111111000",
43533=>"110010111",
43534=>"101111111",
43535=>"111111111",
43536=>"111111111",
43537=>"111111111",
43538=>"000101111",
43539=>"111000101",
43540=>"000101111",
43541=>"111111111",
43542=>"100110110",
43543=>"011110000",
43544=>"001001111",
43545=>"000000000",
43546=>"100111000",
43547=>"011111111",
43548=>"000001101",
43549=>"011010000",
43550=>"001000111",
43551=>"111011010",
43552=>"000000100",
43553=>"111111111",
43554=>"000000010",
43555=>"111111111",
43556=>"000000000",
43557=>"000011001",
43558=>"110111110",
43559=>"000000001",
43560=>"000000100",
43561=>"000111101",
43562=>"000000101",
43563=>"111101111",
43564=>"100110000",
43565=>"000000000",
43566=>"001000111",
43567=>"000000001",
43568=>"000111111",
43569=>"011010100",
43570=>"111111111",
43571=>"000000111",
43572=>"000000000",
43573=>"000100000",
43574=>"100111100",
43575=>"000000111",
43576=>"100111111",
43577=>"000000000",
43578=>"111000111",
43579=>"001101111",
43580=>"001001001",
43581=>"111111010",
43582=>"001101101",
43583=>"101100111",
43584=>"111111110",
43585=>"001111111",
43586=>"111111001",
43587=>"111111111",
43588=>"110111000",
43589=>"001000010",
43590=>"111111111",
43591=>"000000000",
43592=>"011000101",
43593=>"000010111",
43594=>"101110111",
43595=>"001000000",
43596=>"111111000",
43597=>"010000000",
43598=>"000000000",
43599=>"111001000",
43600=>"110111111",
43601=>"111010000",
43602=>"110100000",
43603=>"000100100",
43604=>"000000000",
43605=>"011111111",
43606=>"111011111",
43607=>"011111011",
43608=>"000110110",
43609=>"000000100",
43610=>"000011011",
43611=>"000000000",
43612=>"000111111",
43613=>"010001001",
43614=>"000000000",
43615=>"111111100",
43616=>"110110110",
43617=>"000000001",
43618=>"111110010",
43619=>"001000100",
43620=>"000000101",
43621=>"000000001",
43622=>"000000111",
43623=>"000111111",
43624=>"000001101",
43625=>"111000011",
43626=>"110000000",
43627=>"111111101",
43628=>"001101101",
43629=>"000000110",
43630=>"000001101",
43631=>"000000111",
43632=>"001001011",
43633=>"000000111",
43634=>"111011001",
43635=>"111110111",
43636=>"011000001",
43637=>"000000100",
43638=>"111111000",
43639=>"111111111",
43640=>"001010110",
43641=>"111111000",
43642=>"001001000",
43643=>"110010111",
43644=>"011001001",
43645=>"001000000",
43646=>"111111111",
43647=>"110111111",
43648=>"000111111",
43649=>"111110010",
43650=>"011100100",
43651=>"101111111",
43652=>"111000001",
43653=>"000000000",
43654=>"000110111",
43655=>"100000000",
43656=>"100010100",
43657=>"101000111",
43658=>"000000101",
43659=>"111001011",
43660=>"110111000",
43661=>"111101110",
43662=>"111101011",
43663=>"001001011",
43664=>"100100111",
43665=>"111111111",
43666=>"000111111",
43667=>"111001000",
43668=>"000001100",
43669=>"111111111",
43670=>"111111001",
43671=>"000111111",
43672=>"000000000",
43673=>"010010110",
43674=>"011110010",
43675=>"111111000",
43676=>"000000011",
43677=>"010010011",
43678=>"000111111",
43679=>"000000000",
43680=>"000110110",
43681=>"000011110",
43682=>"111111010",
43683=>"100000000",
43684=>"010111000",
43685=>"000000010",
43686=>"111111110",
43687=>"000001010",
43688=>"110010011",
43689=>"011101011",
43690=>"111111100",
43691=>"000101111",
43692=>"000000001",
43693=>"110011011",
43694=>"011011001",
43695=>"001000110",
43696=>"000000000",
43697=>"000000001",
43698=>"100110010",
43699=>"101101011",
43700=>"111000011",
43701=>"000000000",
43702=>"000000001",
43703=>"001000000",
43704=>"000100100",
43705=>"000000000",
43706=>"001000000",
43707=>"011000000",
43708=>"111000000",
43709=>"111111011",
43710=>"011011011",
43711=>"000000000",
43712=>"000000001",
43713=>"001101111",
43714=>"001001111",
43715=>"000000110",
43716=>"000000111",
43717=>"000000001",
43718=>"000000000",
43719=>"110010000",
43720=>"110000010",
43721=>"010111001",
43722=>"000000011",
43723=>"001000000",
43724=>"000000000",
43725=>"100001100",
43726=>"000101111",
43727=>"110111110",
43728=>"000000010",
43729=>"100100111",
43730=>"000000000",
43731=>"111000000",
43732=>"000001001",
43733=>"000100100",
43734=>"111111111",
43735=>"000000001",
43736=>"000000000",
43737=>"000000010",
43738=>"001001000",
43739=>"110110010",
43740=>"011111001",
43741=>"111111010",
43742=>"000000100",
43743=>"000000000",
43744=>"000111111",
43745=>"110111000",
43746=>"110111111",
43747=>"101100111",
43748=>"111001111",
43749=>"111111001",
43750=>"010010000",
43751=>"000111111",
43752=>"111110100",
43753=>"001000111",
43754=>"100010011",
43755=>"111110000",
43756=>"111111110",
43757=>"000001010",
43758=>"000000000",
43759=>"110111110",
43760=>"110000000",
43761=>"000001000",
43762=>"001001000",
43763=>"101100001",
43764=>"110000000",
43765=>"111111111",
43766=>"111111100",
43767=>"100000000",
43768=>"111111010",
43769=>"011000000",
43770=>"010011000",
43771=>"010000000",
43772=>"111111111",
43773=>"000111001",
43774=>"110000000",
43775=>"001000000",
43776=>"100100110",
43777=>"011100001",
43778=>"000010000",
43779=>"101000000",
43780=>"000111111",
43781=>"001101111",
43782=>"111000101",
43783=>"010011000",
43784=>"101001001",
43785=>"001000000",
43786=>"011000100",
43787=>"111100000",
43788=>"111001100",
43789=>"000110000",
43790=>"101100001",
43791=>"001111101",
43792=>"000000000",
43793=>"010001000",
43794=>"100000100",
43795=>"111111101",
43796=>"001001111",
43797=>"011010001",
43798=>"001111011",
43799=>"110111110",
43800=>"000000000",
43801=>"000001111",
43802=>"110110011",
43803=>"101000101",
43804=>"000101111",
43805=>"010000000",
43806=>"000101111",
43807=>"000000000",
43808=>"000111111",
43809=>"000010111",
43810=>"010010000",
43811=>"000000101",
43812=>"111110111",
43813=>"001001011",
43814=>"001111101",
43815=>"001010111",
43816=>"111111011",
43817=>"011101111",
43818=>"111100110",
43819=>"011010000",
43820=>"011100101",
43821=>"111111111",
43822=>"000110111",
43823=>"000011010",
43824=>"100001111",
43825=>"000011001",
43826=>"110000000",
43827=>"010001011",
43828=>"000000000",
43829=>"001010111",
43830=>"111111001",
43831=>"100000000",
43832=>"010100100",
43833=>"101000000",
43834=>"111101001",
43835=>"110011111",
43836=>"011001011",
43837=>"111110111",
43838=>"100000100",
43839=>"000110000",
43840=>"100101011",
43841=>"000101111",
43842=>"001100101",
43843=>"000100100",
43844=>"011101001",
43845=>"000111111",
43846=>"000111111",
43847=>"101000001",
43848=>"011111111",
43849=>"111100101",
43850=>"101101111",
43851=>"101000000",
43852=>"100000101",
43853=>"111101010",
43854=>"001110110",
43855=>"010010111",
43856=>"111101101",
43857=>"111111111",
43858=>"010000000",
43859=>"010001000",
43860=>"111000000",
43861=>"010110010",
43862=>"001011010",
43863=>"100000001",
43864=>"010000000",
43865=>"011001001",
43866=>"001010000",
43867=>"010111101",
43868=>"111000000",
43869=>"100110000",
43870=>"010011010",
43871=>"000000001",
43872=>"000000000",
43873=>"100100100",
43874=>"000000001",
43875=>"000110110",
43876=>"111001001",
43877=>"000111111",
43878=>"111101010",
43879=>"000000101",
43880=>"011011001",
43881=>"110111101",
43882=>"011111101",
43883=>"111101001",
43884=>"001000001",
43885=>"001000000",
43886=>"001101101",
43887=>"000101011",
43888=>"100110110",
43889=>"000000010",
43890=>"011001100",
43891=>"000000000",
43892=>"000001111",
43893=>"000001101",
43894=>"000000001",
43895=>"011101100",
43896=>"110111010",
43897=>"000100111",
43898=>"010010111",
43899=>"011000001",
43900=>"001001001",
43901=>"000001000",
43902=>"011011000",
43903=>"101001001",
43904=>"111000000",
43905=>"011011010",
43906=>"101111001",
43907=>"101111111",
43908=>"000101111",
43909=>"011000000",
43910=>"000101100",
43911=>"100000101",
43912=>"000011001",
43913=>"110100100",
43914=>"001000100",
43915=>"111101111",
43916=>"000111010",
43917=>"111001011",
43918=>"100101100",
43919=>"001000101",
43920=>"000100101",
43921=>"000110110",
43922=>"101111011",
43923=>"100100010",
43924=>"000010000",
43925=>"000000110",
43926=>"111100100",
43927=>"011001000",
43928=>"111101011",
43929=>"101111111",
43930=>"001100000",
43931=>"000000000",
43932=>"100100100",
43933=>"111000000",
43934=>"000101111",
43935=>"111100111",
43936=>"111011111",
43937=>"111111011",
43938=>"111101111",
43939=>"100000101",
43940=>"110011111",
43941=>"000000001",
43942=>"111101010",
43943=>"111101000",
43944=>"010010111",
43945=>"000000000",
43946=>"100111111",
43947=>"100000000",
43948=>"010011010",
43949=>"000000101",
43950=>"111111001",
43951=>"011101101",
43952=>"000001000",
43953=>"111110100",
43954=>"000100100",
43955=>"000000100",
43956=>"111111011",
43957=>"101000100",
43958=>"000000110",
43959=>"000001110",
43960=>"011100110",
43961=>"011000010",
43962=>"101001101",
43963=>"100000101",
43964=>"111111110",
43965=>"111011000",
43966=>"000101000",
43967=>"000110111",
43968=>"010111001",
43969=>"111000000",
43970=>"111101101",
43971=>"110100110",
43972=>"000000000",
43973=>"110111110",
43974=>"100000000",
43975=>"000000000",
43976=>"010000000",
43977=>"000011011",
43978=>"000000010",
43979=>"000000001",
43980=>"100000000",
43981=>"110100101",
43982=>"000000001",
43983=>"000001010",
43984=>"110111010",
43985=>"010011101",
43986=>"000000101",
43987=>"000011111",
43988=>"000010000",
43989=>"000001011",
43990=>"001000000",
43991=>"111101011",
43992=>"011011000",
43993=>"010010100",
43994=>"111111101",
43995=>"101000000",
43996=>"010011011",
43997=>"110100000",
43998=>"010000000",
43999=>"000111101",
44000=>"010000000",
44001=>"100000101",
44002=>"001111111",
44003=>"001100000",
44004=>"000010011",
44005=>"000000000",
44006=>"110000000",
44007=>"011111111",
44008=>"101000100",
44009=>"000011111",
44010=>"100100001",
44011=>"000000000",
44012=>"101000000",
44013=>"000010111",
44014=>"000000100",
44015=>"000000100",
44016=>"011010000",
44017=>"111111011",
44018=>"100000000",
44019=>"110110000",
44020=>"101001111",
44021=>"011000000",
44022=>"000000001",
44023=>"000011000",
44024=>"000111111",
44025=>"000111111",
44026=>"000010010",
44027=>"111111101",
44028=>"100100101",
44029=>"100000000",
44030=>"111110111",
44031=>"010000111",
44032=>"001100100",
44033=>"000000000",
44034=>"101000000",
44035=>"011111011",
44036=>"000011101",
44037=>"000000001",
44038=>"000111010",
44039=>"000011011",
44040=>"010001001",
44041=>"010010000",
44042=>"001001001",
44043=>"110110111",
44044=>"000000000",
44045=>"001000000",
44046=>"001011011",
44047=>"001111110",
44048=>"010000000",
44049=>"000000000",
44050=>"000000101",
44051=>"000000000",
44052=>"111111111",
44053=>"111011000",
44054=>"011011111",
44055=>"111010000",
44056=>"100100001",
44057=>"111010101",
44058=>"011001001",
44059=>"011010001",
44060=>"111000001",
44061=>"001101001",
44062=>"110000000",
44063=>"000001111",
44064=>"000000000",
44065=>"100011001",
44066=>"000111001",
44067=>"111111000",
44068=>"100101101",
44069=>"110000001",
44070=>"001001001",
44071=>"010000011",
44072=>"000000111",
44073=>"010010000",
44074=>"110010000",
44075=>"010000111",
44076=>"000000000",
44077=>"111000100",
44078=>"011010000",
44079=>"111111011",
44080=>"110000001",
44081=>"100111101",
44082=>"110000000",
44083=>"010000000",
44084=>"000000111",
44085=>"110011011",
44086=>"001011001",
44087=>"000011000",
44088=>"010000000",
44089=>"100000000",
44090=>"001110110",
44091=>"000000101",
44092=>"100110110",
44093=>"111101110",
44094=>"000010000",
44095=>"000110000",
44096=>"111011101",
44097=>"110110000",
44098=>"011111100",
44099=>"000100100",
44100=>"111100000",
44101=>"010010101",
44102=>"000000110",
44103=>"001010111",
44104=>"101011100",
44105=>"111111001",
44106=>"000000100",
44107=>"000110111",
44108=>"010000010",
44109=>"001111101",
44110=>"000101001",
44111=>"111100111",
44112=>"000001111",
44113=>"101000000",
44114=>"111010111",
44115=>"011000110",
44116=>"101110101",
44117=>"000000000",
44118=>"001100000",
44119=>"000111101",
44120=>"100100110",
44121=>"001111110",
44122=>"100101011",
44123=>"011011001",
44124=>"010010000",
44125=>"000001001",
44126=>"111010001",
44127=>"000001111",
44128=>"000111010",
44129=>"000001000",
44130=>"101101001",
44131=>"111111101",
44132=>"000110110",
44133=>"000001100",
44134=>"100110111",
44135=>"001111101",
44136=>"000000111",
44137=>"111010000",
44138=>"011011010",
44139=>"011010000",
44140=>"111000001",
44141=>"111001111",
44142=>"101000000",
44143=>"111000101",
44144=>"001111111",
44145=>"110110000",
44146=>"100100100",
44147=>"101111101",
44148=>"110111101",
44149=>"000000000",
44150=>"000000000",
44151=>"000100000",
44152=>"010010111",
44153=>"000010011",
44154=>"100000010",
44155=>"111011000",
44156=>"100110110",
44157=>"100000000",
44158=>"000001111",
44159=>"111111100",
44160=>"000000110",
44161=>"111000110",
44162=>"111111001",
44163=>"101101010",
44164=>"111000001",
44165=>"010000110",
44166=>"011011000",
44167=>"000110100",
44168=>"100111111",
44169=>"101011010",
44170=>"011110100",
44171=>"000000000",
44172=>"111111111",
44173=>"000011010",
44174=>"010011010",
44175=>"000001010",
44176=>"101100111",
44177=>"010000100",
44178=>"010111111",
44179=>"101101111",
44180=>"011100000",
44181=>"111011000",
44182=>"111010000",
44183=>"000001011",
44184=>"111011000",
44185=>"111011011",
44186=>"111101000",
44187=>"000000011",
44188=>"110001010",
44189=>"010011000",
44190=>"010011100",
44191=>"000111000",
44192=>"000001100",
44193=>"000101111",
44194=>"001001000",
44195=>"001101010",
44196=>"111001111",
44197=>"100110000",
44198=>"010110101",
44199=>"000001010",
44200=>"111010100",
44201=>"000111111",
44202=>"101000101",
44203=>"000101111",
44204=>"010001100",
44205=>"000111111",
44206=>"000001011",
44207=>"010010010",
44208=>"110110111",
44209=>"000001001",
44210=>"010000100",
44211=>"100110110",
44212=>"110111001",
44213=>"001011000",
44214=>"011111010",
44215=>"111010000",
44216=>"001011011",
44217=>"000001000",
44218=>"010011010",
44219=>"010010000",
44220=>"101101010",
44221=>"101011010",
44222=>"101111000",
44223=>"010000110",
44224=>"010110010",
44225=>"010010000",
44226=>"010010111",
44227=>"100101111",
44228=>"110100100",
44229=>"100110111",
44230=>"000000000",
44231=>"111010001",
44232=>"111011011",
44233=>"000000100",
44234=>"101111100",
44235=>"111011001",
44236=>"000001000",
44237=>"001011000",
44238=>"000100000",
44239=>"010001111",
44240=>"101010010",
44241=>"000101111",
44242=>"110100111",
44243=>"000101111",
44244=>"110110111",
44245=>"001101110",
44246=>"110010101",
44247=>"110010001",
44248=>"100000010",
44249=>"111010001",
44250=>"000100000",
44251=>"111000000",
44252=>"110111101",
44253=>"111101001",
44254=>"000011011",
44255=>"010010001",
44256=>"101111111",
44257=>"011111101",
44258=>"111000111",
44259=>"100111111",
44260=>"000111000",
44261=>"000101111",
44262=>"100111110",
44263=>"000100100",
44264=>"011010101",
44265=>"000000000",
44266=>"100100100",
44267=>"111111001",
44268=>"000000000",
44269=>"000000000",
44270=>"000000110",
44271=>"010001000",
44272=>"101001001",
44273=>"001011101",
44274=>"111011010",
44275=>"000011110",
44276=>"000001001",
44277=>"111101001",
44278=>"010110000",
44279=>"010000111",
44280=>"110000000",
44281=>"001010010",
44282=>"011110110",
44283=>"101111111",
44284=>"111111010",
44285=>"111111111",
44286=>"000111111",
44287=>"000011010",
44288=>"000000100",
44289=>"000001011",
44290=>"100100100",
44291=>"010100111",
44292=>"110000001",
44293=>"110100000",
44294=>"111011011",
44295=>"000011011",
44296=>"100100100",
44297=>"110001001",
44298=>"000011011",
44299=>"000000011",
44300=>"110100000",
44301=>"000100001",
44302=>"110101000",
44303=>"111110101",
44304=>"001011000",
44305=>"110001011",
44306=>"110100010",
44307=>"001001011",
44308=>"110110111",
44309=>"110110111",
44310=>"000010001",
44311=>"101011011",
44312=>"110000000",
44313=>"110010110",
44314=>"110000011",
44315=>"001001000",
44316=>"000000110",
44317=>"110000100",
44318=>"100100000",
44319=>"110100100",
44320=>"101101100",
44321=>"110010001",
44322=>"111100000",
44323=>"000000000",
44324=>"011111100",
44325=>"001101101",
44326=>"100001111",
44327=>"001011010",
44328=>"111010100",
44329=>"000000000",
44330=>"110010011",
44331=>"001000000",
44332=>"011110011",
44333=>"110100100",
44334=>"011110111",
44335=>"111010111",
44336=>"001111100",
44337=>"101110000",
44338=>"100000101",
44339=>"001110011",
44340=>"000011111",
44341=>"011011110",
44342=>"010100101",
44343=>"000011011",
44344=>"001100111",
44345=>"110100000",
44346=>"111100100",
44347=>"001011010",
44348=>"011110000",
44349=>"011111111",
44350=>"100001000",
44351=>"001000111",
44352=>"111000010",
44353=>"001011010",
44354=>"111011000",
44355=>"100001001",
44356=>"111100010",
44357=>"100000001",
44358=>"100110101",
44359=>"111101100",
44360=>"111111101",
44361=>"000100011",
44362=>"011001011",
44363=>"000001011",
44364=>"111100111",
44365=>"100101100",
44366=>"000011110",
44367=>"011110000",
44368=>"000000001",
44369=>"011111111",
44370=>"010111100",
44371=>"001001010",
44372=>"111100100",
44373=>"000111110",
44374=>"111110111",
44375=>"110100000",
44376=>"111011111",
44377=>"000000000",
44378=>"001001101",
44379=>"000001000",
44380=>"000001000",
44381=>"110100000",
44382=>"101011001",
44383=>"010100001",
44384=>"110110110",
44385=>"010100001",
44386=>"110100111",
44387=>"111111100",
44388=>"000110100",
44389=>"001000000",
44390=>"000100111",
44391=>"000000110",
44392=>"100100100",
44393=>"111100110",
44394=>"111011000",
44395=>"111011111",
44396=>"001000010",
44397=>"100001011",
44398=>"011000000",
44399=>"110111011",
44400=>"010111000",
44401=>"001000011",
44402=>"000001011",
44403=>"100100100",
44404=>"011011010",
44405=>"110100011",
44406=>"100100010",
44407=>"000100100",
44408=>"111101001",
44409=>"000011111",
44410=>"101011010",
44411=>"111110100",
44412=>"001011011",
44413=>"011110000",
44414=>"001011111",
44415=>"110100100",
44416=>"011010100",
44417=>"100100000",
44418=>"100011011",
44419=>"000111000",
44420=>"100100001",
44421=>"010100100",
44422=>"001001110",
44423=>"000001001",
44424=>"011111101",
44425=>"000000000",
44426=>"110011000",
44427=>"101011010",
44428=>"110001001",
44429=>"000100111",
44430=>"010111100",
44431=>"110000001",
44432=>"011010100",
44433=>"000001011",
44434=>"001011010",
44435=>"000011010",
44436=>"110001000",
44437=>"100000011",
44438=>"100111111",
44439=>"111110000",
44440=>"001011000",
44441=>"110100000",
44442=>"110110100",
44443=>"100100101",
44444=>"011001011",
44445=>"110100100",
44446=>"011001001",
44447=>"000000010",
44448=>"000000110",
44449=>"101100001",
44450=>"000101001",
44451=>"000101010",
44452=>"110010011",
44453=>"101101001",
44454=>"001010011",
44455=>"000000000",
44456=>"011001011",
44457=>"010110110",
44458=>"000100100",
44459=>"111000001",
44460=>"100100000",
44461=>"110100100",
44462=>"111111011",
44463=>"001011010",
44464=>"111000000",
44465=>"000001111",
44466=>"111110110",
44467=>"001010110",
44468=>"000110111",
44469=>"011111000",
44470=>"000001001",
44471=>"011001011",
44472=>"000001000",
44473=>"000001100",
44474=>"011100100",
44475=>"011110100",
44476=>"111111110",
44477=>"111011001",
44478=>"000000000",
44479=>"001010000",
44480=>"110100000",
44481=>"000001001",
44482=>"100110010",
44483=>"000000000",
44484=>"001010000",
44485=>"111110110",
44486=>"000111011",
44487=>"110100100",
44488=>"010110110",
44489=>"010000011",
44490=>"011101110",
44491=>"100111000",
44492=>"000001000",
44493=>"000001000",
44494=>"011001001",
44495=>"110101000",
44496=>"101000000",
44497=>"000000000",
44498=>"100110010",
44499=>"011110000",
44500=>"100100011",
44501=>"001010000",
44502=>"011100000",
44503=>"011111001",
44504=>"001011111",
44505=>"111000000",
44506=>"011110100",
44507=>"111100011",
44508=>"111011010",
44509=>"100100100",
44510=>"010100111",
44511=>"110000001",
44512=>"111010100",
44513=>"101100000",
44514=>"000011111",
44515=>"000111101",
44516=>"000010001",
44517=>"100001111",
44518=>"111101010",
44519=>"001001100",
44520=>"111111111",
44521=>"001011001",
44522=>"000001001",
44523=>"000100100",
44524=>"000010010",
44525=>"010010011",
44526=>"000000000",
44527=>"111000100",
44528=>"001000011",
44529=>"000000010",
44530=>"000011001",
44531=>"111111100",
44532=>"000011000",
44533=>"111010001",
44534=>"100000000",
44535=>"001000100",
44536=>"000011010",
44537=>"111111110",
44538=>"011100111",
44539=>"100110100",
44540=>"010111110",
44541=>"001011110",
44542=>"000000000",
44543=>"000011010",
44544=>"011000001",
44545=>"000110111",
44546=>"101101101",
44547=>"000000110",
44548=>"111000100",
44549=>"010000000",
44550=>"000010111",
44551=>"000000000",
44552=>"101111111",
44553=>"111101000",
44554=>"010100111",
44555=>"000100101",
44556=>"000011111",
44557=>"000100111",
44558=>"100101111",
44559=>"110111110",
44560=>"000000010",
44561=>"000000010",
44562=>"000000101",
44563=>"010010000",
44564=>"111101111",
44565=>"101010111",
44566=>"001111011",
44567=>"000000000",
44568=>"111000101",
44569=>"111100010",
44570=>"011101100",
44571=>"000000100",
44572=>"000001111",
44573=>"111010011",
44574=>"111101001",
44575=>"000010110",
44576=>"111101100",
44577=>"001101111",
44578=>"000010010",
44579=>"010111000",
44580=>"000110100",
44581=>"100000000",
44582=>"100101011",
44583=>"001000101",
44584=>"110010000",
44585=>"001110110",
44586=>"010000000",
44587=>"100001001",
44588=>"110010011",
44589=>"010111101",
44590=>"011111101",
44591=>"111011101",
44592=>"010001000",
44593=>"000110111",
44594=>"000011000",
44595=>"000111110",
44596=>"000000010",
44597=>"011011110",
44598=>"000100000",
44599=>"000110011",
44600=>"000000000",
44601=>"000100101",
44602=>"000111101",
44603=>"001000111",
44604=>"110000111",
44605=>"111101101",
44606=>"001000000",
44607=>"000000110",
44608=>"000000010",
44609=>"000000010",
44610=>"101101001",
44611=>"000000110",
44612=>"111101101",
44613=>"000010000",
44614=>"000000111",
44615=>"010000111",
44616=>"001101000",
44617=>"001001111",
44618=>"000000000",
44619=>"111111101",
44620=>"100101101",
44621=>"001101001",
44622=>"110000111",
44623=>"010000010",
44624=>"000101000",
44625=>"110000100",
44626=>"000000011",
44627=>"001001001",
44628=>"001010010",
44629=>"011010111",
44630=>"000011011",
44631=>"000000000",
44632=>"000111101",
44633=>"001011111",
44634=>"110100100",
44635=>"001011010",
44636=>"000101001",
44637=>"000001111",
44638=>"110111010",
44639=>"000000001",
44640=>"000101111",
44641=>"000000110",
44642=>"000001001",
44643=>"001000001",
44644=>"010000101",
44645=>"000100000",
44646=>"010111110",
44647=>"101111010",
44648=>"000001110",
44649=>"100000101",
44650=>"111111010",
44651=>"111100101",
44652=>"010101111",
44653=>"111010110",
44654=>"000000111",
44655=>"011011111",
44656=>"110111101",
44657=>"000000110",
44658=>"001101000",
44659=>"011011000",
44660=>"111110010",
44661=>"101001001",
44662=>"000010010",
44663=>"111111111",
44664=>"010000000",
44665=>"111100011",
44666=>"010110010",
44667=>"111111101",
44668=>"001001001",
44669=>"110100100",
44670=>"000000011",
44671=>"101111101",
44672=>"010000000",
44673=>"000010111",
44674=>"111000111",
44675=>"010000011",
44676=>"110000000",
44677=>"001000000",
44678=>"000000010",
44679=>"000000000",
44680=>"100110110",
44681=>"000101000",
44682=>"011001000",
44683=>"010000000",
44684=>"111110000",
44685=>"100000111",
44686=>"111100101",
44687=>"001000000",
44688=>"011000000",
44689=>"000000000",
44690=>"111001000",
44691=>"000000010",
44692=>"000000000",
44693=>"111000000",
44694=>"010111111",
44695=>"000011001",
44696=>"110010111",
44697=>"000001101",
44698=>"000010011",
44699=>"101000100",
44700=>"100101111",
44701=>"011001000",
44702=>"001100000",
44703=>"110100110",
44704=>"111111011",
44705=>"000011000",
44706=>"000000111",
44707=>"000000001",
44708=>"111100100",
44709=>"100110110",
44710=>"010110000",
44711=>"000000100",
44712=>"010000110",
44713=>"000111110",
44714=>"111111101",
44715=>"101000000",
44716=>"010010111",
44717=>"000000000",
44718=>"100100100",
44719=>"000000111",
44720=>"110100011",
44721=>"101001111",
44722=>"111101101",
44723=>"000000000",
44724=>"110011001",
44725=>"010011001",
44726=>"111101000",
44727=>"001000001",
44728=>"010000011",
44729=>"000100000",
44730=>"000000001",
44731=>"110110100",
44732=>"111000111",
44733=>"011111101",
44734=>"011011111",
44735=>"000111000",
44736=>"000001101",
44737=>"000000101",
44738=>"000101110",
44739=>"001110111",
44740=>"000000001",
44741=>"010110100",
44742=>"010010001",
44743=>"000000000",
44744=>"101111111",
44745=>"110111000",
44746=>"111101111",
44747=>"101010010",
44748=>"111100100",
44749=>"000100000",
44750=>"111111010",
44751=>"000010000",
44752=>"101000000",
44753=>"110110110",
44754=>"000010110",
44755=>"111010111",
44756=>"101000000",
44757=>"101111111",
44758=>"000101111",
44759=>"100101110",
44760=>"000010011",
44761=>"010010000",
44762=>"111011110",
44763=>"100000000",
44764=>"100011110",
44765=>"111011111",
44766=>"000001000",
44767=>"000010000",
44768=>"000000001",
44769=>"101101100",
44770=>"000000000",
44771=>"001011111",
44772=>"111001000",
44773=>"010101011",
44774=>"000000011",
44775=>"001001011",
44776=>"010000010",
44777=>"000000001",
44778=>"110011011",
44779=>"010010010",
44780=>"000010010",
44781=>"111011000",
44782=>"000000000",
44783=>"000000010",
44784=>"010010110",
44785=>"100010001",
44786=>"000001000",
44787=>"110010100",
44788=>"000110001",
44789=>"101101101",
44790=>"000000000",
44791=>"000111110",
44792=>"000000000",
44793=>"000100000",
44794=>"101101001",
44795=>"010011000",
44796=>"111111010",
44797=>"010000100",
44798=>"100000001",
44799=>"010000010",
44800=>"000010110",
44801=>"000000000",
44802=>"101101101",
44803=>"111011011",
44804=>"100000011",
44805=>"100000101",
44806=>"000110111",
44807=>"111010010",
44808=>"000010010",
44809=>"000111011",
44810=>"100000100",
44811=>"101000000",
44812=>"010100000",
44813=>"000000001",
44814=>"111110110",
44815=>"000011110",
44816=>"110110110",
44817=>"000000110",
44818=>"111000110",
44819=>"000010010",
44820=>"101111110",
44821=>"101001111",
44822=>"101001000",
44823=>"101110111",
44824=>"001000000",
44825=>"110010000",
44826=>"000010010",
44827=>"000110010",
44828=>"000101000",
44829=>"111000010",
44830=>"111101101",
44831=>"111001000",
44832=>"111000000",
44833=>"000010110",
44834=>"000001001",
44835=>"000000000",
44836=>"000111010",
44837=>"011111111",
44838=>"010110111",
44839=>"110111111",
44840=>"000010000",
44841=>"101010110",
44842=>"000110010",
44843=>"100001000",
44844=>"000011111",
44845=>"111111111",
44846=>"111010111",
44847=>"001001111",
44848=>"000101000",
44849=>"110000101",
44850=>"101110111",
44851=>"110111111",
44852=>"111000000",
44853=>"000000010",
44854=>"111000100",
44855=>"110100000",
44856=>"000010111",
44857=>"001100001",
44858=>"100011111",
44859=>"000000000",
44860=>"111111100",
44861=>"111011001",
44862=>"001101000",
44863=>"000010101",
44864=>"111000111",
44865=>"101111111",
44866=>"110000100",
44867=>"000000100",
44868=>"111000011",
44869=>"000101111",
44870=>"111100000",
44871=>"111010000",
44872=>"011110111",
44873=>"010010010",
44874=>"000100101",
44875=>"100011111",
44876=>"110000000",
44877=>"000111111",
44878=>"001100100",
44879=>"100110010",
44880=>"111001000",
44881=>"111011101",
44882=>"011010010",
44883=>"110011001",
44884=>"101000000",
44885=>"011111111",
44886=>"000111000",
44887=>"001001101",
44888=>"001111000",
44889=>"011010000",
44890=>"011000000",
44891=>"000110100",
44892=>"100111111",
44893=>"001011111",
44894=>"101011110",
44895=>"000000001",
44896=>"000000000",
44897=>"111011001",
44898=>"101001101",
44899=>"110100000",
44900=>"000111101",
44901=>"000111000",
44902=>"000110110",
44903=>"100000000",
44904=>"110011111",
44905=>"000010111",
44906=>"000001111",
44907=>"110110001",
44908=>"001110111",
44909=>"000110111",
44910=>"011000100",
44911=>"000111111",
44912=>"001111001",
44913=>"100110110",
44914=>"111101000",
44915=>"101011000",
44916=>"010010101",
44917=>"010001001",
44918=>"000000000",
44919=>"111011000",
44920=>"111000101",
44921=>"010010000",
44922=>"000000000",
44923=>"100111111",
44924=>"111110010",
44925=>"110110100",
44926=>"100111111",
44927=>"111000000",
44928=>"010110001",
44929=>"111100000",
44930=>"000110100",
44931=>"010111111",
44932=>"011110100",
44933=>"010010000",
44934=>"100110111",
44935=>"011000000",
44936=>"001110100",
44937=>"000100011",
44938=>"100111111",
44939=>"010001110",
44940=>"000001001",
44941=>"110111111",
44942=>"111010000",
44943=>"110001001",
44944=>"100011001",
44945=>"010111111",
44946=>"100111110",
44947=>"000000100",
44948=>"111000000",
44949=>"101101111",
44950=>"010011000",
44951=>"000010000",
44952=>"000100001",
44953=>"100000000",
44954=>"001111101",
44955=>"111100001",
44956=>"111111100",
44957=>"111001001",
44958=>"001010000",
44959=>"111101101",
44960=>"110111011",
44961=>"000111101",
44962=>"100010111",
44963=>"000111101",
44964=>"000111111",
44965=>"010110000",
44966=>"100001111",
44967=>"000010000",
44968=>"000000110",
44969=>"010010010",
44970=>"001101101",
44971=>"101000000",
44972=>"110101101",
44973=>"100000000",
44974=>"111110001",
44975=>"010001111",
44976=>"111000110",
44977=>"110001001",
44978=>"110111000",
44979=>"110101000",
44980=>"000011100",
44981=>"010111111",
44982=>"101111010",
44983=>"100110111",
44984=>"111111101",
44985=>"011000000",
44986=>"111010000",
44987=>"000000111",
44988=>"111111110",
44989=>"111101111",
44990=>"011011001",
44991=>"000110000",
44992=>"011001101",
44993=>"000000000",
44994=>"010110011",
44995=>"000110110",
44996=>"000010011",
44997=>"011000110",
44998=>"000000000",
44999=>"011111000",
45000=>"101111111",
45001=>"001001000",
45002=>"111111010",
45003=>"101000010",
45004=>"111010000",
45005=>"111110010",
45006=>"101000000",
45007=>"000000001",
45008=>"011101111",
45009=>"011111100",
45010=>"000000000",
45011=>"101000000",
45012=>"001001000",
45013=>"110000000",
45014=>"110010010",
45015=>"000000000",
45016=>"001000110",
45017=>"001111110",
45018=>"010110101",
45019=>"000000101",
45020=>"110010000",
45021=>"111101101",
45022=>"110000000",
45023=>"100000000",
45024=>"111000100",
45025=>"111100000",
45026=>"101101011",
45027=>"011111001",
45028=>"111000000",
45029=>"011000000",
45030=>"101110111",
45031=>"000110001",
45032=>"010111100",
45033=>"000000000",
45034=>"001001011",
45035=>"100001111",
45036=>"111100110",
45037=>"000000000",
45038=>"111100000",
45039=>"111100000",
45040=>"111000000",
45041=>"110000011",
45042=>"000000000",
45043=>"110110111",
45044=>"000111111",
45045=>"000000000",
45046=>"010000000",
45047=>"000010000",
45048=>"000100110",
45049=>"111110101",
45050=>"010110010",
45051=>"000000010",
45052=>"000110111",
45053=>"100000000",
45054=>"001111100",
45055=>"101111101",
45056=>"101000001",
45057=>"010111111",
45058=>"111111010",
45059=>"000000101",
45060=>"111000100",
45061=>"101001000",
45062=>"111100111",
45063=>"100101100",
45064=>"100101000",
45065=>"110100101",
45066=>"011001110",
45067=>"000100111",
45068=>"111111110",
45069=>"000110110",
45070=>"110000000",
45071=>"111001001",
45072=>"111111110",
45073=>"000000111",
45074=>"010000001",
45075=>"000000000",
45076=>"111000111",
45077=>"111111111",
45078=>"110111110",
45079=>"111000000",
45080=>"000001001",
45081=>"010100111",
45082=>"111111000",
45083=>"001000100",
45084=>"101110111",
45085=>"011111111",
45086=>"111010000",
45087=>"111011000",
45088=>"000100111",
45089=>"111010111",
45090=>"111010101",
45091=>"111001001",
45092=>"111100110",
45093=>"111001100",
45094=>"010010110",
45095=>"000010111",
45096=>"111110110",
45097=>"000110001",
45098=>"001111000",
45099=>"001000011",
45100=>"000000100",
45101=>"111100001",
45102=>"111111110",
45103=>"111001100",
45104=>"000010000",
45105=>"111010110",
45106=>"111111111",
45107=>"001000000",
45108=>"000110111",
45109=>"010010111",
45110=>"100000100",
45111=>"111000000",
45112=>"111001111",
45113=>"000000000",
45114=>"000101111",
45115=>"101000010",
45116=>"111110111",
45117=>"111000001",
45118=>"000000101",
45119=>"111001000",
45120=>"000111111",
45121=>"001000001",
45122=>"101101011",
45123=>"111110001",
45124=>"111111010",
45125=>"001000000",
45126=>"111101101",
45127=>"011000000",
45128=>"100111110",
45129=>"011111101",
45130=>"001011010",
45131=>"100111011",
45132=>"111111111",
45133=>"010001001",
45134=>"111011000",
45135=>"111001011",
45136=>"111111111",
45137=>"111110000",
45138=>"010111001",
45139=>"000000110",
45140=>"111000010",
45141=>"111011110",
45142=>"111100000",
45143=>"001000010",
45144=>"111111000",
45145=>"111011111",
45146=>"001111001",
45147=>"000101111",
45148=>"000000011",
45149=>"100111111",
45150=>"110000110",
45151=>"111011111",
45152=>"111101000",
45153=>"011111111",
45154=>"011101111",
45155=>"110100110",
45156=>"000011101",
45157=>"011001010",
45158=>"000000111",
45159=>"111110000",
45160=>"111111111",
45161=>"111000100",
45162=>"101111000",
45163=>"111001001",
45164=>"011000111",
45165=>"000100101",
45166=>"000111111",
45167=>"110111111",
45168=>"000010011",
45169=>"111010111",
45170=>"011000000",
45171=>"011000000",
45172=>"111111111",
45173=>"101000001",
45174=>"000111100",
45175=>"000101110",
45176=>"000111111",
45177=>"000000100",
45178=>"111111001",
45179=>"001000001",
45180=>"111011100",
45181=>"000000101",
45182=>"000000000",
45183=>"000100101",
45184=>"000000010",
45185=>"111111101",
45186=>"110101111",
45187=>"000010110",
45188=>"000000100",
45189=>"111011010",
45190=>"100100010",
45191=>"111010111",
45192=>"011001000",
45193=>"011000110",
45194=>"000000011",
45195=>"000000000",
45196=>"111111110",
45197=>"001000011",
45198=>"111000000",
45199=>"000010110",
45200=>"111110011",
45201=>"000001011",
45202=>"110110111",
45203=>"000001101",
45204=>"000000000",
45205=>"111111111",
45206=>"000000111",
45207=>"000111100",
45208=>"101100110",
45209=>"111111111",
45210=>"111000100",
45211=>"101000011",
45212=>"111110010",
45213=>"000100111",
45214=>"100111100",
45215=>"111000000",
45216=>"111110100",
45217=>"110001000",
45218=>"111111111",
45219=>"010010000",
45220=>"001000101",
45221=>"110010110",
45222=>"110111000",
45223=>"000000111",
45224=>"001000000",
45225=>"111111000",
45226=>"100101100",
45227=>"000010111",
45228=>"011000000",
45229=>"000000000",
45230=>"111111011",
45231=>"010011010",
45232=>"011001000",
45233=>"101111101",
45234=>"000000111",
45235=>"110011111",
45236=>"111101010",
45237=>"111101111",
45238=>"001100111",
45239=>"100101010",
45240=>"110111111",
45241=>"001001000",
45242=>"000100000",
45243=>"000000000",
45244=>"010000010",
45245=>"111111000",
45246=>"011001000",
45247=>"011000000",
45248=>"000110111",
45249=>"010000001",
45250=>"111011001",
45251=>"110110111",
45252=>"110111111",
45253=>"111010110",
45254=>"110010111",
45255=>"011011100",
45256=>"001101111",
45257=>"111000000",
45258=>"011111111",
45259=>"001000110",
45260=>"000100111",
45261=>"111110000",
45262=>"000111111",
45263=>"111000000",
45264=>"000000000",
45265=>"100011011",
45266=>"100100000",
45267=>"111001110",
45268=>"001101010",
45269=>"000011011",
45270=>"111111111",
45271=>"110111111",
45272=>"111010011",
45273=>"000010010",
45274=>"110000011",
45275=>"111000000",
45276=>"011110011",
45277=>"111111100",
45278=>"110111011",
45279=>"111110110",
45280=>"111010111",
45281=>"110101000",
45282=>"011000000",
45283=>"111000000",
45284=>"111111000",
45285=>"111000001",
45286=>"111001001",
45287=>"110111111",
45288=>"011111101",
45289=>"001000100",
45290=>"100110110",
45291=>"010100000",
45292=>"111001010",
45293=>"011000001",
45294=>"011000000",
45295=>"111001001",
45296=>"111000000",
45297=>"010001001",
45298=>"000000001",
45299=>"000100111",
45300=>"000100100",
45301=>"010100000",
45302=>"000001100",
45303=>"111001111",
45304=>"111111111",
45305=>"111111111",
45306=>"111111000",
45307=>"000011100",
45308=>"111000011",
45309=>"000000000",
45310=>"100100111",
45311=>"000000110",
45312=>"110100100",
45313=>"110111100",
45314=>"101001001",
45315=>"010001000",
45316=>"111101100",
45317=>"110000110",
45318=>"000010100",
45319=>"111011100",
45320=>"000000111",
45321=>"110000011",
45322=>"101000100",
45323=>"111010111",
45324=>"100001011",
45325=>"000000100",
45326=>"110111000",
45327=>"000000100",
45328=>"011010011",
45329=>"011011100",
45330=>"000000100",
45331=>"011100001",
45332=>"111110000",
45333=>"111111111",
45334=>"110110010",
45335=>"101111101",
45336=>"100000000",
45337=>"001010100",
45338=>"000111110",
45339=>"101111000",
45340=>"110100100",
45341=>"001001011",
45342=>"100110001",
45343=>"001000100",
45344=>"001110110",
45345=>"110010010",
45346=>"010100110",
45347=>"011110100",
45348=>"001000100",
45349=>"100100110",
45350=>"001001100",
45351=>"100001011",
45352=>"110111110",
45353=>"000110100",
45354=>"001111000",
45355=>"011010000",
45356=>"011111110",
45357=>"010000100",
45358=>"100110110",
45359=>"011111100",
45360=>"110111111",
45361=>"001001010",
45362=>"100101111",
45363=>"000011011",
45364=>"100100111",
45365=>"011111110",
45366=>"000110110",
45367=>"000001011",
45368=>"000010000",
45369=>"000000011",
45370=>"010000000",
45371=>"101001011",
45372=>"000001110",
45373=>"110000110",
45374=>"000010000",
45375=>"000111000",
45376=>"101000001",
45377=>"110110100",
45378=>"111001010",
45379=>"101100000",
45380=>"011000000",
45381=>"000000011",
45382=>"101010110",
45383=>"000011100",
45384=>"101111111",
45385=>"001010001",
45386=>"000000101",
45387=>"110101001",
45388=>"100100110",
45389=>"111110100",
45390=>"001001100",
45391=>"110110111",
45392=>"010110100",
45393=>"000111111",
45394=>"111100100",
45395=>"010010110",
45396=>"000001001",
45397=>"110010100",
45398=>"001100100",
45399=>"100111001",
45400=>"000000100",
45401=>"001111110",
45402=>"000100110",
45403=>"100110111",
45404=>"100001001",
45405=>"011011001",
45406=>"111000011",
45407=>"000111000",
45408=>"000000010",
45409=>"001011001",
45410=>"100000001",
45411=>"011111110",
45412=>"001100100",
45413=>"001101001",
45414=>"000110001",
45415=>"000100110",
45416=>"001001011",
45417=>"100110000",
45418=>"100000001",
45419=>"100000001",
45420=>"101111110",
45421=>"001010000",
45422=>"000000000",
45423=>"100111111",
45424=>"011001101",
45425=>"110001001",
45426=>"111110110",
45427=>"101001001",
45428=>"000000000",
45429=>"100000100",
45430=>"110011011",
45431=>"000100001",
45432=>"000110010",
45433=>"000000001",
45434=>"001000011",
45435=>"100101001",
45436=>"000001111",
45437=>"001110100",
45438=>"000000000",
45439=>"011111110",
45440=>"000110100",
45441=>"000000100",
45442=>"100000100",
45443=>"100110011",
45444=>"011001001",
45445=>"001100110",
45446=>"110100100",
45447=>"011001001",
45448=>"001101111",
45449=>"011100100",
45450=>"101100100",
45451=>"000001001",
45452=>"110001010",
45453=>"000100101",
45454=>"011111001",
45455=>"000000000",
45456=>"000010110",
45457=>"110110110",
45458=>"010100110",
45459=>"001011011",
45460=>"011011011",
45461=>"110001000",
45462=>"010111111",
45463=>"000110111",
45464=>"100100110",
45465=>"011100110",
45466=>"010100000",
45467=>"001001101",
45468=>"010100111",
45469=>"011011111",
45470=>"100110111",
45471=>"001000000",
45472=>"100111111",
45473=>"111011101",
45474=>"000110111",
45475=>"110110101",
45476=>"000000000",
45477=>"000000100",
45478=>"101101100",
45479=>"001110110",
45480=>"100001011",
45481=>"110100001",
45482=>"111001100",
45483=>"111110000",
45484=>"111001111",
45485=>"111101011",
45486=>"001110111",
45487=>"001000110",
45488=>"010011011",
45489=>"000011110",
45490=>"001111111",
45491=>"000000110",
45492=>"101011110",
45493=>"100011110",
45494=>"110100001",
45495=>"111111100",
45496=>"011011100",
45497=>"000001011",
45498=>"110110110",
45499=>"000000100",
45500=>"011100000",
45501=>"000100110",
45502=>"011011000",
45503=>"011011010",
45504=>"001000011",
45505=>"000000000",
45506=>"100100100",
45507=>"001111010",
45508=>"000010011",
45509=>"111001000",
45510=>"100111000",
45511=>"100010111",
45512=>"001001010",
45513=>"000111010",
45514=>"111011101",
45515=>"110000010",
45516=>"001000110",
45517=>"011011001",
45518=>"011011011",
45519=>"000011011",
45520=>"111110100",
45521=>"011111100",
45522=>"001000011",
45523=>"110100000",
45524=>"101000100",
45525=>"111111000",
45526=>"000010000",
45527=>"100111001",
45528=>"001001100",
45529=>"100000100",
45530=>"111101100",
45531=>"111000001",
45532=>"011011011",
45533=>"110010110",
45534=>"110101000",
45535=>"101101010",
45536=>"000000110",
45537=>"100001111",
45538=>"100100001",
45539=>"001111110",
45540=>"000000000",
45541=>"111110111",
45542=>"001011001",
45543=>"101101001",
45544=>"111000110",
45545=>"100100001",
45546=>"111100000",
45547=>"110001111",
45548=>"000000000",
45549=>"100000000",
45550=>"000000100",
45551=>"000000001",
45552=>"011001011",
45553=>"000010111",
45554=>"110110010",
45555=>"111001000",
45556=>"001001111",
45557=>"000000000",
45558=>"000000110",
45559=>"011011011",
45560=>"110011001",
45561=>"001110000",
45562=>"000000100",
45563=>"001001000",
45564=>"111110110",
45565=>"100011000",
45566=>"101001101",
45567=>"001110010",
45568=>"011001000",
45569=>"000111110",
45570=>"000000100",
45571=>"010110111",
45572=>"000101000",
45573=>"110010010",
45574=>"000001001",
45575=>"011111010",
45576=>"000111110",
45577=>"000000001",
45578=>"000000010",
45579=>"000100011",
45580=>"000000010",
45581=>"010010000",
45582=>"000000001",
45583=>"000001011",
45584=>"011111010",
45585=>"000000000",
45586=>"101101101",
45587=>"000011010",
45588=>"000001010",
45589=>"000011010",
45590=>"000111010",
45591=>"111111111",
45592=>"111000100",
45593=>"011111011",
45594=>"111111011",
45595=>"010111010",
45596=>"111001111",
45597=>"000000000",
45598=>"110100000",
45599=>"000000010",
45600=>"000000000",
45601=>"010111111",
45602=>"111101111",
45603=>"010111010",
45604=>"001111011",
45605=>"110111001",
45606=>"010010010",
45607=>"000110000",
45608=>"010011010",
45609=>"100110110",
45610=>"000011111",
45611=>"010000000",
45612=>"110111011",
45613=>"010100010",
45614=>"111010000",
45615=>"000101011",
45616=>"010111000",
45617=>"000101000",
45618=>"001001100",
45619=>"111000011",
45620=>"000000001",
45621=>"010111011",
45622=>"000011011",
45623=>"000000000",
45624=>"000010010",
45625=>"001000011",
45626=>"001001010",
45627=>"011000000",
45628=>"010110111",
45629=>"111111111",
45630=>"000000101",
45631=>"110110110",
45632=>"000101111",
45633=>"101001000",
45634=>"010010010",
45635=>"001110000",
45636=>"101111010",
45637=>"111010000",
45638=>"111001110",
45639=>"111101101",
45640=>"000001010",
45641=>"110111010",
45642=>"111010011",
45643=>"110000111",
45644=>"101100101",
45645=>"010011010",
45646=>"000001000",
45647=>"111010011",
45648=>"000010111",
45649=>"111111111",
45650=>"110011110",
45651=>"011111010",
45652=>"001000001",
45653=>"000100000",
45654=>"000111110",
45655=>"111111011",
45656=>"110011111",
45657=>"000010001",
45658=>"000010010",
45659=>"000111010",
45660=>"000001010",
45661=>"000001111",
45662=>"010010000",
45663=>"000010010",
45664=>"010110010",
45665=>"010111111",
45666=>"001000101",
45667=>"000011010",
45668=>"010010110",
45669=>"010011000",
45670=>"000000000",
45671=>"000010111",
45672=>"010011010",
45673=>"011001000",
45674=>"000010010",
45675=>"000010110",
45676=>"011011111",
45677=>"001001010",
45678=>"000000001",
45679=>"000011110",
45680=>"000111110",
45681=>"000010010",
45682=>"001100110",
45683=>"000000010",
45684=>"000010010",
45685=>"101000101",
45686=>"010111010",
45687=>"010110110",
45688=>"010010000",
45689=>"010011010",
45690=>"000001010",
45691=>"010111010",
45692=>"100100110",
45693=>"110111000",
45694=>"010111001",
45695=>"100111111",
45696=>"101101000",
45697=>"110100000",
45698=>"010010010",
45699=>"010000001",
45700=>"110010010",
45701=>"000101011",
45702=>"011100000",
45703=>"011111011",
45704=>"000111001",
45705=>"011011010",
45706=>"001010011",
45707=>"000100101",
45708=>"001010000",
45709=>"000000010",
45710=>"011111111",
45711=>"101000101",
45712=>"000001100",
45713=>"110111001",
45714=>"011000111",
45715=>"000110011",
45716=>"110111011",
45717=>"000000010",
45718=>"010111010",
45719=>"110111011",
45720=>"010111001",
45721=>"111111000",
45722=>"000010010",
45723=>"000000000",
45724=>"000000010",
45725=>"111010010",
45726=>"010111010",
45727=>"101000101",
45728=>"010010000",
45729=>"000010010",
45730=>"010110110",
45731=>"110111111",
45732=>"010000011",
45733=>"010011010",
45734=>"001011011",
45735=>"000000101",
45736=>"000111110",
45737=>"000111110",
45738=>"000000000",
45739=>"000000100",
45740=>"101000111",
45741=>"000000101",
45742=>"110110010",
45743=>"011010010",
45744=>"101101101",
45745=>"010011110",
45746=>"000101110",
45747=>"000000110",
45748=>"010111010",
45749=>"010111111",
45750=>"111111100",
45751=>"000000001",
45752=>"011010011",
45753=>"011010011",
45754=>"110000110",
45755=>"011010110",
45756=>"101001001",
45757=>"111111100",
45758=>"001011011",
45759=>"010000010",
45760=>"000011010",
45761=>"000000110",
45762=>"011111010",
45763=>"111111100",
45764=>"001001000",
45765=>"110110110",
45766=>"010010011",
45767=>"000000000",
45768=>"111111111",
45769=>"011111000",
45770=>"111001100",
45771=>"000010000",
45772=>"010011000",
45773=>"000000001",
45774=>"010000111",
45775=>"110110000",
45776=>"010100110",
45777=>"010111010",
45778=>"111011011",
45779=>"010011010",
45780=>"000001010",
45781=>"100111111",
45782=>"000000010",
45783=>"110101010",
45784=>"000011010",
45785=>"010001010",
45786=>"100000100",
45787=>"001000000",
45788=>"010110000",
45789=>"111011010",
45790=>"010010010",
45791=>"010000010",
45792=>"010000000",
45793=>"101000010",
45794=>"010111000",
45795=>"010111000",
45796=>"000000010",
45797=>"000010010",
45798=>"010000000",
45799=>"000111110",
45800=>"010010010",
45801=>"010111010",
45802=>"000000110",
45803=>"000000110",
45804=>"010010000",
45805=>"001111111",
45806=>"010101010",
45807=>"010000011",
45808=>"010010010",
45809=>"011101100",
45810=>"110111011",
45811=>"010011000",
45812=>"110010010",
45813=>"001000010",
45814=>"001000010",
45815=>"000101100",
45816=>"000010010",
45817=>"000010011",
45818=>"000000010",
45819=>"000001000",
45820=>"010111010",
45821=>"000000000",
45822=>"000101000",
45823=>"000000010",
45824=>"011010111",
45825=>"100111011",
45826=>"011100101",
45827=>"010111010",
45828=>"110110110",
45829=>"000010100",
45830=>"100101101",
45831=>"111111101",
45832=>"110010000",
45833=>"111101101",
45834=>"010001001",
45835=>"101111110",
45836=>"100000000",
45837=>"000000000",
45838=>"111110110",
45839=>"111111111",
45840=>"001101101",
45841=>"111110000",
45842=>"000011011",
45843=>"001000000",
45844=>"101101000",
45845=>"111111010",
45846=>"011111000",
45847=>"001101101",
45848=>"001001000",
45849=>"000000110",
45850=>"111111010",
45851=>"111100100",
45852=>"100100100",
45853=>"000111010",
45854=>"000111111",
45855=>"111111000",
45856=>"111101001",
45857=>"110111100",
45858=>"111111111",
45859=>"011111010",
45860=>"001111111",
45861=>"000001111",
45862=>"010011000",
45863=>"111101111",
45864=>"100101010",
45865=>"111111000",
45866=>"111111000",
45867=>"000010111",
45868=>"100110100",
45869=>"010011010",
45870=>"101111111",
45871=>"101000001",
45872=>"000100000",
45873=>"100110100",
45874=>"101010111",
45875=>"011000000",
45876=>"001101101",
45877=>"010101000",
45878=>"011011001",
45879=>"110010110",
45880=>"000000010",
45881=>"111111000",
45882=>"100001001",
45883=>"101001100",
45884=>"100111000",
45885=>"000011111",
45886=>"101000000",
45887=>"001000001",
45888=>"111111000",
45889=>"000010111",
45890=>"111110100",
45891=>"111111110",
45892=>"101000001",
45893=>"100010000",
45894=>"000000100",
45895=>"010111000",
45896=>"011111001",
45897=>"110100000",
45898=>"111111111",
45899=>"111001000",
45900=>"010111111",
45901=>"000111010",
45902=>"011011001",
45903=>"000000000",
45904=>"111000110",
45905=>"000111111",
45906=>"000111110",
45907=>"100111010",
45908=>"111101010",
45909=>"011011011",
45910=>"001011010",
45911=>"111101001",
45912=>"110111100",
45913=>"000110000",
45914=>"010011010",
45915=>"001101000",
45916=>"111111000",
45917=>"100100000",
45918=>"111101000",
45919=>"111111111",
45920=>"111111111",
45921=>"111111110",
45922=>"001000000",
45923=>"010010000",
45924=>"101111000",
45925=>"111100000",
45926=>"111111101",
45927=>"111001101",
45928=>"110101000",
45929=>"001111111",
45930=>"000010000",
45931=>"000011000",
45932=>"000010000",
45933=>"111111000",
45934=>"000011000",
45935=>"101000100",
45936=>"111111000",
45937=>"111011111",
45938=>"111111100",
45939=>"111111000",
45940=>"001111000",
45941=>"111011110",
45942=>"111001000",
45943=>"000111011",
45944=>"000000000",
45945=>"011101000",
45946=>"010000101",
45947=>"000111000",
45948=>"110010100",
45949=>"100011000",
45950=>"000000000",
45951=>"001000000",
45952=>"100000111",
45953=>"000000100",
45954=>"101111000",
45955=>"000111110",
45956=>"011111011",
45957=>"001010000",
45958=>"011110011",
45959=>"111101000",
45960=>"000111100",
45961=>"111101110",
45962=>"111101000",
45963=>"100111111",
45964=>"110111110",
45965=>"000000001",
45966=>"000101000",
45967=>"000010000",
45968=>"001011110",
45969=>"100101000",
45970=>"011011010",
45971=>"111000000",
45972=>"011111000",
45973=>"000101000",
45974=>"101101000",
45975=>"011011000",
45976=>"000000000",
45977=>"000000111",
45978=>"011001000",
45979=>"000000000",
45980=>"101111010",
45981=>"100100000",
45982=>"011011101",
45983=>"110100000",
45984=>"110110010",
45985=>"111101000",
45986=>"111001000",
45987=>"011111111",
45988=>"000110000",
45989=>"000111000",
45990=>"110111111",
45991=>"001100101",
45992=>"101000010",
45993=>"101010010",
45994=>"011011011",
45995=>"000010000",
45996=>"100000111",
45997=>"010011010",
45998=>"110011011",
45999=>"000100000",
46000=>"100100111",
46001=>"111111101",
46002=>"000010000",
46003=>"010011000",
46004=>"000100000",
46005=>"111000000",
46006=>"011001001",
46007=>"010000001",
46008=>"101110100",
46009=>"110110100",
46010=>"000000101",
46011=>"010101000",
46012=>"111011010",
46013=>"011000101",
46014=>"011110100",
46015=>"111101111",
46016=>"101111000",
46017=>"011011010",
46018=>"100111000",
46019=>"000100110",
46020=>"111101111",
46021=>"010011111",
46022=>"011111000",
46023=>"111111101",
46024=>"110111111",
46025=>"101100111",
46026=>"011010010",
46027=>"111111010",
46028=>"111110000",
46029=>"010000001",
46030=>"000000000",
46031=>"000000100",
46032=>"011001111",
46033=>"000000000",
46034=>"101000011",
46035=>"111111011",
46036=>"001111000",
46037=>"110000000",
46038=>"010110000",
46039=>"100101000",
46040=>"100100000",
46041=>"000000000",
46042=>"111001011",
46043=>"111000101",
46044=>"100111100",
46045=>"000001101",
46046=>"111011001",
46047=>"010100001",
46048=>"100100000",
46049=>"111101101",
46050=>"010011001",
46051=>"111111000",
46052=>"111101001",
46053=>"000111000",
46054=>"101000000",
46055=>"111110010",
46056=>"111010000",
46057=>"111111001",
46058=>"100100000",
46059=>"111011100",
46060=>"010000111",
46061=>"110111111",
46062=>"000111011",
46063=>"011011000",
46064=>"010111010",
46065=>"110101011",
46066=>"101111000",
46067=>"101111000",
46068=>"111111010",
46069=>"001001101",
46070=>"001010010",
46071=>"111011111",
46072=>"100100000",
46073=>"000110000",
46074=>"000111010",
46075=>"010100000",
46076=>"010010010",
46077=>"010010000",
46078=>"011011001",
46079=>"101010000",
46080=>"000000011",
46081=>"010000111",
46082=>"101101000",
46083=>"111101101",
46084=>"111111010",
46085=>"001001000",
46086=>"110010011",
46087=>"010010111",
46088=>"000000111",
46089=>"000111111",
46090=>"100011000",
46091=>"100111011",
46092=>"000111101",
46093=>"011011111",
46094=>"111010011",
46095=>"000100101",
46096=>"000010110",
46097=>"001111010",
46098=>"110111000",
46099=>"100100111",
46100=>"101010110",
46101=>"111111010",
46102=>"101100111",
46103=>"000000101",
46104=>"101101101",
46105=>"110110111",
46106=>"111000111",
46107=>"111011111",
46108=>"110101101",
46109=>"101111101",
46110=>"010100101",
46111=>"001100000",
46112=>"110010010",
46113=>"111011111",
46114=>"111001000",
46115=>"111101001",
46116=>"001011000",
46117=>"000000100",
46118=>"111000111",
46119=>"001111001",
46120=>"111000011",
46121=>"111010010",
46122=>"111001111",
46123=>"011011111",
46124=>"111001001",
46125=>"101001101",
46126=>"111111000",
46127=>"000000000",
46128=>"000000000",
46129=>"111101101",
46130=>"101100100",
46131=>"111000000",
46132=>"000000111",
46133=>"101101111",
46134=>"000100110",
46135=>"000111111",
46136=>"000111101",
46137=>"011101100",
46138=>"010110000",
46139=>"110000000",
46140=>"110001001",
46141=>"000110011",
46142=>"000101101",
46143=>"011010001",
46144=>"000000111",
46145=>"010110111",
46146=>"001010101",
46147=>"000100101",
46148=>"000000000",
46149=>"000001101",
46150=>"110010101",
46151=>"001100011",
46152=>"000000101",
46153=>"111000000",
46154=>"000010001",
46155=>"000011111",
46156=>"001111010",
46157=>"101111010",
46158=>"001010010",
46159=>"001110000",
46160=>"111010010",
46161=>"101000011",
46162=>"011000010",
46163=>"000001011",
46164=>"000111111",
46165=>"000000101",
46166=>"011001011",
46167=>"101111111",
46168=>"110110000",
46169=>"110110110",
46170=>"011000000",
46171=>"110110000",
46172=>"010110111",
46173=>"011001001",
46174=>"100000101",
46175=>"000001101",
46176=>"010010111",
46177=>"100110010",
46178=>"000011111",
46179=>"110100000",
46180=>"111111000",
46181=>"111011111",
46182=>"010000000",
46183=>"111111100",
46184=>"010111101",
46185=>"101100000",
46186=>"000010010",
46187=>"010011111",
46188=>"010111000",
46189=>"111111000",
46190=>"000001000",
46191=>"000010101",
46192=>"110110010",
46193=>"000110000",
46194=>"000000011",
46195=>"111101101",
46196=>"000000010",
46197=>"000001011",
46198=>"111001111",
46199=>"000111111",
46200=>"000001001",
46201=>"010010101",
46202=>"110000000",
46203=>"101101000",
46204=>"001111111",
46205=>"110100100",
46206=>"010111111",
46207=>"111011000",
46208=>"000000001",
46209=>"000101100",
46210=>"111100101",
46211=>"111111000",
46212=>"000010010",
46213=>"010000100",
46214=>"001000101",
46215=>"011000001",
46216=>"111010000",
46217=>"111000000",
46218=>"110110111",
46219=>"000000001",
46220=>"111001000",
46221=>"000101100",
46222=>"010000101",
46223=>"010000110",
46224=>"011011011",
46225=>"000100010",
46226=>"001001000",
46227=>"000011111",
46228=>"111000000",
46229=>"101101101",
46230=>"110000101",
46231=>"100000011",
46232=>"100011101",
46233=>"101001110",
46234=>"101100010",
46235=>"010101100",
46236=>"001101111",
46237=>"110111010",
46238=>"001100000",
46239=>"100011111",
46240=>"001000101",
46241=>"001001111",
46242=>"111011101",
46243=>"111111000",
46244=>"110110000",
46245=>"010011001",
46246=>"101001001",
46247=>"000010111",
46248=>"100111111",
46249=>"001000010",
46250=>"101000010",
46251=>"001001010",
46252=>"011000101",
46253=>"011110010",
46254=>"001111011",
46255=>"111111101",
46256=>"010001001",
46257=>"111011001",
46258=>"101111111",
46259=>"001011101",
46260=>"111111101",
46261=>"111111101",
46262=>"100000100",
46263=>"101000011",
46264=>"011100100",
46265=>"110010110",
46266=>"000000001",
46267=>"000111100",
46268=>"111100000",
46269=>"110111111",
46270=>"000111011",
46271=>"111111101",
46272=>"000010000",
46273=>"000000001",
46274=>"000001111",
46275=>"111111001",
46276=>"000000000",
46277=>"001001000",
46278=>"000100110",
46279=>"001000100",
46280=>"111000000",
46281=>"001001111",
46282=>"100011101",
46283=>"101001111",
46284=>"000100101",
46285=>"100111111",
46286=>"100111111",
46287=>"000111000",
46288=>"111111010",
46289=>"011010000",
46290=>"011111111",
46291=>"000000000",
46292=>"100000010",
46293=>"110100100",
46294=>"101111000",
46295=>"011011111",
46296=>"000100101",
46297=>"000000110",
46298=>"111010101",
46299=>"111000000",
46300=>"000000000",
46301=>"001100000",
46302=>"100110101",
46303=>"001000111",
46304=>"011111111",
46305=>"101101000",
46306=>"111000000",
46307=>"111011100",
46308=>"000001010",
46309=>"000000000",
46310=>"110011111",
46311=>"010111111",
46312=>"000010000",
46313=>"111100000",
46314=>"000010010",
46315=>"010101111",
46316=>"000010111",
46317=>"000000000",
46318=>"100010010",
46319=>"000000000",
46320=>"010100100",
46321=>"100100001",
46322=>"100111001",
46323=>"110000001",
46324=>"000000111",
46325=>"111000000",
46326=>"000100001",
46327=>"111111001",
46328=>"000001111",
46329=>"000100100",
46330=>"111110011",
46331=>"011110101",
46332=>"000010110",
46333=>"110101001",
46334=>"011000101",
46335=>"011111111",
46336=>"101000000",
46337=>"000000111",
46338=>"000000000",
46339=>"001101111",
46340=>"110001010",
46341=>"001001000",
46342=>"010100100",
46343=>"000111111",
46344=>"111001001",
46345=>"111000000",
46346=>"000000100",
46347=>"010000101",
46348=>"010010111",
46349=>"111000111",
46350=>"001010010",
46351=>"000000000",
46352=>"000001000",
46353=>"101000101",
46354=>"000110111",
46355=>"111000100",
46356=>"100000110",
46357=>"000010010",
46358=>"000101111",
46359=>"010000000",
46360=>"101000001",
46361=>"000000000",
46362=>"000000100",
46363=>"110111110",
46364=>"110111001",
46365=>"111000001",
46366=>"101110011",
46367=>"111101111",
46368=>"000000000",
46369=>"000000111",
46370=>"100101100",
46371=>"000101111",
46372=>"001001000",
46373=>"010110001",
46374=>"000111010",
46375=>"010111111",
46376=>"111000000",
46377=>"000111111",
46378=>"000011000",
46379=>"100000000",
46380=>"000111111",
46381=>"011111000",
46382=>"111010111",
46383=>"101110001",
46384=>"001111001",
46385=>"111010000",
46386=>"100100110",
46387=>"111111101",
46388=>"000000101",
46389=>"101101001",
46390=>"100100001",
46391=>"101111001",
46392=>"000110000",
46393=>"101001111",
46394=>"111101111",
46395=>"101111010",
46396=>"000111110",
46397=>"010111111",
46398=>"101100100",
46399=>"011001111",
46400=>"101000010",
46401=>"110010111",
46402=>"100111111",
46403=>"000000000",
46404=>"011000000",
46405=>"110001000",
46406=>"110000001",
46407=>"100110101",
46408=>"000111111",
46409=>"010000110",
46410=>"101101101",
46411=>"111111011",
46412=>"101110010",
46413=>"110100000",
46414=>"010011100",
46415=>"111000000",
46416=>"101101101",
46417=>"010111111",
46418=>"010010111",
46419=>"110010110",
46420=>"011000110",
46421=>"001100100",
46422=>"100111011",
46423=>"001000100",
46424=>"001101111",
46425=>"110110000",
46426=>"000110111",
46427=>"111100100",
46428=>"000100111",
46429=>"010000000",
46430=>"111111000",
46431=>"100100000",
46432=>"000110111",
46433=>"010000000",
46434=>"111111110",
46435=>"001111101",
46436=>"000100010",
46437=>"010110000",
46438=>"100000000",
46439=>"100011000",
46440=>"001000010",
46441=>"011100000",
46442=>"111111000",
46443=>"000110110",
46444=>"000110110",
46445=>"000000010",
46446=>"111110111",
46447=>"111010000",
46448=>"101111010",
46449=>"010010010",
46450=>"001001100",
46451=>"101101001",
46452=>"000011010",
46453=>"111001000",
46454=>"110100111",
46455=>"000010000",
46456=>"011111110",
46457=>"110010000",
46458=>"110001001",
46459=>"000000000",
46460=>"101000100",
46461=>"111100100",
46462=>"111000110",
46463=>"111000000",
46464=>"000000000",
46465=>"000000010",
46466=>"111101000",
46467=>"110010101",
46468=>"010000111",
46469=>"111101001",
46470=>"110111110",
46471=>"000000000",
46472=>"000110000",
46473=>"000111010",
46474=>"010000000",
46475=>"111101000",
46476=>"111001000",
46477=>"000000001",
46478=>"110010000",
46479=>"001001000",
46480=>"010111001",
46481=>"000000010",
46482=>"000101110",
46483=>"110000110",
46484=>"111111010",
46485=>"001000000",
46486=>"000111111",
46487=>"010010010",
46488=>"010111101",
46489=>"101111111",
46490=>"111000000",
46491=>"000100010",
46492=>"010101000",
46493=>"001101000",
46494=>"101101000",
46495=>"000111110",
46496=>"100001011",
46497=>"110100001",
46498=>"110000010",
46499=>"000101110",
46500=>"111011110",
46501=>"001001000",
46502=>"011111010",
46503=>"011110111",
46504=>"111000110",
46505=>"000000111",
46506=>"111000111",
46507=>"111110101",
46508=>"111111010",
46509=>"111100000",
46510=>"100101101",
46511=>"010001000",
46512=>"010110111",
46513=>"011011000",
46514=>"110000000",
46515=>"100011000",
46516=>"111000001",
46517=>"100111111",
46518=>"000000100",
46519=>"111000000",
46520=>"011111111",
46521=>"000010100",
46522=>"111011000",
46523=>"011111000",
46524=>"100110011",
46525=>"100000110",
46526=>"100000100",
46527=>"000000010",
46528=>"111000000",
46529=>"111000000",
46530=>"000110011",
46531=>"100000000",
46532=>"000110011",
46533=>"011111100",
46534=>"000000111",
46535=>"000110100",
46536=>"010010000",
46537=>"000110010",
46538=>"000001000",
46539=>"100000000",
46540=>"111101000",
46541=>"000100000",
46542=>"111100000",
46543=>"011011000",
46544=>"111000101",
46545=>"001111111",
46546=>"011111010",
46547=>"111101110",
46548=>"010010000",
46549=>"100100101",
46550=>"000000111",
46551=>"000111111",
46552=>"001111000",
46553=>"001000000",
46554=>"011100011",
46555=>"111000000",
46556=>"100111011",
46557=>"000000000",
46558=>"000001101",
46559=>"101000010",
46560=>"110011000",
46561=>"011001000",
46562=>"111111101",
46563=>"000001100",
46564=>"000001000",
46565=>"010000000",
46566=>"111000110",
46567=>"001111101",
46568=>"100111111",
46569=>"100000111",
46570=>"111001000",
46571=>"111000010",
46572=>"000111111",
46573=>"101001000",
46574=>"000000010",
46575=>"010100100",
46576=>"111101111",
46577=>"100011000",
46578=>"111111010",
46579=>"111111111",
46580=>"011110111",
46581=>"100000101",
46582=>"011001000",
46583=>"000111100",
46584=>"111000000",
46585=>"000001000",
46586=>"111101101",
46587=>"111111100",
46588=>"100111111",
46589=>"001000000",
46590=>"111000000",
46591=>"000110110",
46592=>"011011010",
46593=>"000000110",
46594=>"000000000",
46595=>"111111000",
46596=>"100000100",
46597=>"010110000",
46598=>"110010111",
46599=>"000111111",
46600=>"111101001",
46601=>"101101111",
46602=>"100000000",
46603=>"111111011",
46604=>"010010011",
46605=>"101101111",
46606=>"110101011",
46607=>"000000011",
46608=>"100000000",
46609=>"111111100",
46610=>"110110000",
46611=>"010000101",
46612=>"111111111",
46613=>"000000000",
46614=>"011011011",
46615=>"111110111",
46616=>"000110100",
46617=>"000000001",
46618=>"000000000",
46619=>"111111100",
46620=>"111111110",
46621=>"011101000",
46622=>"110100000",
46623=>"111111011",
46624=>"000010010",
46625=>"010011110",
46626=>"100110101",
46627=>"010111010",
46628=>"110111000",
46629=>"110100000",
46630=>"111110110",
46631=>"111010000",
46632=>"101000111",
46633=>"111111000",
46634=>"111011110",
46635=>"111111110",
46636=>"110111000",
46637=>"110010000",
46638=>"010110111",
46639=>"001000000",
46640=>"101000100",
46641=>"110100111",
46642=>"110100111",
46643=>"111011011",
46644=>"111110001",
46645=>"111111111",
46646=>"111111110",
46647=>"110000011",
46648=>"111110111",
46649=>"111000000",
46650=>"101000100",
46651=>"111111010",
46652=>"100100111",
46653=>"110111111",
46654=>"101000111",
46655=>"111101110",
46656=>"111011111",
46657=>"111000000",
46658=>"110110100",
46659=>"100100100",
46660=>"111010010",
46661=>"010000000",
46662=>"000100111",
46663=>"110110101",
46664=>"000110110",
46665=>"001001110",
46666=>"000000011",
46667=>"000000000",
46668=>"000000000",
46669=>"000111111",
46670=>"010000000",
46671=>"110111011",
46672=>"111111111",
46673=>"000111111",
46674=>"000000010",
46675=>"011001000",
46676=>"001000000",
46677=>"100010000",
46678=>"001001101",
46679=>"000000000",
46680=>"000101111",
46681=>"111111011",
46682=>"111111110",
46683=>"001000000",
46684=>"000000000",
46685=>"011001111",
46686=>"111111010",
46687=>"001111010",
46688=>"001001110",
46689=>"001100110",
46690=>"000000001",
46691=>"100111111",
46692=>"101110000",
46693=>"000000101",
46694=>"000100101",
46695=>"011011000",
46696=>"000110100",
46697=>"110001000",
46698=>"110000110",
46699=>"111000000",
46700=>"111000000",
46701=>"100110111",
46702=>"000000011",
46703=>"000001111",
46704=>"101100000",
46705=>"111111000",
46706=>"111111111",
46707=>"000000000",
46708=>"111000000",
46709=>"000000000",
46710=>"000000101",
46711=>"111111110",
46712=>"001000111",
46713=>"110101100",
46714=>"010010111",
46715=>"000110111",
46716=>"100110011",
46717=>"100100000",
46718=>"111101110",
46719=>"000001101",
46720=>"010000000",
46721=>"100100100",
46722=>"000000100",
46723=>"010000100",
46724=>"111111111",
46725=>"100000001",
46726=>"111011001",
46727=>"001011011",
46728=>"011011111",
46729=>"000000000",
46730=>"000000000",
46731=>"111000000",
46732=>"000000000",
46733=>"000011111",
46734=>"111111111",
46735=>"001000001",
46736=>"101111001",
46737=>"111111000",
46738=>"000000110",
46739=>"000000000",
46740=>"000101111",
46741=>"111111010",
46742=>"000000000",
46743=>"000110000",
46744=>"010010100",
46745=>"111111111",
46746=>"000111110",
46747=>"000000000",
46748=>"110110000",
46749=>"000111111",
46750=>"110010010",
46751=>"001001101",
46752=>"000111001",
46753=>"111110010",
46754=>"111110000",
46755=>"111101101",
46756=>"111111111",
46757=>"110100000",
46758=>"111110111",
46759=>"111110000",
46760=>"000111111",
46761=>"110000000",
46762=>"000000111",
46763=>"111101110",
46764=>"110100000",
46765=>"000000000",
46766=>"100000011",
46767=>"010010010",
46768=>"011010100",
46769=>"010010110",
46770=>"000000000",
46771=>"101101110",
46772=>"111011011",
46773=>"000000111",
46774=>"001000000",
46775=>"000010101",
46776=>"001011001",
46777=>"000110110",
46778=>"111110001",
46779=>"000000000",
46780=>"001001000",
46781=>"100111111",
46782=>"111100101",
46783=>"111111010",
46784=>"000000000",
46785=>"111111111",
46786=>"010111010",
46787=>"011001000",
46788=>"000000000",
46789=>"111110110",
46790=>"101100010",
46791=>"000000110",
46792=>"000000110",
46793=>"000000000",
46794=>"010000000",
46795=>"010111000",
46796=>"001001000",
46797=>"001011011",
46798=>"111011001",
46799=>"111110110",
46800=>"111111111",
46801=>"111000000",
46802=>"010110111",
46803=>"000100110",
46804=>"000000101",
46805=>"100110111",
46806=>"100000000",
46807=>"000111000",
46808=>"001000000",
46809=>"011111110",
46810=>"000111111",
46811=>"000000110",
46812=>"111011000",
46813=>"010000111",
46814=>"000000000",
46815=>"011100001",
46816=>"000000000",
46817=>"000000011",
46818=>"111100000",
46819=>"000000000",
46820=>"000000000",
46821=>"001000000",
46822=>"011101101",
46823=>"011010111",
46824=>"000000110",
46825=>"100111011",
46826=>"000000000",
46827=>"000000000",
46828=>"111110010",
46829=>"011000000",
46830=>"000001010",
46831=>"110000000",
46832=>"111100000",
46833=>"111011011",
46834=>"010011110",
46835=>"111100000",
46836=>"111010000",
46837=>"000111110",
46838=>"000000000",
46839=>"111111001",
46840=>"010111000",
46841=>"110111111",
46842=>"010110000",
46843=>"010001001",
46844=>"111110000",
46845=>"100010000",
46846=>"001011011",
46847=>"011111011",
46848=>"110111100",
46849=>"010101101",
46850=>"000000101",
46851=>"000010010",
46852=>"000000001",
46853=>"111110000",
46854=>"000010010",
46855=>"111111100",
46856=>"000000001",
46857=>"000000000",
46858=>"000001000",
46859=>"000000000",
46860=>"010010000",
46861=>"010111111",
46862=>"110001001",
46863=>"111111000",
46864=>"001011100",
46865=>"100111111",
46866=>"010010010",
46867=>"000000000",
46868=>"000000111",
46869=>"110101100",
46870=>"010110110",
46871=>"101111011",
46872=>"011111000",
46873=>"011011001",
46874=>"111111111",
46875=>"000001000",
46876=>"000000000",
46877=>"011000000",
46878=>"111010000",
46879=>"111000000",
46880=>"000010101",
46881=>"010010101",
46882=>"111000011",
46883=>"001100010",
46884=>"111110000",
46885=>"010110010",
46886=>"000011010",
46887=>"000001000",
46888=>"111111101",
46889=>"001110101",
46890=>"100000110",
46891=>"010111101",
46892=>"011011011",
46893=>"111110010",
46894=>"111111001",
46895=>"011001111",
46896=>"000000111",
46897=>"110001001",
46898=>"001010000",
46899=>"111001101",
46900=>"000110111",
46901=>"000000111",
46902=>"110110001",
46903=>"101000000",
46904=>"000001111",
46905=>"011100000",
46906=>"000100100",
46907=>"000001111",
46908=>"100110101",
46909=>"000111011",
46910=>"000001110",
46911=>"000000110",
46912=>"011000101",
46913=>"111111101",
46914=>"111111011",
46915=>"111101111",
46916=>"000000111",
46917=>"101000010",
46918=>"000000000",
46919=>"111101000",
46920=>"111001100",
46921=>"111111000",
46922=>"111000001",
46923=>"101000000",
46924=>"101100000",
46925=>"011111000",
46926=>"000100000",
46927=>"111110111",
46928=>"000010101",
46929=>"010000000",
46930=>"011010000",
46931=>"001000100",
46932=>"010000000",
46933=>"011000111",
46934=>"011001001",
46935=>"111111011",
46936=>"110111101",
46937=>"111001000",
46938=>"010000011",
46939=>"110111000",
46940=>"000000011",
46941=>"000001001",
46942=>"001000100",
46943=>"101101101",
46944=>"000111111",
46945=>"111100110",
46946=>"111010000",
46947=>"000000100",
46948=>"100100000",
46949=>"111100000",
46950=>"110110000",
46951=>"101101111",
46952=>"000100110",
46953=>"111111101",
46954=>"100011011",
46955=>"001010000",
46956=>"011111111",
46957=>"000101000",
46958=>"000000111",
46959=>"010111111",
46960=>"010111011",
46961=>"111111111",
46962=>"011101100",
46963=>"101111010",
46964=>"000111111",
46965=>"000000101",
46966=>"001111111",
46967=>"011011001",
46968=>"111111100",
46969=>"010100000",
46970=>"111001000",
46971=>"000101101",
46972=>"011110101",
46973=>"000100000",
46974=>"000001111",
46975=>"010000110",
46976=>"101111010",
46977=>"010111000",
46978=>"110000000",
46979=>"111001001",
46980=>"111111111",
46981=>"101001000",
46982=>"011111111",
46983=>"111110110",
46984=>"001111011",
46985=>"101101101",
46986=>"101111111",
46987=>"100000000",
46988=>"000101000",
46989=>"110001111",
46990=>"010001111",
46991=>"000001010",
46992=>"110110011",
46993=>"001101111",
46994=>"000101111",
46995=>"011100100",
46996=>"010000000",
46997=>"111010000",
46998=>"101000100",
46999=>"110000111",
47000=>"000101110",
47001=>"000111111",
47002=>"001101111",
47003=>"000001101",
47004=>"000011011",
47005=>"011000100",
47006=>"000100111",
47007=>"000000001",
47008=>"000100000",
47009=>"110000000",
47010=>"111100000",
47011=>"010100111",
47012=>"010000100",
47013=>"010011011",
47014=>"101001000",
47015=>"101000011",
47016=>"111111010",
47017=>"000110111",
47018=>"100110111",
47019=>"110111110",
47020=>"101000011",
47021=>"111111110",
47022=>"100100100",
47023=>"111010000",
47024=>"100000000",
47025=>"110001001",
47026=>"000000100",
47027=>"111000100",
47028=>"110110110",
47029=>"101100100",
47030=>"110100000",
47031=>"001010000",
47032=>"001010111",
47033=>"110010001",
47034=>"010000000",
47035=>"000011111",
47036=>"101100000",
47037=>"111111110",
47038=>"000000001",
47039=>"101101111",
47040=>"000110111",
47041=>"000000000",
47042=>"000111111",
47043=>"110110111",
47044=>"011000000",
47045=>"101001000",
47046=>"111010000",
47047=>"000100010",
47048=>"111010101",
47049=>"100001110",
47050=>"100101100",
47051=>"001000100",
47052=>"000000000",
47053=>"000001111",
47054=>"101101001",
47055=>"000001011",
47056=>"100111000",
47057=>"000100110",
47058=>"011000000",
47059=>"001101011",
47060=>"110011101",
47061=>"111100100",
47062=>"010010000",
47063=>"001111101",
47064=>"101101111",
47065=>"000000111",
47066=>"111100000",
47067=>"000000000",
47068=>"111011110",
47069=>"000011111",
47070=>"111111010",
47071=>"011111000",
47072=>"100111001",
47073=>"100010100",
47074=>"110000000",
47075=>"001111111",
47076=>"000000000",
47077=>"011101111",
47078=>"000000000",
47079=>"010100000",
47080=>"101100111",
47081=>"100111111",
47082=>"101100001",
47083=>"000000111",
47084=>"101100000",
47085=>"010111101",
47086=>"000000000",
47087=>"000000000",
47088=>"000000111",
47089=>"100000100",
47090=>"000010000",
47091=>"011001000",
47092=>"110111001",
47093=>"010111111",
47094=>"000000000",
47095=>"110000000",
47096=>"000000101",
47097=>"000111111",
47098=>"010011000",
47099=>"110010000",
47100=>"101000001",
47101=>"000000100",
47102=>"110111000",
47103=>"000000000",
47104=>"110111001",
47105=>"100101010",
47106=>"001001111",
47107=>"101000000",
47108=>"100000100",
47109=>"010001100",
47110=>"100000001",
47111=>"101011011",
47112=>"100101111",
47113=>"000011011",
47114=>"010010100",
47115=>"000010111",
47116=>"111000000",
47117=>"010111111",
47118=>"100100100",
47119=>"000100110",
47120=>"000110111",
47121=>"111111000",
47122=>"111010000",
47123=>"001001001",
47124=>"001111101",
47125=>"111101101",
47126=>"110010000",
47127=>"001010010",
47128=>"100000001",
47129=>"101111111",
47130=>"000111111",
47131=>"000000000",
47132=>"000000111",
47133=>"111111011",
47134=>"011010000",
47135=>"011010111",
47136=>"011001101",
47137=>"111011000",
47138=>"000010110",
47139=>"011010000",
47140=>"000110100",
47141=>"100000100",
47142=>"111001000",
47143=>"100111101",
47144=>"111101111",
47145=>"001010010",
47146=>"000000110",
47147=>"010000001",
47148=>"011111101",
47149=>"010010111",
47150=>"000001000",
47151=>"001000111",
47152=>"111101000",
47153=>"101100110",
47154=>"100010000",
47155=>"010000101",
47156=>"111111100",
47157=>"111101100",
47158=>"011011001",
47159=>"000111110",
47160=>"011000001",
47161=>"101100101",
47162=>"000010000",
47163=>"100010010",
47164=>"000000100",
47165=>"111111110",
47166=>"000110100",
47167=>"100000011",
47168=>"101000000",
47169=>"010100110",
47170=>"000000010",
47171=>"000000100",
47172=>"111111000",
47173=>"000000110",
47174=>"000000000",
47175=>"101000000",
47176=>"001111111",
47177=>"100000000",
47178=>"101100111",
47179=>"000000001",
47180=>"000010010",
47181=>"111111111",
47182=>"111111001",
47183=>"010111111",
47184=>"111011000",
47185=>"101011111",
47186=>"000001010",
47187=>"111001011",
47188=>"110000101",
47189=>"100010110",
47190=>"110010011",
47191=>"010000001",
47192=>"000101001",
47193=>"101000000",
47194=>"011001100",
47195=>"000000001",
47196=>"111010000",
47197=>"010001100",
47198=>"111111010",
47199=>"001000001",
47200=>"000010000",
47201=>"001100000",
47202=>"000111000",
47203=>"000100001",
47204=>"110010111",
47205=>"001011001",
47206=>"111000110",
47207=>"011101111",
47208=>"000000011",
47209=>"100000000",
47210=>"000010011",
47211=>"111000000",
47212=>"110011000",
47213=>"010010111",
47214=>"000010000",
47215=>"000001111",
47216=>"011011011",
47217=>"100010111",
47218=>"100100100",
47219=>"010010010",
47220=>"000010111",
47221=>"000000101",
47222=>"000100011",
47223=>"111111000",
47224=>"011000001",
47225=>"000000000",
47226=>"100010010",
47227=>"101100101",
47228=>"110101110",
47229=>"011110001",
47230=>"010000001",
47231=>"000000101",
47232=>"101010000",
47233=>"111000000",
47234=>"100000101",
47235=>"111111000",
47236=>"111000000",
47237=>"000001000",
47238=>"000000001",
47239=>"000001011",
47240=>"011110110",
47241=>"110100101",
47242=>"000011011",
47243=>"101000000",
47244=>"000000101",
47245=>"101001101",
47246=>"000000101",
47247=>"000000100",
47248=>"100101001",
47249=>"100000000",
47250=>"000000101",
47251=>"100000001",
47252=>"000000001",
47253=>"000000000",
47254=>"001010000",
47255=>"111111000",
47256=>"110111111",
47257=>"101000001",
47258=>"001011111",
47259=>"000000101",
47260=>"011111110",
47261=>"000010000",
47262=>"000101111",
47263=>"011010000",
47264=>"000011001",
47265=>"101011101",
47266=>"101000100",
47267=>"111110010",
47268=>"011000100",
47269=>"000110110",
47270=>"111111000",
47271=>"000000111",
47272=>"110010111",
47273=>"001101000",
47274=>"101101101",
47275=>"010111000",
47276=>"110001000",
47277=>"111110010",
47278=>"111111100",
47279=>"111010110",
47280=>"111001010",
47281=>"010001101",
47282=>"111101111",
47283=>"100110010",
47284=>"111111011",
47285=>"110001000",
47286=>"111011011",
47287=>"000010111",
47288=>"000000001",
47289=>"100100100",
47290=>"011000001",
47291=>"111010010",
47292=>"100011110",
47293=>"001111010",
47294=>"001001101",
47295=>"010000010",
47296=>"100000000",
47297=>"111000000",
47298=>"000001000",
47299=>"111110110",
47300=>"011000000",
47301=>"101000000",
47302=>"100110111",
47303=>"110101111",
47304=>"100011111",
47305=>"011000001",
47306=>"101111111",
47307=>"111011111",
47308=>"000100100",
47309=>"011101000",
47310=>"010000000",
47311=>"010000000",
47312=>"001100101",
47313=>"110110110",
47314=>"101011111",
47315=>"000010010",
47316=>"100100101",
47317=>"011110011",
47318=>"000001101",
47319=>"101101111",
47320=>"111000010",
47321=>"010000101",
47322=>"101110101",
47323=>"110000000",
47324=>"011011101",
47325=>"010010100",
47326=>"111111111",
47327=>"010000000",
47328=>"000001000",
47329=>"000000000",
47330=>"111000110",
47331=>"000101111",
47332=>"110100001",
47333=>"000111001",
47334=>"000111111",
47335=>"100101001",
47336=>"000111011",
47337=>"111110000",
47338=>"100011001",
47339=>"111011010",
47340=>"111000001",
47341=>"000000000",
47342=>"010011110",
47343=>"010110001",
47344=>"101101101",
47345=>"011000000",
47346=>"110100011",
47347=>"100110111",
47348=>"001111111",
47349=>"000000000",
47350=>"000101000",
47351=>"010000000",
47352=>"000000000",
47353=>"001111010",
47354=>"111111011",
47355=>"001000000",
47356=>"111111010",
47357=>"111101110",
47358=>"011010001",
47359=>"100100001",
47360=>"100100100",
47361=>"011001100",
47362=>"110111001",
47363=>"000000000",
47364=>"110111100",
47365=>"000000000",
47366=>"100000000",
47367=>"100101111",
47368=>"111110000",
47369=>"111111010",
47370=>"110111011",
47371=>"000000000",
47372=>"100000000",
47373=>"110100111",
47374=>"001011110",
47375=>"011101111",
47376=>"000110000",
47377=>"011111001",
47378=>"010111010",
47379=>"001100000",
47380=>"110111111",
47381=>"000110000",
47382=>"010101100",
47383=>"110000111",
47384=>"111000000",
47385=>"111000101",
47386=>"011001000",
47387=>"000111011",
47388=>"011001111",
47389=>"100111111",
47390=>"100111000",
47391=>"111001000",
47392=>"010111111",
47393=>"000000000",
47394=>"111100100",
47395=>"010000000",
47396=>"110111110",
47397=>"000011011",
47398=>"010011010",
47399=>"000111111",
47400=>"111111111",
47401=>"111011111",
47402=>"000000000",
47403=>"000000000",
47404=>"000001001",
47405=>"001100010",
47406=>"100000101",
47407=>"011001111",
47408=>"000000111",
47409=>"110110111",
47410=>"111110111",
47411=>"000000011",
47412=>"000000000",
47413=>"000000000",
47414=>"011111011",
47415=>"100000010",
47416=>"100100011",
47417=>"101101000",
47418=>"100100101",
47419=>"000111110",
47420=>"010000111",
47421=>"111111011",
47422=>"010101101",
47423=>"000110110",
47424=>"000011000",
47425=>"000011101",
47426=>"111110111",
47427=>"010010010",
47428=>"010010010",
47429=>"101001000",
47430=>"001111101",
47431=>"011000011",
47432=>"000000010",
47433=>"000111111",
47434=>"111101001",
47435=>"000000000",
47436=>"010110010",
47437=>"001011011",
47438=>"111010111",
47439=>"111111111",
47440=>"000010010",
47441=>"111111111",
47442=>"000000000",
47443=>"001001011",
47444=>"000011000",
47445=>"000000000",
47446=>"011001011",
47447=>"111011111",
47448=>"111101000",
47449=>"111111111",
47450=>"001011000",
47451=>"000000010",
47452=>"100000000",
47453=>"101001001",
47454=>"110111011",
47455=>"110011111",
47456=>"010111111",
47457=>"110000010",
47458=>"000100100",
47459=>"010111110",
47460=>"100000100",
47461=>"110111111",
47462=>"000111110",
47463=>"011111100",
47464=>"000000010",
47465=>"000111111",
47466=>"111111111",
47467=>"001000110",
47468=>"111111111",
47469=>"000011111",
47470=>"000000101",
47471=>"010110100",
47472=>"011011111",
47473=>"000000101",
47474=>"011111010",
47475=>"100000000",
47476=>"111101111",
47477=>"100100100",
47478=>"111001111",
47479=>"010010010",
47480=>"101001000",
47481=>"000000000",
47482=>"000000000",
47483=>"101110010",
47484=>"001000101",
47485=>"110101110",
47486=>"000101111",
47487=>"111011010",
47488=>"100111111",
47489=>"111000000",
47490=>"000100000",
47491=>"011011111",
47492=>"000000000",
47493=>"111111111",
47494=>"100110110",
47495=>"100000100",
47496=>"100111111",
47497=>"100110110",
47498=>"111111111",
47499=>"000001111",
47500=>"110000000",
47501=>"000000100",
47502=>"101000000",
47503=>"000000000",
47504=>"001001001",
47505=>"001010000",
47506=>"010111011",
47507=>"011000000",
47508=>"111000010",
47509=>"011001001",
47510=>"000111011",
47511=>"110100110",
47512=>"110111101",
47513=>"101000000",
47514=>"011010011",
47515=>"000000000",
47516=>"000000000",
47517=>"000010000",
47518=>"000001000",
47519=>"001000000",
47520=>"000000000",
47521=>"011110000",
47522=>"111101111",
47523=>"111111000",
47524=>"100100101",
47525=>"011001010",
47526=>"111001100",
47527=>"000010000",
47528=>"101111110",
47529=>"100010111",
47530=>"100000100",
47531=>"110101001",
47532=>"111101111",
47533=>"011111011",
47534=>"100001011",
47535=>"100000100",
47536=>"000000100",
47537=>"000001011",
47538=>"000000001",
47539=>"111000000",
47540=>"111110011",
47541=>"111000100",
47542=>"111111111",
47543=>"000100111",
47544=>"000000001",
47545=>"011011010",
47546=>"000111111",
47547=>"000100110",
47548=>"101111011",
47549=>"111111111",
47550=>"110000010",
47551=>"000100001",
47552=>"101000000",
47553=>"000000000",
47554=>"000000111",
47555=>"100110110",
47556=>"000000010",
47557=>"001000100",
47558=>"000010101",
47559=>"000000000",
47560=>"100100000",
47561=>"111000000",
47562=>"111111011",
47563=>"011011010",
47564=>"001111011",
47565=>"100100000",
47566=>"000000000",
47567=>"111110000",
47568=>"011011010",
47569=>"110110110",
47570=>"011000000",
47571=>"101100100",
47572=>"000000000",
47573=>"000101100",
47574=>"000010011",
47575=>"001101111",
47576=>"000000100",
47577=>"001010010",
47578=>"111110101",
47579=>"100000100",
47580=>"100000000",
47581=>"000001101",
47582=>"011000000",
47583=>"001000000",
47584=>"000110000",
47585=>"100000000",
47586=>"101000000",
47587=>"000010001",
47588=>"000010000",
47589=>"000000001",
47590=>"111000000",
47591=>"000000100",
47592=>"000101111",
47593=>"000000101",
47594=>"011111110",
47595=>"001000101",
47596=>"111101101",
47597=>"000000000",
47598=>"101001000",
47599=>"111000000",
47600=>"111111111",
47601=>"110001101",
47602=>"100100111",
47603=>"111111110",
47604=>"011010111",
47605=>"000111010",
47606=>"000000010",
47607=>"000100111",
47608=>"000000101",
47609=>"100001011",
47610=>"110000000",
47611=>"000001101",
47612=>"000010000",
47613=>"000000100",
47614=>"100111010",
47615=>"000100100",
47616=>"011011111",
47617=>"000000000",
47618=>"010010010",
47619=>"111110000",
47620=>"101001000",
47621=>"000010001",
47622=>"000101111",
47623=>"110111111",
47624=>"111000101",
47625=>"001101111",
47626=>"001000000",
47627=>"000000000",
47628=>"110010011",
47629=>"111111111",
47630=>"100000001",
47631=>"010101011",
47632=>"000111110",
47633=>"101101000",
47634=>"000100000",
47635=>"000000000",
47636=>"000000100",
47637=>"110111100",
47638=>"000011000",
47639=>"101111111",
47640=>"000000000",
47641=>"000000000",
47642=>"000000000",
47643=>"101001111",
47644=>"101101101",
47645=>"101111001",
47646=>"100010011",
47647=>"111111101",
47648=>"101000000",
47649=>"000100000",
47650=>"100110010",
47651=>"000000101",
47652=>"001000101",
47653=>"100111001",
47654=>"000010000",
47655=>"001001111",
47656=>"101111111",
47657=>"101010101",
47658=>"000000001",
47659=>"000000000",
47660=>"000000111",
47661=>"100111011",
47662=>"111100100",
47663=>"100100011",
47664=>"111001011",
47665=>"111000111",
47666=>"000101100",
47667=>"100010010",
47668=>"000101110",
47669=>"110010010",
47670=>"000001000",
47671=>"111101101",
47672=>"101110110",
47673=>"111111111",
47674=>"100101101",
47675=>"000000001",
47676=>"101111100",
47677=>"000111111",
47678=>"000001011",
47679=>"111111111",
47680=>"111010000",
47681=>"000000110",
47682=>"111101101",
47683=>"001001101",
47684=>"000010111",
47685=>"110000000",
47686=>"000011010",
47687=>"000111010",
47688=>"111111111",
47689=>"000000101",
47690=>"100101101",
47691=>"110010111",
47692=>"111111111",
47693=>"000010111",
47694=>"110100111",
47695=>"001000010",
47696=>"000001101",
47697=>"001111000",
47698=>"101001010",
47699=>"001011111",
47700=>"000010111",
47701=>"000000010",
47702=>"000100110",
47703=>"001001010",
47704=>"100110000",
47705=>"001010110",
47706=>"000100111",
47707=>"011011110",
47708=>"001000100",
47709=>"001000001",
47710=>"111011010",
47711=>"100100101",
47712=>"000000000",
47713=>"000111111",
47714=>"000010000",
47715=>"101111111",
47716=>"110001111",
47717=>"111001100",
47718=>"110000001",
47719=>"111001000",
47720=>"011111111",
47721=>"101000000",
47722=>"011100000",
47723=>"111111011",
47724=>"000111001",
47725=>"000000000",
47726=>"000011001",
47727=>"111101010",
47728=>"001101111",
47729=>"101000100",
47730=>"000110010",
47731=>"100110110",
47732=>"111111111",
47733=>"001001101",
47734=>"111111000",
47735=>"000001110",
47736=>"000000110",
47737=>"000000000",
47738=>"000110111",
47739=>"000101111",
47740=>"100000000",
47741=>"100100101",
47742=>"000110110",
47743=>"010111101",
47744=>"000000111",
47745=>"010010010",
47746=>"111000000",
47747=>"110101100",
47748=>"010000010",
47749=>"110111000",
47750=>"001010110",
47751=>"000100001",
47752=>"000111111",
47753=>"000001011",
47754=>"111111111",
47755=>"011000110",
47756=>"011010000",
47757=>"000011011",
47758=>"010110010",
47759=>"000110101",
47760=>"001000100",
47761=>"010110101",
47762=>"101111101",
47763=>"111011010",
47764=>"111111110",
47765=>"000000000",
47766=>"010010010",
47767=>"111000101",
47768=>"000000000",
47769=>"011000001",
47770=>"000110000",
47771=>"000000000",
47772=>"001001000",
47773=>"000001101",
47774=>"101101011",
47775=>"000000000",
47776=>"100001111",
47777=>"111111011",
47778=>"000111111",
47779=>"000010010",
47780=>"000000110",
47781=>"000001001",
47782=>"010000100",
47783=>"000111111",
47784=>"000000010",
47785=>"110010000",
47786=>"000000000",
47787=>"000000000",
47788=>"000001001",
47789=>"101101111",
47790=>"110100001",
47791=>"011111110",
47792=>"111111101",
47793=>"001101101",
47794=>"100000111",
47795=>"000001000",
47796=>"111000100",
47797=>"111111001",
47798=>"000011001",
47799=>"101111111",
47800=>"100101101",
47801=>"110100000",
47802=>"111111100",
47803=>"101010001",
47804=>"111000000",
47805=>"011000000",
47806=>"000000010",
47807=>"000100100",
47808=>"111111111",
47809=>"010000000",
47810=>"101111111",
47811=>"001001100",
47812=>"000100100",
47813=>"001000110",
47814=>"111000011",
47815=>"101111010",
47816=>"000101111",
47817=>"111111110",
47818=>"000000000",
47819=>"011010000",
47820=>"011001100",
47821=>"001100000",
47822=>"000000000",
47823=>"111101100",
47824=>"111111111",
47825=>"100000011",
47826=>"111010000",
47827=>"101000000",
47828=>"010000000",
47829=>"000100000",
47830=>"100100111",
47831=>"101001111",
47832=>"000000111",
47833=>"010001011",
47834=>"110100010",
47835=>"101000000",
47836=>"001010010",
47837=>"000001100",
47838=>"110010011",
47839=>"111111110",
47840=>"000010011",
47841=>"100011011",
47842=>"010011111",
47843=>"000100100",
47844=>"011010001",
47845=>"010110111",
47846=>"001011110",
47847=>"101011100",
47848=>"000001010",
47849=>"000000010",
47850=>"000000100",
47851=>"000011000",
47852=>"111000000",
47853=>"000001100",
47854=>"000000001",
47855=>"101000101",
47856=>"111110000",
47857=>"100000110",
47858=>"001100110",
47859=>"101000011",
47860=>"110101000",
47861=>"000100101",
47862=>"000000000",
47863=>"100000011",
47864=>"010011010",
47865=>"100101100",
47866=>"100110100",
47867=>"111000000",
47868=>"101101010",
47869=>"000100101",
47870=>"110100001",
47871=>"000101000",
47872=>"011011100",
47873=>"000000000",
47874=>"101000000",
47875=>"010010011",
47876=>"000100000",
47877=>"010011000",
47878=>"000001000",
47879=>"011010010",
47880=>"011110100",
47881=>"010011110",
47882=>"000000111",
47883=>"000000010",
47884=>"011000001",
47885=>"000010011",
47886=>"100100001",
47887=>"110001000",
47888=>"000011011",
47889=>"100000111",
47890=>"101100101",
47891=>"100000010",
47892=>"011010011",
47893=>"000100111",
47894=>"000000000",
47895=>"111101111",
47896=>"100000001",
47897=>"011000101",
47898=>"011111111",
47899=>"000011011",
47900=>"111100101",
47901=>"101000000",
47902=>"010010000",
47903=>"111000101",
47904=>"111111000",
47905=>"011100100",
47906=>"111111101",
47907=>"000000111",
47908=>"001111001",
47909=>"011110000",
47910=>"100110110",
47911=>"101001000",
47912=>"011001010",
47913=>"111111000",
47914=>"111011011",
47915=>"111011000",
47916=>"001011111",
47917=>"101101110",
47918=>"011011100",
47919=>"000000000",
47920=>"010011000",
47921=>"101101101",
47922=>"111101110",
47923=>"101000000",
47924=>"000111011",
47925=>"101001110",
47926=>"000000000",
47927=>"010110000",
47928=>"010101000",
47929=>"000000111",
47930=>"101100111",
47931=>"000100000",
47932=>"000100000",
47933=>"111000000",
47934=>"000011011",
47935=>"010111111",
47936=>"010001010",
47937=>"111011000",
47938=>"111111000",
47939=>"000011010",
47940=>"111000010",
47941=>"010100010",
47942=>"101010011",
47943=>"101000101",
47944=>"000001110",
47945=>"010011100",
47946=>"000000011",
47947=>"100010010",
47948=>"111111111",
47949=>"000111111",
47950=>"001111110",
47951=>"101111110",
47952=>"100010111",
47953=>"111101111",
47954=>"000110100",
47955=>"001001010",
47956=>"100111111",
47957=>"001000110",
47958=>"001100100",
47959=>"000111111",
47960=>"001000111",
47961=>"010110001",
47962=>"101101101",
47963=>"011011010",
47964=>"001000000",
47965=>"100001000",
47966=>"000000111",
47967=>"000010010",
47968=>"000010111",
47969=>"111000011",
47970=>"000010111",
47971=>"011100100",
47972=>"000111100",
47973=>"111001000",
47974=>"111110000",
47975=>"111100100",
47976=>"111010110",
47977=>"111101101",
47978=>"010011111",
47979=>"111010101",
47980=>"110000001",
47981=>"000111111",
47982=>"000011011",
47983=>"011111100",
47984=>"000111100",
47985=>"011011000",
47986=>"000000000",
47987=>"111100100",
47988=>"010110111",
47989=>"001000100",
47990=>"101010010",
47991=>"010011101",
47992=>"000000000",
47993=>"111101001",
47994=>"111101101",
47995=>"011001000",
47996=>"100000000",
47997=>"010110000",
47998=>"000101011",
47999=>"000010010",
48000=>"000000000",
48001=>"100100110",
48002=>"011010000",
48003=>"111110111",
48004=>"011101000",
48005=>"101000000",
48006=>"110111000",
48007=>"000110110",
48008=>"010111001",
48009=>"100100111",
48010=>"100011011",
48011=>"000000100",
48012=>"101001011",
48013=>"001111010",
48014=>"010001011",
48015=>"000000001",
48016=>"111101101",
48017=>"111111000",
48018=>"100100110",
48019=>"000010100",
48020=>"000010010",
48021=>"000000010",
48022=>"110111001",
48023=>"001101000",
48024=>"000010010",
48025=>"101001111",
48026=>"100100011",
48027=>"100100111",
48028=>"000010000",
48029=>"001010000",
48030=>"010000111",
48031=>"100101100",
48032=>"100100110",
48033=>"001000000",
48034=>"010000011",
48035=>"100000001",
48036=>"111100101",
48037=>"100011011",
48038=>"010101000",
48039=>"000111111",
48040=>"100000000",
48041=>"001101011",
48042=>"010101111",
48043=>"000000000",
48044=>"011110100",
48045=>"010011110",
48046=>"011110111",
48047=>"111110010",
48048=>"010111111",
48049=>"100000001",
48050=>"101111000",
48051=>"101101000",
48052=>"001111100",
48053=>"101011100",
48054=>"011010000",
48055=>"111011000",
48056=>"000001000",
48057=>"000110101",
48058=>"011011100",
48059=>"000101100",
48060=>"011000001",
48061=>"111110111",
48062=>"001111000",
48063=>"001101111",
48064=>"100010110",
48065=>"010011111",
48066=>"111001011",
48067=>"000011101",
48068=>"011101101",
48069=>"000100001",
48070=>"010000000",
48071=>"111011110",
48072=>"111011111",
48073=>"000110000",
48074=>"011000000",
48075=>"011011010",
48076=>"100010010",
48077=>"000000000",
48078=>"100011011",
48079=>"011001000",
48080=>"100100111",
48081=>"011111000",
48082=>"010000100",
48083=>"111101110",
48084=>"000001011",
48085=>"000110110",
48086=>"100001101",
48087=>"010001000",
48088=>"110101111",
48089=>"000000111",
48090=>"011011111",
48091=>"101000001",
48092=>"000100000",
48093=>"111011111",
48094=>"000000101",
48095=>"011000000",
48096=>"000011111",
48097=>"111001101",
48098=>"111101100",
48099=>"000011110",
48100=>"000000000",
48101=>"110100100",
48102=>"111011010",
48103=>"000011111",
48104=>"000011010",
48105=>"000010000",
48106=>"100000111",
48107=>"011111111",
48108=>"100000110",
48109=>"010110110",
48110=>"000000000",
48111=>"000000000",
48112=>"111000111",
48113=>"000101111",
48114=>"011011000",
48115=>"001101101",
48116=>"010110000",
48117=>"101000111",
48118=>"000000001",
48119=>"011111000",
48120=>"100000010",
48121=>"101100111",
48122=>"010000111",
48123=>"000000111",
48124=>"100011011",
48125=>"111100101",
48126=>"011110110",
48127=>"101011000",
48128=>"000100000",
48129=>"000001010",
48130=>"100000000",
48131=>"000001000",
48132=>"111111011",
48133=>"000000001",
48134=>"000000111",
48135=>"000000001",
48136=>"100010110",
48137=>"111101111",
48138=>"111111111",
48139=>"110010000",
48140=>"110010111",
48141=>"111101111",
48142=>"000101000",
48143=>"110111111",
48144=>"111110011",
48145=>"000000100",
48146=>"011010010",
48147=>"000000110",
48148=>"100001000",
48149=>"111010000",
48150=>"111111111",
48151=>"110011111",
48152=>"001001001",
48153=>"101111001",
48154=>"000010001",
48155=>"100100101",
48156=>"000001000",
48157=>"000000001",
48158=>"010011110",
48159=>"000000001",
48160=>"000001000",
48161=>"000000001",
48162=>"001000011",
48163=>"111001001",
48164=>"100000101",
48165=>"100110000",
48166=>"111011010",
48167=>"111111111",
48168=>"111000111",
48169=>"001000100",
48170=>"000000110",
48171=>"110110011",
48172=>"011111111",
48173=>"011000000",
48174=>"100100100",
48175=>"100001001",
48176=>"101100000",
48177=>"000000000",
48178=>"000000011",
48179=>"000000011",
48180=>"111111000",
48181=>"000000000",
48182=>"110100100",
48183=>"000000000",
48184=>"000000000",
48185=>"001001001",
48186=>"010010010",
48187=>"110111111",
48188=>"000000000",
48189=>"111111111",
48190=>"000101111",
48191=>"110110111",
48192=>"100110111",
48193=>"111110010",
48194=>"000011111",
48195=>"110111011",
48196=>"100101111",
48197=>"011000100",
48198=>"100110111",
48199=>"111111111",
48200=>"000000000",
48201=>"111111111",
48202=>"111000101",
48203=>"010111111",
48204=>"001000000",
48205=>"011011011",
48206=>"111111111",
48207=>"111111111",
48208=>"100000101",
48209=>"111111011",
48210=>"111101111",
48211=>"000000000",
48212=>"000111111",
48213=>"000000010",
48214=>"010100110",
48215=>"101001111",
48216=>"000001001",
48217=>"111111111",
48218=>"000100100",
48219=>"111110111",
48220=>"000000001",
48221=>"000000000",
48222=>"010000010",
48223=>"111111110",
48224=>"111001111",
48225=>"110111111",
48226=>"000000001",
48227=>"001111011",
48228=>"000001101",
48229=>"011111000",
48230=>"000110111",
48231=>"010000000",
48232=>"001111110",
48233=>"101111010",
48234=>"000000110",
48235=>"000000100",
48236=>"101000111",
48237=>"101101001",
48238=>"110111110",
48239=>"100101001",
48240=>"110110110",
48241=>"000000100",
48242=>"001001100",
48243=>"110110111",
48244=>"011011111",
48245=>"000000111",
48246=>"000000000",
48247=>"010011111",
48248=>"111111111",
48249=>"011111111",
48250=>"000000110",
48251=>"100000100",
48252=>"010110110",
48253=>"000000000",
48254=>"111011111",
48255=>"101111101",
48256=>"000101011",
48257=>"111111111",
48258=>"000000000",
48259=>"001100111",
48260=>"000000000",
48261=>"000001111",
48262=>"011011010",
48263=>"010010000",
48264=>"101001011",
48265=>"101111111",
48266=>"111111010",
48267=>"000000110",
48268=>"000111011",
48269=>"111110110",
48270=>"000110110",
48271=>"000000101",
48272=>"001001111",
48273=>"000000000",
48274=>"000000000",
48275=>"011010111",
48276=>"000110111",
48277=>"000000110",
48278=>"111110110",
48279=>"000000011",
48280=>"111100010",
48281=>"111111111",
48282=>"011110110",
48283=>"110110110",
48284=>"000111111",
48285=>"111110000",
48286=>"000000000",
48287=>"000101101",
48288=>"110110011",
48289=>"111111111",
48290=>"101000101",
48291=>"011111011",
48292=>"111000000",
48293=>"110111111",
48294=>"111111001",
48295=>"001001001",
48296=>"000001011",
48297=>"000000000",
48298=>"001000000",
48299=>"101101111",
48300=>"111111111",
48301=>"000000000",
48302=>"101101101",
48303=>"111111110",
48304=>"111111111",
48305=>"000000100",
48306=>"000110000",
48307=>"011011100",
48308=>"111001111",
48309=>"001111010",
48310=>"000011111",
48311=>"000010000",
48312=>"001001000",
48313=>"000111110",
48314=>"001110100",
48315=>"100111110",
48316=>"100000001",
48317=>"111011100",
48318=>"111110110",
48319=>"001001110",
48320=>"110110010",
48321=>"111110000",
48322=>"110101000",
48323=>"010010110",
48324=>"000000000",
48325=>"100000000",
48326=>"100000111",
48327=>"010111110",
48328=>"001000000",
48329=>"111111110",
48330=>"010011111",
48331=>"110111000",
48332=>"100100011",
48333=>"000010010",
48334=>"000000001",
48335=>"000111001",
48336=>"111111000",
48337=>"110110110",
48338=>"101000000",
48339=>"000000000",
48340=>"011011001",
48341=>"001001000",
48342=>"000000001",
48343=>"111100000",
48344=>"111001001",
48345=>"111100000",
48346=>"001011011",
48347=>"111111110",
48348=>"011111110",
48349=>"001111111",
48350=>"110111111",
48351=>"000000000",
48352=>"111110000",
48353=>"010001111",
48354=>"001000000",
48355=>"111111111",
48356=>"101001001",
48357=>"111000111",
48358=>"100000101",
48359=>"111111111",
48360=>"000000000",
48361=>"000101111",
48362=>"111111111",
48363=>"111111111",
48364=>"111101001",
48365=>"000011000",
48366=>"000000001",
48367=>"000000000",
48368=>"000000001",
48369=>"001001000",
48370=>"101110101",
48371=>"110000000",
48372=>"001111111",
48373=>"110111001",
48374=>"000001111",
48375=>"110000000",
48376=>"010000000",
48377=>"000000000",
48378=>"111111111",
48379=>"000101000",
48380=>"000010000",
48381=>"000100111",
48382=>"100100100",
48383=>"000111111",
48384=>"001001001",
48385=>"000100111",
48386=>"101100101",
48387=>"011010011",
48388=>"110100111",
48389=>"010010010",
48390=>"111100100",
48391=>"000010011",
48392=>"000100101",
48393=>"000000001",
48394=>"101100100",
48395=>"111100000",
48396=>"000011010",
48397=>"000010000",
48398=>"100111011",
48399=>"001100111",
48400=>"110000101",
48401=>"000000111",
48402=>"101000111",
48403=>"111100100",
48404=>"000000101",
48405=>"000000010",
48406=>"111111111",
48407=>"111101100",
48408=>"111100100",
48409=>"110001101",
48410=>"000000010",
48411=>"111101111",
48412=>"000100101",
48413=>"100000000",
48414=>"111111011",
48415=>"101000000",
48416=>"000000000",
48417=>"010011011",
48418=>"101101111",
48419=>"000010010",
48420=>"001011010",
48421=>"010110100",
48422=>"000010010",
48423=>"000000111",
48424=>"101010111",
48425=>"001010000",
48426=>"101000100",
48427=>"110000000",
48428=>"111001001",
48429=>"111100111",
48430=>"011000100",
48431=>"111111110",
48432=>"011011111",
48433=>"011110101",
48434=>"000111111",
48435=>"111000000",
48436=>"111000000",
48437=>"000100000",
48438=>"000010011",
48439=>"010111100",
48440=>"010010000",
48441=>"000001001",
48442=>"011100111",
48443=>"100100000",
48444=>"000111110",
48445=>"110111010",
48446=>"000000000",
48447=>"100110110",
48448=>"000000110",
48449=>"101011001",
48450=>"011111111",
48451=>"011011000",
48452=>"000000010",
48453=>"011000100",
48454=>"000000000",
48455=>"000010000",
48456=>"000001010",
48457=>"000011111",
48458=>"101000000",
48459=>"111100100",
48460=>"111011000",
48461=>"100110011",
48462=>"011011010",
48463=>"101000111",
48464=>"101110000",
48465=>"111010000",
48466=>"111101111",
48467=>"010000000",
48468=>"111101100",
48469=>"010111111",
48470=>"010011001",
48471=>"111000000",
48472=>"111000100",
48473=>"100110100",
48474=>"100010010",
48475=>"000011001",
48476=>"000011011",
48477=>"111001001",
48478=>"100011111",
48479=>"000000010",
48480=>"000011111",
48481=>"000000111",
48482=>"111000000",
48483=>"111101101",
48484=>"000100000",
48485=>"111110010",
48486=>"111100000",
48487=>"001011000",
48488=>"111011111",
48489=>"010111000",
48490=>"000010010",
48491=>"001000000",
48492=>"100100000",
48493=>"011000101",
48494=>"010000000",
48495=>"111000010",
48496=>"000000100",
48497=>"010011000",
48498=>"000010111",
48499=>"111011011",
48500=>"000111111",
48501=>"100100100",
48502=>"010011010",
48503=>"000111010",
48504=>"101111000",
48505=>"011011011",
48506=>"111000000",
48507=>"000101100",
48508=>"100110100",
48509=>"010100000",
48510=>"111100111",
48511=>"100000000",
48512=>"111011010",
48513=>"000000000",
48514=>"000111011",
48515=>"000000011",
48516=>"101001000",
48517=>"111000000",
48518=>"100111000",
48519=>"110101100",
48520=>"000000100",
48521=>"101100000",
48522=>"111100110",
48523=>"111011000",
48524=>"000000101",
48525=>"101101111",
48526=>"110111110",
48527=>"001000000",
48528=>"100100000",
48529=>"100100101",
48530=>"111100111",
48531=>"111011100",
48532=>"100110000",
48533=>"110110000",
48534=>"011111011",
48535=>"000011011",
48536=>"010100100",
48537=>"011100111",
48538=>"000111011",
48539=>"100100110",
48540=>"001111000",
48541=>"110111100",
48542=>"011010000",
48543=>"111000000",
48544=>"000100111",
48545=>"110111010",
48546=>"000011001",
48547=>"011100011",
48548=>"000000000",
48549=>"000011100",
48550=>"101111010",
48551=>"000011011",
48552=>"100111111",
48553=>"000010111",
48554=>"111000000",
48555=>"110100100",
48556=>"111010000",
48557=>"000011011",
48558=>"111110110",
48559=>"111111011",
48560=>"000100100",
48561=>"011001001",
48562=>"111111100",
48563=>"000111100",
48564=>"000011011",
48565=>"111111111",
48566=>"000100110",
48567=>"000011001",
48568=>"101111011",
48569=>"001111000",
48570=>"111010001",
48571=>"111000010",
48572=>"011000001",
48573=>"000111111",
48574=>"000011111",
48575=>"111100011",
48576=>"111000000",
48577=>"001000000",
48578=>"001101111",
48579=>"011011010",
48580=>"110101101",
48581=>"001011101",
48582=>"111110100",
48583=>"111001101",
48584=>"000000100",
48585=>"000011010",
48586=>"010111011",
48587=>"000100111",
48588=>"100100000",
48589=>"000001111",
48590=>"101001000",
48591=>"001001000",
48592=>"000000111",
48593=>"000110110",
48594=>"111000000",
48595=>"000111011",
48596=>"111100110",
48597=>"110100110",
48598=>"100000000",
48599=>"000001111",
48600=>"111000000",
48601=>"000100000",
48602=>"001111100",
48603=>"111000000",
48604=>"110011111",
48605=>"100101111",
48606=>"000100000",
48607=>"111111000",
48608=>"000111111",
48609=>"011000010",
48610=>"111000000",
48611=>"000000110",
48612=>"000100000",
48613=>"111000100",
48614=>"110000101",
48615=>"000001011",
48616=>"010011111",
48617=>"001000001",
48618=>"100100000",
48619=>"111000100",
48620=>"000111111",
48621=>"000000000",
48622=>"000100000",
48623=>"000100100",
48624=>"111000000",
48625=>"000111101",
48626=>"100011000",
48627=>"000011110",
48628=>"010110011",
48629=>"111111111",
48630=>"000000110",
48631=>"000101011",
48632=>"110000000",
48633=>"101001111",
48634=>"010100010",
48635=>"101001001",
48636=>"000111000",
48637=>"011100100",
48638=>"001001001",
48639=>"101100000",
48640=>"110101000",
48641=>"100010101",
48642=>"101000111",
48643=>"000000010",
48644=>"111101101",
48645=>"101100111",
48646=>"000111000",
48647=>"111111010",
48648=>"001000000",
48649=>"111000100",
48650=>"001000101",
48651=>"011000110",
48652=>"111000101",
48653=>"000101101",
48654=>"100100100",
48655=>"111111011",
48656=>"000010101",
48657=>"000000000",
48658=>"011001010",
48659=>"111111000",
48660=>"010011011",
48661=>"000000000",
48662=>"110111100",
48663=>"111011101",
48664=>"110000111",
48665=>"000111000",
48666=>"111101111",
48667=>"000000111",
48668=>"011000010",
48669=>"000000000",
48670=>"000000111",
48671=>"111000000",
48672=>"000111001",
48673=>"111000111",
48674=>"000100101",
48675=>"001100111",
48676=>"110011001",
48677=>"000001111",
48678=>"000010000",
48679=>"111111110",
48680=>"001001000",
48681=>"011110101",
48682=>"111111011",
48683=>"010011000",
48684=>"111010011",
48685=>"111000000",
48686=>"101110100",
48687=>"100000011",
48688=>"110000111",
48689=>"111111101",
48690=>"101000000",
48691=>"000000001",
48692=>"001000111",
48693=>"000000000",
48694=>"100111011",
48695=>"110000110",
48696=>"111111010",
48697=>"010000111",
48698=>"111010101",
48699=>"111000111",
48700=>"000000000",
48701=>"111010001",
48702=>"111000000",
48703=>"111111001",
48704=>"010000000",
48705=>"111000001",
48706=>"110111000",
48707=>"111000110",
48708=>"010000000",
48709=>"000001000",
48710=>"000111000",
48711=>"100000000",
48712=>"110000000",
48713=>"111000111",
48714=>"110110000",
48715=>"101010100",
48716=>"111000111",
48717=>"001011100",
48718=>"111111011",
48719=>"000000111",
48720=>"000000010",
48721=>"111011101",
48722=>"101010000",
48723=>"001001010",
48724=>"101000110",
48725=>"101001100",
48726=>"111110001",
48727=>"110000101",
48728=>"111010010",
48729=>"111111000",
48730=>"111110011",
48731=>"011111100",
48732=>"000111000",
48733=>"010000010",
48734=>"010111000",
48735=>"110000111",
48736=>"001001111",
48737=>"000111110",
48738=>"111000111",
48739=>"110111111",
48740=>"011000001",
48741=>"000010100",
48742=>"111001111",
48743=>"000011001",
48744=>"010000111",
48745=>"111010111",
48746=>"111111000",
48747=>"000000000",
48748=>"111101101",
48749=>"000011000",
48750=>"010111100",
48751=>"010011101",
48752=>"001000010",
48753=>"101000100",
48754=>"001111100",
48755=>"110110000",
48756=>"111011000",
48757=>"000001011",
48758=>"100010001",
48759=>"110001000",
48760=>"000111111",
48761=>"000111110",
48762=>"000000000",
48763=>"111000000",
48764=>"010000011",
48765=>"001001010",
48766=>"011111010",
48767=>"111000111",
48768=>"000100000",
48769=>"111000000",
48770=>"000000000",
48771=>"000111110",
48772=>"000100000",
48773=>"001000000",
48774=>"100101111",
48775=>"110000100",
48776=>"000000000",
48777=>"111000100",
48778=>"010111000",
48779=>"100000000",
48780=>"000111000",
48781=>"100111000",
48782=>"101000001",
48783=>"100000000",
48784=>"010000111",
48785=>"010000010",
48786=>"001111111",
48787=>"010111010",
48788=>"111100000",
48789=>"100110101",
48790=>"000000000",
48791=>"110010000",
48792=>"011101111",
48793=>"111111000",
48794=>"000000111",
48795=>"000000001",
48796=>"111111111",
48797=>"000111110",
48798=>"000111110",
48799=>"111000111",
48800=>"110000110",
48801=>"011010110",
48802=>"110111111",
48803=>"100000000",
48804=>"000111101",
48805=>"000000011",
48806=>"100000000",
48807=>"111111111",
48808=>"000000101",
48809=>"111011111",
48810=>"111000111",
48811=>"110010111",
48812=>"101111000",
48813=>"010111010",
48814=>"100000000",
48815=>"000111011",
48816=>"100100000",
48817=>"011000001",
48818=>"111111111",
48819=>"010001011",
48820=>"010000100",
48821=>"000000110",
48822=>"001000100",
48823=>"000000000",
48824=>"001000111",
48825=>"111001011",
48826=>"111111000",
48827=>"010000111",
48828=>"000111000",
48829=>"111111111",
48830=>"001111111",
48831=>"000100000",
48832=>"110010000",
48833=>"010000110",
48834=>"000100000",
48835=>"011101000",
48836=>"111000000",
48837=>"001000000",
48838=>"000110100",
48839=>"111111111",
48840=>"111111000",
48841=>"110000111",
48842=>"100111000",
48843=>"000000000",
48844=>"000010000",
48845=>"111100100",
48846=>"000000111",
48847=>"000001111",
48848=>"111011111",
48849=>"010011111",
48850=>"100101001",
48851=>"111000000",
48852=>"010010000",
48853=>"000000110",
48854=>"111000111",
48855=>"011011111",
48856=>"000000000",
48857=>"111111100",
48858=>"010111011",
48859=>"010010110",
48860=>"001110111",
48861=>"100010111",
48862=>"000000001",
48863=>"101101100",
48864=>"111110111",
48865=>"110000111",
48866=>"000000000",
48867=>"001010000",
48868=>"001101001",
48869=>"010000111",
48870=>"000011111",
48871=>"110001110",
48872=>"000100000",
48873=>"111111110",
48874=>"111000011",
48875=>"000000111",
48876=>"000000111",
48877=>"111111111",
48878=>"011011000",
48879=>"111101100",
48880=>"111111110",
48881=>"110000000",
48882=>"110110000",
48883=>"010111111",
48884=>"001111000",
48885=>"110000110",
48886=>"011000111",
48887=>"101000001",
48888=>"110110100",
48889=>"111111000",
48890=>"011000000",
48891=>"000001000",
48892=>"111111111",
48893=>"000111000",
48894=>"111101111",
48895=>"000010011",
48896=>"110110110",
48897=>"111100000",
48898=>"000000000",
48899=>"111001000",
48900=>"110110110",
48901=>"000000100",
48902=>"101111111",
48903=>"100100101",
48904=>"000000100",
48905=>"010111111",
48906=>"100010011",
48907=>"000000000",
48908=>"000000000",
48909=>"010000111",
48910=>"011110000",
48911=>"010001000",
48912=>"000000000",
48913=>"100000101",
48914=>"111100000",
48915=>"000110011",
48916=>"011000000",
48917=>"110111111",
48918=>"111011010",
48919=>"100100110",
48920=>"100000000",
48921=>"111111111",
48922=>"100100111",
48923=>"011011100",
48924=>"010100000",
48925=>"011111100",
48926=>"111001111",
48927=>"000000000",
48928=>"010111000",
48929=>"100000000",
48930=>"000000000",
48931=>"100000110",
48932=>"000000111",
48933=>"111100000",
48934=>"000000101",
48935=>"000000000",
48936=>"110111111",
48937=>"100001001",
48938=>"101111001",
48939=>"100000000",
48940=>"100100110",
48941=>"000000000",
48942=>"000111111",
48943=>"000100110",
48944=>"000000000",
48945=>"000110111",
48946=>"000110000",
48947=>"110111111",
48948=>"111001101",
48949=>"111011101",
48950=>"100000001",
48951=>"011011100",
48952=>"111100000",
48953=>"101000000",
48954=>"000000000",
48955=>"111100100",
48956=>"110111000",
48957=>"111111100",
48958=>"000000100",
48959=>"010011101",
48960=>"001001101",
48961=>"101111111",
48962=>"100101110",
48963=>"100000100",
48964=>"000010000",
48965=>"101001000",
48966=>"000111010",
48967=>"000000111",
48968=>"100100100",
48969=>"001000011",
48970=>"101100111",
48971=>"101100110",
48972=>"000100000",
48973=>"000000000",
48974=>"001001101",
48975=>"000000011",
48976=>"100000000",
48977=>"111110111",
48978=>"100110000",
48979=>"001000100",
48980=>"001000001",
48981=>"010111101",
48982=>"011011110",
48983=>"000000100",
48984=>"100000000",
48985=>"100110111",
48986=>"001011101",
48987=>"100110011",
48988=>"000100100",
48989=>"000001000",
48990=>"011111000",
48991=>"001001001",
48992=>"101100111",
48993=>"001111010",
48994=>"000000101",
48995=>"000100001",
48996=>"111111010",
48997=>"111110111",
48998=>"101111111",
48999=>"010110111",
49000=>"010011010",
49001=>"000010011",
49002=>"010011011",
49003=>"011110100",
49004=>"001000000",
49005=>"011111010",
49006=>"111100101",
49007=>"100000010",
49008=>"110110110",
49009=>"111101101",
49010=>"001100100",
49011=>"000000000",
49012=>"011111111",
49013=>"100000111",
49014=>"000000000",
49015=>"111111111",
49016=>"011011000",
49017=>"111111000",
49018=>"011111011",
49019=>"011101110",
49020=>"110110111",
49021=>"000000000",
49022=>"000110111",
49023=>"000001111",
49024=>"000101101",
49025=>"111100111",
49026=>"011010011",
49027=>"011111000",
49028=>"011111001",
49029=>"010111000",
49030=>"000011100",
49031=>"101100100",
49032=>"011011001",
49033=>"001000000",
49034=>"011011011",
49035=>"000100000",
49036=>"111111000",
49037=>"000000000",
49038=>"011011100",
49039=>"001000000",
49040=>"111111111",
49041=>"111101000",
49042=>"000000000",
49043=>"101100101",
49044=>"110010100",
49045=>"000000101",
49046=>"111011000",
49047=>"000011110",
49048=>"011010010",
49049=>"010000110",
49050=>"111111011",
49051=>"000000011",
49052=>"001000111",
49053=>"011011000",
49054=>"100100111",
49055=>"100100111",
49056=>"100100110",
49057=>"011011000",
49058=>"111101101",
49059=>"001111000",
49060=>"000101111",
49061=>"000000111",
49062=>"100010001",
49063=>"000000100",
49064=>"001111111",
49065=>"100010000",
49066=>"001100001",
49067=>"000100000",
49068=>"110100100",
49069=>"000000000",
49070=>"010001001",
49071=>"111111010",
49072=>"000101001",
49073=>"000100110",
49074=>"001101001",
49075=>"100000001",
49076=>"001011111",
49077=>"100100000",
49078=>"100100001",
49079=>"011111101",
49080=>"001001100",
49081=>"111010101",
49082=>"011001010",
49083=>"111100100",
49084=>"011111001",
49085=>"010011010",
49086=>"000100100",
49087=>"100000000",
49088=>"100000100",
49089=>"000100111",
49090=>"000111100",
49091=>"001101111",
49092=>"011110000",
49093=>"010110000",
49094=>"111011100",
49095=>"111111000",
49096=>"010100000",
49097=>"100000111",
49098=>"001101111",
49099=>"111111111",
49100=>"000100100",
49101=>"011011010",
49102=>"000001111",
49103=>"111111100",
49104=>"101100111",
49105=>"010110010",
49106=>"100001111",
49107=>"011001000",
49108=>"100100111",
49109=>"100001001",
49110=>"100000111",
49111=>"111011110",
49112=>"100000101",
49113=>"001111010",
49114=>"001001011",
49115=>"000010111",
49116=>"101000001",
49117=>"110010011",
49118=>"000100000",
49119=>"111011010",
49120=>"100000111",
49121=>"101100100",
49122=>"000000011",
49123=>"001111011",
49124=>"101000111",
49125=>"000000111",
49126=>"000100000",
49127=>"010110100",
49128=>"001100100",
49129=>"001000000",
49130=>"100100100",
49131=>"101100100",
49132=>"000000101",
49133=>"000010111",
49134=>"101100110",
49135=>"000100111",
49136=>"000000000",
49137=>"000011110",
49138=>"100100111",
49139=>"001111110",
49140=>"011011101",
49141=>"101111101",
49142=>"001000010",
49143=>"001001011",
49144=>"100000111",
49145=>"001011011",
49146=>"000000000",
49147=>"001111011",
49148=>"111111000",
49149=>"111111110",
49150=>"000000100",
49151=>"100100111",
49152=>"010000100",
49153=>"001110110",
49154=>"001001111",
49155=>"111000001",
49156=>"000000110",
49157=>"001000111",
49158=>"000000000",
49159=>"000000110",
49160=>"100101110",
49161=>"000000000",
49162=>"101000110",
49163=>"001000000",
49164=>"011001101",
49165=>"001001000",
49166=>"000110011",
49167=>"100010001",
49168=>"110110111",
49169=>"000011111",
49170=>"000000110",
49171=>"001110000",
49172=>"011001001",
49173=>"001000000",
49174=>"100000000",
49175=>"010111111",
49176=>"000000111",
49177=>"110010000",
49178=>"110110000",
49179=>"001000000",
49180=>"001000101",
49181=>"000000000",
49182=>"111000000",
49183=>"110110000",
49184=>"001111111",
49185=>"101110100",
49186=>"100101100",
49187=>"110110110",
49188=>"000000011",
49189=>"011111011",
49190=>"001000111",
49191=>"111111000",
49192=>"000001111",
49193=>"111001010",
49194=>"000100000",
49195=>"110111000",
49196=>"110111011",
49197=>"000000111",
49198=>"000101010",
49199=>"001000110",
49200=>"000000001",
49201=>"000000110",
49202=>"011111110",
49203=>"000001111",
49204=>"110000001",
49205=>"000001001",
49206=>"111111011",
49207=>"001000110",
49208=>"110000000",
49209=>"001000000",
49210=>"001000000",
49211=>"010100111",
49212=>"110011010",
49213=>"110111010",
49214=>"000000001",
49215=>"010111001",
49216=>"000110111",
49217=>"001111000",
49218=>"110111011",
49219=>"001110110",
49220=>"111010010",
49221=>"001000001",
49222=>"000000111",
49223=>"110000001",
49224=>"011111000",
49225=>"110110111",
49226=>"001000110",
49227=>"111110100",
49228=>"111000001",
49229=>"000100010",
49230=>"100010011",
49231=>"110110000",
49232=>"110000010",
49233=>"010010000",
49234=>"111111011",
49235=>"011000000",
49236=>"001001101",
49237=>"010010110",
49238=>"111010110",
49239=>"110110000",
49240=>"111000101",
49241=>"110010111",
49242=>"101101111",
49243=>"111110010",
49244=>"010110000",
49245=>"001001010",
49246=>"101101111",
49247=>"010110111",
49248=>"111000110",
49249=>"110110000",
49250=>"001001111",
49251=>"011001111",
49252=>"100000000",
49253=>"111011011",
49254=>"110110010",
49255=>"010111000",
49256=>"000010111",
49257=>"000000110",
49258=>"000100110",
49259=>"111110011",
49260=>"000000000",
49261=>"000001111",
49262=>"010010000",
49263=>"000001110",
49264=>"110111110",
49265=>"110110110",
49266=>"111110100",
49267=>"000000111",
49268=>"111111110",
49269=>"000000010",
49270=>"000010010",
49271=>"111001011",
49272=>"000001000",
49273=>"101110111",
49274=>"001110111",
49275=>"100001000",
49276=>"100110010",
49277=>"100000001",
49278=>"010110001",
49279=>"110010100",
49280=>"000000000",
49281=>"000000000",
49282=>"101000110",
49283=>"001101000",
49284=>"001000001",
49285=>"110001001",
49286=>"110110000",
49287=>"010100100",
49288=>"101101111",
49289=>"110000010",
49290=>"100101110",
49291=>"000000111",
49292=>"000010000",
49293=>"001001111",
49294=>"011001111",
49295=>"000000110",
49296=>"100000100",
49297=>"111111010",
49298=>"111110000",
49299=>"110000110",
49300=>"000110101",
49301=>"001001011",
49302=>"100100110",
49303=>"000001000",
49304=>"110111001",
49305=>"110110000",
49306=>"001001111",
49307=>"000000000",
49308=>"001000001",
49309=>"001001101",
49310=>"110000000",
49311=>"000010110",
49312=>"111001011",
49313=>"001001011",
49314=>"111110000",
49315=>"110100111",
49316=>"001000000",
49317=>"110000010",
49318=>"001010000",
49319=>"110111110",
49320=>"000000101",
49321=>"001100110",
49322=>"000000000",
49323=>"001001011",
49324=>"101110110",
49325=>"111001001",
49326=>"100010000",
49327=>"111111111",
49328=>"100111110",
49329=>"011001001",
49330=>"011001111",
49331=>"000100000",
49332=>"111111110",
49333=>"101111111",
49334=>"111111111",
49335=>"000101001",
49336=>"111110100",
49337=>"110110010",
49338=>"010111110",
49339=>"111000101",
49340=>"000000000",
49341=>"011011111",
49342=>"110000010",
49343=>"111111000",
49344=>"000000001",
49345=>"111000000",
49346=>"110010110",
49347=>"001000010",
49348=>"100001001",
49349=>"100000000",
49350=>"001111110",
49351=>"001101111",
49352=>"111001100",
49353=>"110110000",
49354=>"110001110",
49355=>"110110000",
49356=>"110110010",
49357=>"011010100",
49358=>"000000001",
49359=>"000110110",
49360=>"000000011",
49361=>"110110110",
49362=>"010010100",
49363=>"110111110",
49364=>"000000001",
49365=>"100100110",
49366=>"101001110",
49367=>"001000000",
49368=>"111000000",
49369=>"000110000",
49370=>"100100001",
49371=>"000000111",
49372=>"000000111",
49373=>"111101100",
49374=>"110000000",
49375=>"110000000",
49376=>"000110010",
49377=>"001000111",
49378=>"000000000",
49379=>"101100111",
49380=>"110110000",
49381=>"101001001",
49382=>"000001100",
49383=>"010000000",
49384=>"110110100",
49385=>"001001101",
49386=>"001011001",
49387=>"000000011",
49388=>"110110110",
49389=>"110001100",
49390=>"010011000",
49391=>"000000000",
49392=>"110110000",
49393=>"011001000",
49394=>"000000001",
49395=>"100100000",
49396=>"000001001",
49397=>"101111111",
49398=>"000000110",
49399=>"000000000",
49400=>"000000001",
49401=>"000001011",
49402=>"001001011",
49403=>"000001111",
49404=>"111001010",
49405=>"110110000",
49406=>"011011110",
49407=>"000010110",
49408=>"011001000",
49409=>"000011010",
49410=>"100000000",
49411=>"100101011",
49412=>"001111111",
49413=>"011000000",
49414=>"100110110",
49415=>"000011111",
49416=>"000100111",
49417=>"000100000",
49418=>"100000001",
49419=>"101100111",
49420=>"011011001",
49421=>"111101101",
49422=>"000010111",
49423=>"000100111",
49424=>"000111011",
49425=>"100101111",
49426=>"000110000",
49427=>"110001011",
49428=>"111111111",
49429=>"110101100",
49430=>"000001000",
49431=>"101110010",
49432=>"000000000",
49433=>"111111101",
49434=>"011101010",
49435=>"000100101",
49436=>"101011011",
49437=>"101100000",
49438=>"110000000",
49439=>"000111000",
49440=>"000101101",
49441=>"000111001",
49442=>"001011010",
49443=>"011111000",
49444=>"111111110",
49445=>"011000000",
49446=>"111100100",
49447=>"000000000",
49448=>"011111111",
49449=>"001110010",
49450=>"100000011",
49451=>"010010000",
49452=>"000001110",
49453=>"111111111",
49454=>"111110000",
49455=>"000001000",
49456=>"111000000",
49457=>"110110011",
49458=>"111101000",
49459=>"000011011",
49460=>"000000000",
49461=>"010111010",
49462=>"110000001",
49463=>"100100100",
49464=>"111000000",
49465=>"000000101",
49466=>"000000100",
49467=>"010010011",
49468=>"110110100",
49469=>"111111000",
49470=>"010000000",
49471=>"100000000",
49472=>"101100111",
49473=>"011000011",
49474=>"000100100",
49475=>"001100100",
49476=>"110011000",
49477=>"101100011",
49478=>"000010000",
49479=>"111010010",
49480=>"101101101",
49481=>"000000000",
49482=>"101000011",
49483=>"011011011",
49484=>"100000000",
49485=>"010010011",
49486=>"011011111",
49487=>"001011101",
49488=>"100101000",
49489=>"111101111",
49490=>"110100011",
49491=>"011000001",
49492=>"010100000",
49493=>"100111101",
49494=>"011000000",
49495=>"000110010",
49496=>"110100001",
49497=>"000001001",
49498=>"110110000",
49499=>"010010011",
49500=>"111010000",
49501=>"001001001",
49502=>"000011111",
49503=>"000000000",
49504=>"111011000",
49505=>"101111111",
49506=>"000000100",
49507=>"100100000",
49508=>"000000100",
49509=>"100110000",
49510=>"000001000",
49511=>"011000100",
49512=>"010000101",
49513=>"000000111",
49514=>"010111011",
49515=>"100000010",
49516=>"111010000",
49517=>"000000000",
49518=>"011100000",
49519=>"011010100",
49520=>"001110111",
49521=>"000000101",
49522=>"001010111",
49523=>"000011011",
49524=>"010010011",
49525=>"100000000",
49526=>"000111111",
49527=>"011011000",
49528=>"000010010",
49529=>"001000011",
49530=>"000111111",
49531=>"000011001",
49532=>"101110011",
49533=>"100000000",
49534=>"111000100",
49535=>"000000100",
49536=>"111001010",
49537=>"111011000",
49538=>"100100010",
49539=>"111101000",
49540=>"000000011",
49541=>"111101111",
49542=>"011000100",
49543=>"000011001",
49544=>"010001111",
49545=>"111111111",
49546=>"111000000",
49547=>"110000010",
49548=>"000100101",
49549=>"100100111",
49550=>"000000100",
49551=>"000000001",
49552=>"000000111",
49553=>"000000000",
49554=>"000000000",
49555=>"000011111",
49556=>"000011101",
49557=>"000000111",
49558=>"110000101",
49559=>"100001111",
49560=>"000011011",
49561=>"000000111",
49562=>"111100000",
49563=>"000000111",
49564=>"100000000",
49565=>"010000101",
49566=>"111111011",
49567=>"111010000",
49568=>"101011000",
49569=>"100000010",
49570=>"001000000",
49571=>"011000000",
49572=>"000000000",
49573=>"100110110",
49574=>"000110000",
49575=>"110111011",
49576=>"000010111",
49577=>"000010011",
49578=>"110000101",
49579=>"000011000",
49580=>"101111101",
49581=>"100100011",
49582=>"001001111",
49583=>"011111101",
49584=>"000000000",
49585=>"001000110",
49586=>"100001111",
49587=>"000100001",
49588=>"000000000",
49589=>"111111111",
49590=>"011011011",
49591=>"011011000",
49592=>"001010000",
49593=>"001111111",
49594=>"011111010",
49595=>"111100000",
49596=>"011001000",
49597=>"111111000",
49598=>"001000001",
49599=>"000000001",
49600=>"100000000",
49601=>"111000111",
49602=>"000000011",
49603=>"000110000",
49604=>"000011000",
49605=>"110111101",
49606=>"101000010",
49607=>"010011000",
49608=>"101111000",
49609=>"111100110",
49610=>"111111011",
49611=>"001011011",
49612=>"110000100",
49613=>"101011010",
49614=>"011111010",
49615=>"100110001",
49616=>"110101111",
49617=>"001000110",
49618=>"010000100",
49619=>"100011011",
49620=>"000000100",
49621=>"110011001",
49622=>"100000000",
49623=>"000011000",
49624=>"111111000",
49625=>"011101111",
49626=>"011011010",
49627=>"000000110",
49628=>"111100000",
49629=>"011000011",
49630=>"011100110",
49631=>"000000000",
49632=>"000011000",
49633=>"100000100",
49634=>"000100111",
49635=>"010100111",
49636=>"101000000",
49637=>"110101000",
49638=>"111101110",
49639=>"010000010",
49640=>"100101111",
49641=>"101101000",
49642=>"000100000",
49643=>"100111001",
49644=>"000100111",
49645=>"001011111",
49646=>"000100000",
49647=>"010010000",
49648=>"100110111",
49649=>"001111100",
49650=>"100100000",
49651=>"100000110",
49652=>"110111101",
49653=>"100111100",
49654=>"000111000",
49655=>"001000000",
49656=>"000001111",
49657=>"101101110",
49658=>"011011010",
49659=>"100100011",
49660=>"010001000",
49661=>"101001001",
49662=>"111111011",
49663=>"000000000",
49664=>"001001010",
49665=>"000111011",
49666=>"101001101",
49667=>"001001010",
49668=>"110100110",
49669=>"000000101",
49670=>"111101101",
49671=>"111101000",
49672=>"110000000",
49673=>"000000100",
49674=>"111111001",
49675=>"011000000",
49676=>"000000100",
49677=>"010011110",
49678=>"010011010",
49679=>"111111111",
49680=>"110000100",
49681=>"100000101",
49682=>"010111011",
49683=>"001000001",
49684=>"101101101",
49685=>"001000011",
49686=>"111111011",
49687=>"001000010",
49688=>"101100000",
49689=>"111101100",
49690=>"110000000",
49691=>"000000000",
49692=>"111111010",
49693=>"001000100",
49694=>"111111111",
49695=>"011110010",
49696=>"011111001",
49697=>"000000001",
49698=>"001010111",
49699=>"000000000",
49700=>"100100100",
49701=>"000001111",
49702=>"111010010",
49703=>"000100100",
49704=>"110111000",
49705=>"101001101",
49706=>"101101111",
49707=>"000111111",
49708=>"010101100",
49709=>"111111001",
49710=>"001000101",
49711=>"111001000",
49712=>"110011000",
49713=>"111100000",
49714=>"000110011",
49715=>"111101101",
49716=>"001001000",
49717=>"011001001",
49718=>"000000111",
49719=>"100000100",
49720=>"010101000",
49721=>"000000100",
49722=>"101101111",
49723=>"011000000",
49724=>"011011000",
49725=>"011111011",
49726=>"000000000",
49727=>"110110100",
49728=>"101000101",
49729=>"000111110",
49730=>"010000000",
49731=>"011001000",
49732=>"111111010",
49733=>"100100000",
49734=>"010111000",
49735=>"010010001",
49736=>"001011011",
49737=>"111001001",
49738=>"000101101",
49739=>"110000110",
49740=>"000000111",
49741=>"001010000",
49742=>"111011001",
49743=>"111101100",
49744=>"000010010",
49745=>"000110110",
49746=>"111111101",
49747=>"111100000",
49748=>"000000110",
49749=>"100001011",
49750=>"011011001",
49751=>"000100101",
49752=>"000111011",
49753=>"100100101",
49754=>"101001011",
49755=>"100001111",
49756=>"111001000",
49757=>"101001101",
49758=>"000111111",
49759=>"001000000",
49760=>"111111010",
49761=>"010000000",
49762=>"111111101",
49763=>"001100000",
49764=>"111111000",
49765=>"100111110",
49766=>"010011111",
49767=>"111011011",
49768=>"010111011",
49769=>"101100100",
49770=>"000010010",
49771=>"111111000",
49772=>"111101101",
49773=>"100110111",
49774=>"111010010",
49775=>"000100101",
49776=>"110110000",
49777=>"000001000",
49778=>"000100000",
49779=>"111000100",
49780=>"101111011",
49781=>"000000111",
49782=>"000001101",
49783=>"110000000",
49784=>"000001111",
49785=>"011011001",
49786=>"100110000",
49787=>"000000000",
49788=>"111000000",
49789=>"110000000",
49790=>"010010111",
49791=>"101000001",
49792=>"101101111",
49793=>"100010000",
49794=>"111100010",
49795=>"111011000",
49796=>"001000000",
49797=>"010000000",
49798=>"100110110",
49799=>"000000111",
49800=>"111001000",
49801=>"000101101",
49802=>"100111101",
49803=>"111000100",
49804=>"110111111",
49805=>"001000100",
49806=>"000011111",
49807=>"001001101",
49808=>"100110110",
49809=>"010110011",
49810=>"101000010",
49811=>"110000000",
49812=>"011011001",
49813=>"100000100",
49814=>"000000101",
49815=>"001011001",
49816=>"010110110",
49817=>"000010111",
49818=>"010000110",
49819=>"000100000",
49820=>"001101100",
49821=>"110111101",
49822=>"100000000",
49823=>"000000101",
49824=>"100100110",
49825=>"101101000",
49826=>"111000000",
49827=>"000100111",
49828=>"000000101",
49829=>"111001011",
49830=>"111010000",
49831=>"000000110",
49832=>"010000001",
49833=>"110110111",
49834=>"000100000",
49835=>"000000000",
49836=>"010000000",
49837=>"111111000",
49838=>"000011001",
49839=>"111010000",
49840=>"000010011",
49841=>"010001001",
49842=>"100100111",
49843=>"000010110",
49844=>"011011110",
49845=>"110101111",
49846=>"111100000",
49847=>"010111000",
49848=>"101100000",
49849=>"011000000",
49850=>"010010010",
49851=>"000101111",
49852=>"100000110",
49853=>"010111011",
49854=>"101001000",
49855=>"000101000",
49856=>"101001101",
49857=>"101100100",
49858=>"100110110",
49859=>"110100100",
49860=>"111101111",
49861=>"111110000",
49862=>"011011101",
49863=>"000000111",
49864=>"010000110",
49865=>"001000010",
49866=>"101111101",
49867=>"111111110",
49868=>"001000000",
49869=>"110110000",
49870=>"100000011",
49871=>"000001111",
49872=>"101001000",
49873=>"110110100",
49874=>"111101100",
49875=>"011000100",
49876=>"000000100",
49877=>"000100110",
49878=>"100100000",
49879=>"101110011",
49880=>"100101111",
49881=>"001010000",
49882=>"011000000",
49883=>"000000111",
49884=>"111011100",
49885=>"111010010",
49886=>"101001010",
49887=>"111111000",
49888=>"111000000",
49889=>"111110110",
49890=>"101111110",
49891=>"110110000",
49892=>"111111111",
49893=>"101000000",
49894=>"011000000",
49895=>"000100100",
49896=>"000000000",
49897=>"101111000",
49898=>"100100000",
49899=>"100000010",
49900=>"000000010",
49901=>"111111110",
49902=>"001000000",
49903=>"111010001",
49904=>"111000000",
49905=>"011011101",
49906=>"111000000",
49907=>"110011010",
49908=>"100011101",
49909=>"100010010",
49910=>"000000000",
49911=>"100111111",
49912=>"000000111",
49913=>"100001111",
49914=>"000000000",
49915=>"111111100",
49916=>"111111110",
49917=>"011111010",
49918=>"000000000",
49919=>"000101101",
49920=>"111111111",
49921=>"111011100",
49922=>"100100110",
49923=>"010100001",
49924=>"111110111",
49925=>"110000101",
49926=>"101000101",
49927=>"000111111",
49928=>"011001001",
49929=>"000000001",
49930=>"001010000",
49931=>"000000000",
49932=>"000100000",
49933=>"000000100",
49934=>"101100010",
49935=>"100111110",
49936=>"000000000",
49937=>"110010011",
49938=>"111111011",
49939=>"000101010",
49940=>"010111111",
49941=>"100111010",
49942=>"000001101",
49943=>"101111010",
49944=>"100000000",
49945=>"111111111",
49946=>"111100100",
49947=>"000000100",
49948=>"110100111",
49949=>"010111000",
49950=>"111100011",
49951=>"001000000",
49952=>"111000001",
49953=>"010100010",
49954=>"000000010",
49955=>"111100000",
49956=>"100110100",
49957=>"011111111",
49958=>"111110000",
49959=>"000000101",
49960=>"111101000",
49961=>"000000000",
49962=>"000000000",
49963=>"111010111",
49964=>"000110000",
49965=>"111011010",
49966=>"011011110",
49967=>"111100011",
49968=>"010010101",
49969=>"011110111",
49970=>"101101111",
49971=>"010111011",
49972=>"000111111",
49973=>"001111111",
49974=>"000011010",
49975=>"000111111",
49976=>"010101111",
49977=>"101111111",
49978=>"011101101",
49979=>"000001111",
49980=>"011111111",
49981=>"111111010",
49982=>"101000001",
49983=>"101001011",
49984=>"111111101",
49985=>"101111101",
49986=>"000000011",
49987=>"100101110",
49988=>"001000000",
49989=>"000101111",
49990=>"000100000",
49991=>"000110001",
49992=>"001111001",
49993=>"010001100",
49994=>"001100000",
49995=>"011110111",
49996=>"111111111",
49997=>"000111111",
49998=>"000001001",
49999=>"000111111",
50000=>"000100111",
50001=>"111111110",
50002=>"101100101",
50003=>"001101100",
50004=>"000000000",
50005=>"001110110",
50006=>"010001000",
50007=>"101000101",
50008=>"000000000",
50009=>"101110001",
50010=>"101000000",
50011=>"111011111",
50012=>"110110000",
50013=>"010000001",
50014=>"000000111",
50015=>"101101101",
50016=>"001000101",
50017=>"111000000",
50018=>"000000100",
50019=>"000100000",
50020=>"000101100",
50021=>"111100000",
50022=>"110101111",
50023=>"100101111",
50024=>"000100111",
50025=>"111101111",
50026=>"000000000",
50027=>"111111100",
50028=>"000111101",
50029=>"000111000",
50030=>"000100101",
50031=>"100000010",
50032=>"000001101",
50033=>"111011000",
50034=>"111011011",
50035=>"111001010",
50036=>"000101011",
50037=>"000001111",
50038=>"111000000",
50039=>"001010001",
50040=>"000001000",
50041=>"010000001",
50042=>"010000101",
50043=>"000000000",
50044=>"110000010",
50045=>"111110011",
50046=>"010101111",
50047=>"101000000",
50048=>"110110101",
50049=>"000000010",
50050=>"000010111",
50051=>"000010010",
50052=>"000011010",
50053=>"011000010",
50054=>"100111110",
50055=>"111111011",
50056=>"000100111",
50057=>"000010011",
50058=>"111001000",
50059=>"010001010",
50060=>"000101101",
50061=>"000000101",
50062=>"010111111",
50063=>"011000000",
50064=>"111111011",
50065=>"011110001",
50066=>"010000011",
50067=>"111000000",
50068=>"110111111",
50069=>"100101101",
50070=>"110111010",
50071=>"010100100",
50072=>"001010100",
50073=>"101111101",
50074=>"010010110",
50075=>"100000000",
50076=>"101000000",
50077=>"000000101",
50078=>"011011010",
50079=>"111101111",
50080=>"100111010",
50081=>"110011111",
50082=>"011000000",
50083=>"111000000",
50084=>"011000010",
50085=>"111111010",
50086=>"110001011",
50087=>"000000010",
50088=>"110010010",
50089=>"000000011",
50090=>"011111111",
50091=>"100100111",
50092=>"010011101",
50093=>"111000100",
50094=>"011111101",
50095=>"100000010",
50096=>"000000001",
50097=>"100000100",
50098=>"110111000",
50099=>"111001000",
50100=>"101111001",
50101=>"111010010",
50102=>"111111000",
50103=>"110000011",
50104=>"111011001",
50105=>"101111011",
50106=>"011011011",
50107=>"010110000",
50108=>"000100000",
50109=>"000000000",
50110=>"100000100",
50111=>"000000101",
50112=>"111000000",
50113=>"010111011",
50114=>"110110000",
50115=>"000001000",
50116=>"010010000",
50117=>"000111100",
50118=>"111111100",
50119=>"111100011",
50120=>"000000000",
50121=>"000000000",
50122=>"000000011",
50123=>"000111111",
50124=>"111000000",
50125=>"001010110",
50126=>"111010010",
50127=>"011111111",
50128=>"101000000",
50129=>"001111111",
50130=>"110110111",
50131=>"001101111",
50132=>"000101010",
50133=>"111110110",
50134=>"101000001",
50135=>"000000011",
50136=>"111111000",
50137=>"000000000",
50138=>"011100100",
50139=>"111100101",
50140=>"100101111",
50141=>"100101100",
50142=>"001010000",
50143=>"100000101",
50144=>"111000000",
50145=>"111000001",
50146=>"000000000",
50147=>"101111111",
50148=>"111000000",
50149=>"111100101",
50150=>"100000000",
50151=>"111010110",
50152=>"100100000",
50153=>"001100100",
50154=>"110011010",
50155=>"111100101",
50156=>"000000000",
50157=>"111001101",
50158=>"111101000",
50159=>"000000000",
50160=>"000000011",
50161=>"001111000",
50162=>"001001100",
50163=>"100001111",
50164=>"001110111",
50165=>"100001011",
50166=>"110000000",
50167=>"111001011",
50168=>"010000000",
50169=>"010111010",
50170=>"100000101",
50171=>"011110111",
50172=>"111111111",
50173=>"111101111",
50174=>"000011011",
50175=>"110111111",
50176=>"101101110",
50177=>"111111111",
50178=>"011010101",
50179=>"000000011",
50180=>"011011011",
50181=>"010111000",
50182=>"101000000",
50183=>"100110000",
50184=>"110111100",
50185=>"000001001",
50186=>"001111111",
50187=>"010100000",
50188=>"011110000",
50189=>"000100111",
50190=>"110100001",
50191=>"000000001",
50192=>"100000000",
50193=>"101111111",
50194=>"111110000",
50195=>"001000000",
50196=>"111111111",
50197=>"000011011",
50198=>"110101111",
50199=>"010010011",
50200=>"000000111",
50201=>"001011000",
50202=>"111111111",
50203=>"011000000",
50204=>"000100100",
50205=>"011001100",
50206=>"011011010",
50207=>"001101111",
50208=>"100110000",
50209=>"100111111",
50210=>"111101001",
50211=>"011000000",
50212=>"010000000",
50213=>"000000011",
50214=>"000011111",
50215=>"000000000",
50216=>"000011111",
50217=>"000111111",
50218=>"100001111",
50219=>"000101000",
50220=>"000001001",
50221=>"101110111",
50222=>"110011111",
50223=>"000000000",
50224=>"000110111",
50225=>"001000000",
50226=>"101110100",
50227=>"010111000",
50228=>"111011001",
50229=>"100001111",
50230=>"010111111",
50231=>"001000000",
50232=>"010111010",
50233=>"111100000",
50234=>"100000000",
50235=>"111000001",
50236=>"001011110",
50237=>"110111111",
50238=>"100000000",
50239=>"111010110",
50240=>"111111000",
50241=>"000000000",
50242=>"100011100",
50243=>"101000000",
50244=>"000111111",
50245=>"000100100",
50246=>"101000000",
50247=>"001001101",
50248=>"001110000",
50249=>"000100100",
50250=>"000000000",
50251=>"000000100",
50252=>"100000000",
50253=>"000000000",
50254=>"111110000",
50255=>"111001111",
50256=>"000010011",
50257=>"111011101",
50258=>"011001000",
50259=>"100111000",
50260=>"001000000",
50261=>"011111111",
50262=>"010011000",
50263=>"001000000",
50264=>"101000100",
50265=>"001101001",
50266=>"110111111",
50267=>"010110110",
50268=>"000010100",
50269=>"111111010",
50270=>"000011111",
50271=>"001000011",
50272=>"101000000",
50273=>"000000000",
50274=>"000000100",
50275=>"011101001",
50276=>"000111111",
50277=>"111111100",
50278=>"100000000",
50279=>"111111111",
50280=>"111111111",
50281=>"001000111",
50282=>"010111111",
50283=>"001110000",
50284=>"111110000",
50285=>"000011111",
50286=>"010000100",
50287=>"110000000",
50288=>"111110111",
50289=>"111111011",
50290=>"101111011",
50291=>"111100000",
50292=>"000011110",
50293=>"000000100",
50294=>"111111010",
50295=>"000111010",
50296=>"001111111",
50297=>"000000000",
50298=>"101010111",
50299=>"011000101",
50300=>"111011010",
50301=>"011111001",
50302=>"001111111",
50303=>"000000000",
50304=>"000000000",
50305=>"011111111",
50306=>"000000111",
50307=>"000000000",
50308=>"011000000",
50309=>"111101001",
50310=>"000000000",
50311=>"001000000",
50312=>"110011001",
50313=>"111100100",
50314=>"111100100",
50315=>"001001000",
50316=>"000000101",
50317=>"010011111",
50318=>"000000000",
50319=>"100000000",
50320=>"000000000",
50321=>"011010000",
50322=>"000011111",
50323=>"111111000",
50324=>"110010010",
50325=>"110111000",
50326=>"111100100",
50327=>"011000000",
50328=>"000110000",
50329=>"000111001",
50330=>"111000000",
50331=>"111000000",
50332=>"111101000",
50333=>"111000000",
50334=>"011010000",
50335=>"111000000",
50336=>"110100010",
50337=>"111111000",
50338=>"000000111",
50339=>"001000000",
50340=>"010111011",
50341=>"000000010",
50342=>"010011111",
50343=>"111101100",
50344=>"101011101",
50345=>"100000011",
50346=>"110000000",
50347=>"000000110",
50348=>"101000001",
50349=>"000000110",
50350=>"000010001",
50351=>"100000001",
50352=>"100000000",
50353=>"100110000",
50354=>"000000101",
50355=>"111110110",
50356=>"000111000",
50357=>"101000111",
50358=>"000010111",
50359=>"000000000",
50360=>"110101011",
50361=>"111001000",
50362=>"000000010",
50363=>"000100110",
50364=>"011001010",
50365=>"011111011",
50366=>"111111110",
50367=>"101111101",
50368=>"000000000",
50369=>"100000100",
50370=>"011011000",
50371=>"110110110",
50372=>"111000100",
50373=>"101110111",
50374=>"101000011",
50375=>"010000000",
50376=>"111111100",
50377=>"111101101",
50378=>"000111111",
50379=>"110000111",
50380=>"000000000",
50381=>"111110101",
50382=>"101101111",
50383=>"010111000",
50384=>"011010010",
50385=>"000100000",
50386=>"000000000",
50387=>"000000000",
50388=>"111000100",
50389=>"001011011",
50390=>"111000000",
50391=>"000001011",
50392=>"101000000",
50393=>"111101111",
50394=>"111011001",
50395=>"000100100",
50396=>"011011010",
50397=>"000000111",
50398=>"100000000",
50399=>"001010001",
50400=>"010110100",
50401=>"001010100",
50402=>"111111011",
50403=>"111100000",
50404=>"000000100",
50405=>"111000000",
50406=>"111000000",
50407=>"000011100",
50408=>"000111111",
50409=>"000111110",
50410=>"000110011",
50411=>"100100000",
50412=>"111010000",
50413=>"111101000",
50414=>"010010111",
50415=>"011011000",
50416=>"111101000",
50417=>"001011111",
50418=>"010000000",
50419=>"110111111",
50420=>"000111011",
50421=>"111000101",
50422=>"100000000",
50423=>"001001001",
50424=>"000111011",
50425=>"101111110",
50426=>"000011000",
50427=>"010000000",
50428=>"101000000",
50429=>"001000000",
50430=>"000100110",
50431=>"111000000",
50432=>"011000000",
50433=>"010110011",
50434=>"001000000",
50435=>"110001111",
50436=>"111111011",
50437=>"111110000",
50438=>"110111110",
50439=>"111111111",
50440=>"111001000",
50441=>"111001101",
50442=>"100100010",
50443=>"000000000",
50444=>"111111101",
50445=>"011111001",
50446=>"011000111",
50447=>"000011100",
50448=>"110111010",
50449=>"000000100",
50450=>"111000111",
50451=>"111000000",
50452=>"111101100",
50453=>"111111000",
50454=>"000000000",
50455=>"111101111",
50456=>"010110010",
50457=>"111011000",
50458=>"101111011",
50459=>"000111111",
50460=>"011010010",
50461=>"101001001",
50462=>"111000100",
50463=>"000011111",
50464=>"000000000",
50465=>"111111111",
50466=>"000001001",
50467=>"000111101",
50468=>"000000111",
50469=>"111001000",
50470=>"111100000",
50471=>"000000000",
50472=>"101111001",
50473=>"101111111",
50474=>"111000101",
50475=>"000111110",
50476=>"001111011",
50477=>"111110111",
50478=>"111111000",
50479=>"100111111",
50480=>"111111111",
50481=>"001001000",
50482=>"000000001",
50483=>"110111110",
50484=>"000000000",
50485=>"010001100",
50486=>"000000000",
50487=>"111001000",
50488=>"111000000",
50489=>"101000111",
50490=>"000110111",
50491=>"000000010",
50492=>"100001000",
50493=>"111111011",
50494=>"010000110",
50495=>"000100100",
50496=>"000000000",
50497=>"110010000",
50498=>"111111111",
50499=>"100000000",
50500=>"111111000",
50501=>"111111101",
50502=>"000000000",
50503=>"010110000",
50504=>"110001010",
50505=>"111111000",
50506=>"111111111",
50507=>"000000010",
50508=>"111111111",
50509=>"100100000",
50510=>"110110110",
50511=>"011111111",
50512=>"001101101",
50513=>"000110101",
50514=>"111110111",
50515=>"111010000",
50516=>"000000000",
50517=>"000000000",
50518=>"110110000",
50519=>"111011111",
50520=>"010011000",
50521=>"010010111",
50522=>"100101100",
50523=>"000000011",
50524=>"000110110",
50525=>"010011011",
50526=>"000000000",
50527=>"001000000",
50528=>"111001111",
50529=>"001011110",
50530=>"101101101",
50531=>"000111110",
50532=>"111111111",
50533=>"100100110",
50534=>"111111011",
50535=>"111000000",
50536=>"011010010",
50537=>"110111110",
50538=>"110110100",
50539=>"000110010",
50540=>"100101101",
50541=>"111111111",
50542=>"111010000",
50543=>"010010010",
50544=>"000000101",
50545=>"110010010",
50546=>"000000000",
50547=>"111111111",
50548=>"011000111",
50549=>"101000000",
50550=>"111111010",
50551=>"000111111",
50552=>"001100111",
50553=>"100000101",
50554=>"000001111",
50555=>"111101111",
50556=>"000000000",
50557=>"111101100",
50558=>"000000111",
50559=>"101111101",
50560=>"001001001",
50561=>"000000000",
50562=>"110000101",
50563=>"010110100",
50564=>"010011000",
50565=>"000000011",
50566=>"111010010",
50567=>"011011011",
50568=>"001111000",
50569=>"000100000",
50570=>"011010010",
50571=>"000111001",
50572=>"111001000",
50573=>"001000110",
50574=>"111011101",
50575=>"110100000",
50576=>"011101111",
50577=>"000000000",
50578=>"010000010",
50579=>"010000010",
50580=>"000110110",
50581=>"111110111",
50582=>"111000000",
50583=>"101101100",
50584=>"111111001",
50585=>"111111110",
50586=>"101110111",
50587=>"101111111",
50588=>"111000010",
50589=>"000000000",
50590=>"011011000",
50591=>"000110100",
50592=>"001000011",
50593=>"010000111",
50594=>"111111111",
50595=>"111000000",
50596=>"110100000",
50597=>"101111111",
50598=>"111111101",
50599=>"111001001",
50600=>"110000111",
50601=>"011001011",
50602=>"000000101",
50603=>"001110111",
50604=>"000000101",
50605=>"111111000",
50606=>"000000000",
50607=>"100111111",
50608=>"000000001",
50609=>"100101111",
50610=>"111111111",
50611=>"100000000",
50612=>"100101110",
50613=>"111111010",
50614=>"001000100",
50615=>"101111100",
50616=>"001000000",
50617=>"000111111",
50618=>"111111111",
50619=>"010111111",
50620=>"111111010",
50621=>"001100101",
50622=>"011000101",
50623=>"000111000",
50624=>"000000000",
50625=>"011111110",
50626=>"111110001",
50627=>"101111011",
50628=>"111111111",
50629=>"000000100",
50630=>"010111011",
50631=>"101100111",
50632=>"111000101",
50633=>"000011001",
50634=>"110111100",
50635=>"111001000",
50636=>"101000011",
50637=>"000000000",
50638=>"000000000",
50639=>"000001101",
50640=>"100110110",
50641=>"010100010",
50642=>"010101001",
50643=>"110011111",
50644=>"000000000",
50645=>"010110000",
50646=>"000000000",
50647=>"111001111",
50648=>"000000000",
50649=>"000000000",
50650=>"100000000",
50651=>"111111110",
50652=>"000000000",
50653=>"111111011",
50654=>"000011010",
50655=>"111101111",
50656=>"111111010",
50657=>"101111111",
50658=>"000000101",
50659=>"100100000",
50660=>"000111111",
50661=>"101011111",
50662=>"111111111",
50663=>"000000001",
50664=>"111001000",
50665=>"010010111",
50666=>"000010001",
50667=>"000111001",
50668=>"101001111",
50669=>"000101101",
50670=>"001001001",
50671=>"110111001",
50672=>"000000001",
50673=>"010000010",
50674=>"111001110",
50675=>"110110110",
50676=>"010001000",
50677=>"000111001",
50678=>"111000011",
50679=>"000000010",
50680=>"111000000",
50681=>"010111111",
50682=>"111000010",
50683=>"000000001",
50684=>"111000000",
50685=>"111000000",
50686=>"111111101",
50687=>"100000000",
50688=>"000111011",
50689=>"010000101",
50690=>"000011110",
50691=>"110000000",
50692=>"011100100",
50693=>"010000110",
50694=>"101000000",
50695=>"111010111",
50696=>"000000001",
50697=>"010000000",
50698=>"000000000",
50699=>"101111100",
50700=>"111000000",
50701=>"011000000",
50702=>"011100100",
50703=>"011000000",
50704=>"101110000",
50705=>"110000000",
50706=>"001101100",
50707=>"000000101",
50708=>"000011111",
50709=>"010000010",
50710=>"100111011",
50711=>"100000000",
50712=>"111101000",
50713=>"010111111",
50714=>"001000000",
50715=>"011110110",
50716=>"100111011",
50717=>"111111011",
50718=>"010000001",
50719=>"010111111",
50720=>"100010110",
50721=>"111111111",
50722=>"111000100",
50723=>"000000010",
50724=>"001001101",
50725=>"000100100",
50726=>"010010010",
50727=>"010000000",
50728=>"011010010",
50729=>"101000001",
50730=>"010000000",
50731=>"110111100",
50732=>"111101101",
50733=>"111110000",
50734=>"110111001",
50735=>"111110011",
50736=>"101000000",
50737=>"101101100",
50738=>"000001111",
50739=>"100110110",
50740=>"000000000",
50741=>"011110110",
50742=>"001000100",
50743=>"000001111",
50744=>"111000000",
50745=>"100100000",
50746=>"000101001",
50747=>"000010101",
50748=>"001011111",
50749=>"111111111",
50750=>"000000000",
50751=>"001100111",
50752=>"000001100",
50753=>"010000110",
50754=>"101101001",
50755=>"001000100",
50756=>"111000100",
50757=>"010011101",
50758=>"000000000",
50759=>"010000100",
50760=>"101100000",
50761=>"111110111",
50762=>"101100000",
50763=>"111001010",
50764=>"010000000",
50765=>"001100000",
50766=>"011011001",
50767=>"100110000",
50768=>"000000101",
50769=>"000000000",
50770=>"110000111",
50771=>"110110001",
50772=>"011010000",
50773=>"100001001",
50774=>"000000101",
50775=>"000000000",
50776=>"101001001",
50777=>"100101100",
50778=>"000001111",
50779=>"111001000",
50780=>"010100000",
50781=>"001101001",
50782=>"000000110",
50783=>"101001000",
50784=>"101111111",
50785=>"010001100",
50786=>"101000101",
50787=>"000001101",
50788=>"110111000",
50789=>"011111111",
50790=>"110111111",
50791=>"010101110",
50792=>"111010111",
50793=>"010000000",
50794=>"110100101",
50795=>"000000000",
50796=>"101001001",
50797=>"111111000",
50798=>"010000000",
50799=>"000111101",
50800=>"111111100",
50801=>"111000000",
50802=>"100100001",
50803=>"010101000",
50804=>"000001101",
50805=>"000001000",
50806=>"111010000",
50807=>"000110111",
50808=>"000000111",
50809=>"100011111",
50810=>"111101111",
50811=>"101111010",
50812=>"110011000",
50813=>"001001100",
50814=>"010110111",
50815=>"000111101",
50816=>"010100000",
50817=>"001111101",
50818=>"110011000",
50819=>"110111011",
50820=>"000101111",
50821=>"100000010",
50822=>"000101001",
50823=>"000100001",
50824=>"101111100",
50825=>"111000000",
50826=>"111111111",
50827=>"000000110",
50828=>"000010010",
50829=>"100111101",
50830=>"111110010",
50831=>"001100010",
50832=>"111111100",
50833=>"111110101",
50834=>"010000001",
50835=>"011010010",
50836=>"101111010",
50837=>"011000000",
50838=>"000011000",
50839=>"101101100",
50840=>"010110110",
50841=>"010110110",
50842=>"000111001",
50843=>"000010110",
50844=>"111010000",
50845=>"000010010",
50846=>"000000111",
50847=>"111101000",
50848=>"111100100",
50849=>"010000111",
50850=>"000001000",
50851=>"000000000",
50852=>"001100000",
50853=>"110001101",
50854=>"000001000",
50855=>"000010111",
50856=>"010000000",
50857=>"111011110",
50858=>"111111101",
50859=>"001001000",
50860=>"011111011",
50861=>"000000000",
50862=>"011100100",
50863=>"000010010",
50864=>"111010010",
50865=>"101001010",
50866=>"111101100",
50867=>"100001000",
50868=>"101111111",
50869=>"111110101",
50870=>"010000100",
50871=>"010111011",
50872=>"110110100",
50873=>"100110000",
50874=>"000111111",
50875=>"111000111",
50876=>"111111011",
50877=>"110111111",
50878=>"100000100",
50879=>"010000011",
50880=>"000100000",
50881=>"111110010",
50882=>"111010111",
50883=>"101001001",
50884=>"011000000",
50885=>"110100100",
50886=>"010000000",
50887=>"010111011",
50888=>"110111001",
50889=>"010010110",
50890=>"110111101",
50891=>"010000010",
50892=>"000001111",
50893=>"011001000",
50894=>"000001011",
50895=>"000101111",
50896=>"001000001",
50897=>"100111011",
50898=>"110000000",
50899=>"111000101",
50900=>"001001011",
50901=>"101101111",
50902=>"101101101",
50903=>"111001110",
50904=>"000011000",
50905=>"001111101",
50906=>"111101001",
50907=>"010000000",
50908=>"001101110",
50909=>"011111000",
50910=>"110101101",
50911=>"111110110",
50912=>"111010111",
50913=>"101000000",
50914=>"000000111",
50915=>"110011100",
50916=>"000101111",
50917=>"101111111",
50918=>"010000000",
50919=>"100000011",
50920=>"111000100",
50921=>"000000111",
50922=>"100000001",
50923=>"001010100",
50924=>"111000000",
50925=>"000101000",
50926=>"011010000",
50927=>"000101010",
50928=>"000110101",
50929=>"011001001",
50930=>"110000000",
50931=>"001111101",
50932=>"001011110",
50933=>"000001111",
50934=>"000000101",
50935=>"110110011",
50936=>"000000000",
50937=>"111111111",
50938=>"111101101",
50939=>"111001111",
50940=>"101111101",
50941=>"010111011",
50942=>"001000011",
50943=>"111011010",
50944=>"011111010",
50945=>"111110000",
50946=>"101000000",
50947=>"001000010",
50948=>"000100001",
50949=>"111000001",
50950=>"000101111",
50951=>"000110010",
50952=>"001001111",
50953=>"110000000",
50954=>"110110111",
50955=>"110100011",
50956=>"100000100",
50957=>"001001000",
50958=>"100100011",
50959=>"101111100",
50960=>"001000010",
50961=>"011000100",
50962=>"001000000",
50963=>"111010010",
50964=>"000010000",
50965=>"101000001",
50966=>"101000001",
50967=>"100111011",
50968=>"101101110",
50969=>"110110101",
50970=>"111111001",
50971=>"011100101",
50972=>"111101111",
50973=>"101001111",
50974=>"000010010",
50975=>"001101100",
50976=>"110001101",
50977=>"000010000",
50978=>"000000000",
50979=>"000000000",
50980=>"000111111",
50981=>"000110100",
50982=>"010000010",
50983=>"000010011",
50984=>"110111111",
50985=>"110000000",
50986=>"100100000",
50987=>"101101101",
50988=>"100111111",
50989=>"101100000",
50990=>"000000011",
50991=>"011101111",
50992=>"010110000",
50993=>"011101001",
50994=>"000111111",
50995=>"000000111",
50996=>"000100110",
50997=>"111000001",
50998=>"110100001",
50999=>"000000010",
51000=>"010111000",
51001=>"101000000",
51002=>"111101101",
51003=>"011000111",
51004=>"001110110",
51005=>"111111111",
51006=>"000010011",
51007=>"110111001",
51008=>"011000100",
51009=>"101110000",
51010=>"001000000",
51011=>"011001001",
51012=>"111001101",
51013=>"010000000",
51014=>"010111111",
51015=>"111000010",
51016=>"011000000",
51017=>"001111101",
51018=>"000001101",
51019=>"111110111",
51020=>"110101101",
51021=>"101110000",
51022=>"101111111",
51023=>"100101111",
51024=>"001001000",
51025=>"111000000",
51026=>"000010011",
51027=>"001001001",
51028=>"010010000",
51029=>"001111111",
51030=>"001111111",
51031=>"001010010",
51032=>"101111001",
51033=>"101101011",
51034=>"000100100",
51035=>"000011111",
51036=>"000110010",
51037=>"111001001",
51038=>"011111000",
51039=>"100100000",
51040=>"111100000",
51041=>"101011011",
51042=>"111000000",
51043=>"000000101",
51044=>"000111101",
51045=>"101011100",
51046=>"100110111",
51047=>"101001101",
51048=>"101001001",
51049=>"000101111",
51050=>"010010011",
51051=>"111111101",
51052=>"101001001",
51053=>"001011000",
51054=>"000000000",
51055=>"000011011",
51056=>"010110111",
51057=>"111010111",
51058=>"011001110",
51059=>"100000111",
51060=>"101011010",
51061=>"101001000",
51062=>"111111110",
51063=>"100100000",
51064=>"011000000",
51065=>"000010010",
51066=>"000110110",
51067=>"011101101",
51068=>"000111110",
51069=>"011101101",
51070=>"111101111",
51071=>"000001101",
51072=>"010000000",
51073=>"110000000",
51074=>"000000010",
51075=>"000001000",
51076=>"111010010",
51077=>"010101001",
51078=>"110001111",
51079=>"000011011",
51080=>"000000100",
51081=>"000000000",
51082=>"000011010",
51083=>"010000000",
51084=>"100100010",
51085=>"110100000",
51086=>"111001001",
51087=>"000000000",
51088=>"111001101",
51089=>"111011101",
51090=>"110110000",
51091=>"000000000",
51092=>"001110010",
51093=>"111000000",
51094=>"000000000",
51095=>"010100000",
51096=>"010111111",
51097=>"000000000",
51098=>"110111011",
51099=>"000100000",
51100=>"111101111",
51101=>"111011011",
51102=>"111011110",
51103=>"000000101",
51104=>"111000000",
51105=>"111000000",
51106=>"010101101",
51107=>"110000101",
51108=>"010100111",
51109=>"110110010",
51110=>"110000111",
51111=>"010000000",
51112=>"010101001",
51113=>"000110110",
51114=>"010000001",
51115=>"000000000",
51116=>"110111000",
51117=>"000100101",
51118=>"110100011",
51119=>"000100110",
51120=>"100110011",
51121=>"000100110",
51122=>"111100100",
51123=>"001000101",
51124=>"111001001",
51125=>"100000100",
51126=>"001100000",
51127=>"111111001",
51128=>"010111011",
51129=>"000110111",
51130=>"110101101",
51131=>"111101010",
51132=>"110000010",
51133=>"111111011",
51134=>"011001000",
51135=>"000000111",
51136=>"001000001",
51137=>"000000101",
51138=>"111001111",
51139=>"011110111",
51140=>"010010001",
51141=>"100100110",
51142=>"111111111",
51143=>"101111111",
51144=>"010101111",
51145=>"010100101",
51146=>"110001111",
51147=>"101101000",
51148=>"110011010",
51149=>"000111010",
51150=>"100111111",
51151=>"111101111",
51152=>"100101000",
51153=>"101101100",
51154=>"000011000",
51155=>"011111100",
51156=>"000010000",
51157=>"000011011",
51158=>"111000000",
51159=>"111111111",
51160=>"110101111",
51161=>"000010010",
51162=>"100000001",
51163=>"000001101",
51164=>"000100111",
51165=>"000110101",
51166=>"010011001",
51167=>"010110010",
51168=>"000010000",
51169=>"101001001",
51170=>"111101111",
51171=>"000001101",
51172=>"000010000",
51173=>"110101110",
51174=>"001001000",
51175=>"110011000",
51176=>"000010010",
51177=>"000000000",
51178=>"001011111",
51179=>"111100111",
51180=>"100110111",
51181=>"000000010",
51182=>"000000000",
51183=>"000010011",
51184=>"100100010",
51185=>"000001000",
51186=>"000001011",
51187=>"110100101",
51188=>"110010001",
51189=>"000101100",
51190=>"000000110",
51191=>"111101101",
51192=>"010000000",
51193=>"101101011",
51194=>"111101001",
51195=>"000111010",
51196=>"010111111",
51197=>"000010010",
51198=>"011011001",
51199=>"001110010",
51200=>"010010000",
51201=>"111101111",
51202=>"111010101",
51203=>"000000111",
51204=>"011001000",
51205=>"000000000",
51206=>"110100000",
51207=>"000110111",
51208=>"001001111",
51209=>"010010000",
51210=>"011001000",
51211=>"010110110",
51212=>"000000000",
51213=>"000000000",
51214=>"001011011",
51215=>"001000010",
51216=>"000000010",
51217=>"111001000",
51218=>"001001001",
51219=>"101010111",
51220=>"111101111",
51221=>"111000101",
51222=>"101011100",
51223=>"000000000",
51224=>"111000110",
51225=>"010111111",
51226=>"011111111",
51227=>"110010000",
51228=>"111100100",
51229=>"110101011",
51230=>"001000001",
51231=>"001001111",
51232=>"010000000",
51233=>"011101111",
51234=>"100011111",
51235=>"010000000",
51236=>"111100000",
51237=>"000000100",
51238=>"000101111",
51239=>"101101101",
51240=>"101000001",
51241=>"000001000",
51242=>"010011001",
51243=>"110000010",
51244=>"011011001",
51245=>"010000111",
51246=>"000101101",
51247=>"000000100",
51248=>"010101111",
51249=>"101001001",
51250=>"001100111",
51251=>"010111111",
51252=>"111110000",
51253=>"001101111",
51254=>"111000000",
51255=>"000111010",
51256=>"000111110",
51257=>"000000100",
51258=>"100100111",
51259=>"011111110",
51260=>"000100100",
51261=>"111111001",
51262=>"000000010",
51263=>"000000101",
51264=>"111010000",
51265=>"000000000",
51266=>"101010110",
51267=>"001001011",
51268=>"000000110",
51269=>"001101001",
51270=>"011010010",
51271=>"010000000",
51272=>"001101111",
51273=>"000001011",
51274=>"000000010",
51275=>"010000000",
51276=>"000111110",
51277=>"111011001",
51278=>"111000000",
51279=>"001011110",
51280=>"111111000",
51281=>"111010001",
51282=>"011000011",
51283=>"011111110",
51284=>"001001010",
51285=>"000000100",
51286=>"111111100",
51287=>"010010000",
51288=>"000000100",
51289=>"100100011",
51290=>"100101111",
51291=>"110110001",
51292=>"001001101",
51293=>"001001011",
51294=>"011101101",
51295=>"111100100",
51296=>"111000110",
51297=>"000001111",
51298=>"110111110",
51299=>"001111110",
51300=>"100111100",
51301=>"011111111",
51302=>"000000110",
51303=>"111111100",
51304=>"001001111",
51305=>"001101001",
51306=>"110101011",
51307=>"000001001",
51308=>"000101101",
51309=>"111111000",
51310=>"111110100",
51311=>"000000111",
51312=>"011011001",
51313=>"001000110",
51314=>"111000000",
51315=>"000000100",
51316=>"000000010",
51317=>"101101111",
51318=>"110110110",
51319=>"101000010",
51320=>"010100010",
51321=>"110110000",
51322=>"101101101",
51323=>"000001111",
51324=>"110110110",
51325=>"110100000",
51326=>"111010010",
51327=>"000000010",
51328=>"111111011",
51329=>"101000111",
51330=>"000101101",
51331=>"111010111",
51332=>"001101001",
51333=>"100100111",
51334=>"000000001",
51335=>"111000011",
51336=>"101101001",
51337=>"110110110",
51338=>"000101011",
51339=>"111100000",
51340=>"101000001",
51341=>"001001000",
51342=>"110010000",
51343=>"001000001",
51344=>"110100101",
51345=>"000000000",
51346=>"111100101",
51347=>"010000101",
51348=>"111010011",
51349=>"000000000",
51350=>"000111000",
51351=>"100110001",
51352=>"111110100",
51353=>"000001110",
51354=>"111110010",
51355=>"000000110",
51356=>"010010011",
51357=>"011111010",
51358=>"111111110",
51359=>"000001010",
51360=>"010100001",
51361=>"000001111",
51362=>"101001000",
51363=>"000011011",
51364=>"000001111",
51365=>"011011010",
51366=>"101001001",
51367=>"001111110",
51368=>"110011111",
51369=>"000010111",
51370=>"101101111",
51371=>"111001000",
51372=>"001100101",
51373=>"000011111",
51374=>"111111011",
51375=>"110111111",
51376=>"000000110",
51377=>"001111100",
51378=>"111111000",
51379=>"001100110",
51380=>"100110101",
51381=>"000110111",
51382=>"100000100",
51383=>"000100001",
51384=>"000011011",
51385=>"110010110",
51386=>"010000010",
51387=>"011001000",
51388=>"001001000",
51389=>"111111010",
51390=>"000001011",
51391=>"000000100",
51392=>"000001101",
51393=>"110111000",
51394=>"000000111",
51395=>"101011000",
51396=>"010001000",
51397=>"000011001",
51398=>"010100111",
51399=>"010110110",
51400=>"100111110",
51401=>"000000000",
51402=>"000010001",
51403=>"010110110",
51404=>"001000000",
51405=>"011011111",
51406=>"111011000",
51407=>"100101000",
51408=>"000111110",
51409=>"111101000",
51410=>"000110111",
51411=>"101101100",
51412=>"101101100",
51413=>"111100000",
51414=>"000000110",
51415=>"111101001",
51416=>"101001011",
51417=>"011000111",
51418=>"100100100",
51419=>"000100000",
51420=>"110100011",
51421=>"000000000",
51422=>"111110001",
51423=>"001101111",
51424=>"000000000",
51425=>"001111011",
51426=>"001001110",
51427=>"100110110",
51428=>"101000100",
51429=>"110100101",
51430=>"111110000",
51431=>"111100100",
51432=>"001111111",
51433=>"110100110",
51434=>"110010001",
51435=>"111110111",
51436=>"111010000",
51437=>"101101101",
51438=>"110010000",
51439=>"000101111",
51440=>"001010010",
51441=>"010000100",
51442=>"000000101",
51443=>"000000110",
51444=>"000100011",
51445=>"101111010",
51446=>"101000000",
51447=>"100110110",
51448=>"101000101",
51449=>"111111111",
51450=>"111111000",
51451=>"001011111",
51452=>"000001101",
51453=>"010001000",
51454=>"100100100",
51455=>"000111111",
51456=>"000001100",
51457=>"010000000",
51458=>"000000000",
51459=>"000000000",
51460=>"100011111",
51461=>"111010001",
51462=>"011111110",
51463=>"000011011",
51464=>"000110000",
51465=>"101000000",
51466=>"000000000",
51467=>"101100010",
51468=>"010100000",
51469=>"000111110",
51470=>"000001011",
51471=>"000000000",
51472=>"010011111",
51473=>"110000110",
51474=>"111000000",
51475=>"000000101",
51476=>"111110110",
51477=>"010011111",
51478=>"011101001",
51479=>"000010111",
51480=>"100000000",
51481=>"111111111",
51482=>"111111111",
51483=>"101001000",
51484=>"101000010",
51485=>"000101000",
51486=>"001010000",
51487=>"000111111",
51488=>"110000000",
51489=>"001010010",
51490=>"000000010",
51491=>"101111111",
51492=>"100110111",
51493=>"001111111",
51494=>"101000000",
51495=>"011000000",
51496=>"000111000",
51497=>"001000110",
51498=>"000000000",
51499=>"000000010",
51500=>"111110001",
51501=>"111010100",
51502=>"110110100",
51503=>"111111110",
51504=>"100000111",
51505=>"001011100",
51506=>"000111111",
51507=>"111001110",
51508=>"001000000",
51509=>"001000000",
51510=>"110000001",
51511=>"000000000",
51512=>"111010000",
51513=>"000111111",
51514=>"000000100",
51515=>"000011111",
51516=>"011110110",
51517=>"111111111",
51518=>"000000001",
51519=>"000111100",
51520=>"110000000",
51521=>"001111001",
51522=>"111010000",
51523=>"101010000",
51524=>"101000001",
51525=>"000000010",
51526=>"001101011",
51527=>"111111111",
51528=>"110111111",
51529=>"101000001",
51530=>"101000000",
51531=>"101000110",
51532=>"111010000",
51533=>"001111000",
51534=>"000011010",
51535=>"010111101",
51536=>"001101100",
51537=>"110110110",
51538=>"110110111",
51539=>"011001100",
51540=>"000000000",
51541=>"111111001",
51542=>"011111111",
51543=>"110110111",
51544=>"000100000",
51545=>"000000001",
51546=>"100111111",
51547=>"011111111",
51548=>"111011000",
51549=>"001001001",
51550=>"000111010",
51551=>"110110001",
51552=>"000000000",
51553=>"101101100",
51554=>"000000000",
51555=>"001011100",
51556=>"000000100",
51557=>"000100000",
51558=>"000000010",
51559=>"111010000",
51560=>"000010010",
51561=>"000000000",
51562=>"010000000",
51563=>"111101111",
51564=>"100001001",
51565=>"000000000",
51566=>"000000000",
51567=>"000000000",
51568=>"100100101",
51569=>"110000000",
51570=>"001001100",
51571=>"100000101",
51572=>"111001111",
51573=>"011000000",
51574=>"000110110",
51575=>"010111010",
51576=>"000010110",
51577=>"001001111",
51578=>"001000101",
51579=>"000111011",
51580=>"000100000",
51581=>"000100001",
51582=>"000000000",
51583=>"101101100",
51584=>"101111111",
51585=>"111111001",
51586=>"000011000",
51587=>"000000010",
51588=>"110000000",
51589=>"011001001",
51590=>"100111111",
51591=>"100101100",
51592=>"101011011",
51593=>"111010111",
51594=>"110000110",
51595=>"111000001",
51596=>"000111111",
51597=>"101110101",
51598=>"000001001",
51599=>"101001001",
51600=>"101111101",
51601=>"111111111",
51602=>"000000110",
51603=>"111000100",
51604=>"111000101",
51605=>"110010000",
51606=>"111000101",
51607=>"001001000",
51608=>"111111111",
51609=>"000010010",
51610=>"111001101",
51611=>"111010000",
51612=>"111111010",
51613=>"111111111",
51614=>"010000000",
51615=>"111000001",
51616=>"011111111",
51617=>"110010111",
51618=>"011111111",
51619=>"110000000",
51620=>"010000001",
51621=>"110111011",
51622=>"011100001",
51623=>"010001100",
51624=>"111110010",
51625=>"000000000",
51626=>"000000000",
51627=>"011001111",
51628=>"000011000",
51629=>"000010000",
51630=>"010101101",
51631=>"010110010",
51632=>"000111110",
51633=>"000111100",
51634=>"000100000",
51635=>"000000000",
51636=>"001101001",
51637=>"000000000",
51638=>"000010001",
51639=>"000000000",
51640=>"011000011",
51641=>"111000111",
51642=>"010110100",
51643=>"010010111",
51644=>"101101111",
51645=>"111011000",
51646=>"000011000",
51647=>"110111111",
51648=>"010111011",
51649=>"000111101",
51650=>"111001100",
51651=>"001111001",
51652=>"000000000",
51653=>"100010110",
51654=>"111111001",
51655=>"010111110",
51656=>"001000000",
51657=>"011111101",
51658=>"000000000",
51659=>"000111011",
51660=>"000011010",
51661=>"000000000",
51662=>"010100101",
51663=>"000000011",
51664=>"101111110",
51665=>"000001010",
51666=>"000111110",
51667=>"100001001",
51668=>"010111010",
51669=>"000000110",
51670=>"111000000",
51671=>"100000000",
51672=>"010111111",
51673=>"000000101",
51674=>"110111110",
51675=>"111000001",
51676=>"110000011",
51677=>"000111000",
51678=>"110110111",
51679=>"000010111",
51680=>"010111111",
51681=>"111010110",
51682=>"000111000",
51683=>"100100101",
51684=>"000110110",
51685=>"010001000",
51686=>"101001101",
51687=>"000100100",
51688=>"111111001",
51689=>"111100000",
51690=>"001000000",
51691=>"001000001",
51692=>"111111111",
51693=>"110111111",
51694=>"000000000",
51695=>"010110111",
51696=>"101101101",
51697=>"111001100",
51698=>"111010000",
51699=>"000000000",
51700=>"000000000",
51701=>"101101101",
51702=>"101001111",
51703=>"100101111",
51704=>"000111111",
51705=>"011000000",
51706=>"111101111",
51707=>"111000001",
51708=>"000000101",
51709=>"001000010",
51710=>"110110010",
51711=>"010000110",
51712=>"001001100",
51713=>"111000001",
51714=>"111110101",
51715=>"000010110",
51716=>"000100100",
51717=>"100000000",
51718=>"001101000",
51719=>"000000110",
51720=>"000110110",
51721=>"111010010",
51722=>"000000000",
51723=>"111110111",
51724=>"101111101",
51725=>"101011111",
51726=>"100001001",
51727=>"111110000",
51728=>"000000010",
51729=>"110000011",
51730=>"010111011",
51731=>"110000000",
51732=>"000111001",
51733=>"110010000",
51734=>"111011111",
51735=>"111111111",
51736=>"101101111",
51737=>"111101001",
51738=>"011000000",
51739=>"100101111",
51740=>"100000111",
51741=>"000110111",
51742=>"110000011",
51743=>"000010000",
51744=>"101111111",
51745=>"001110101",
51746=>"110010000",
51747=>"010010000",
51748=>"101100100",
51749=>"101101100",
51750=>"110111000",
51751=>"000000000",
51752=>"010111000",
51753=>"101101101",
51754=>"101101100",
51755=>"010000111",
51756=>"101100101",
51757=>"101010000",
51758=>"110100101",
51759=>"111110111",
51760=>"010000010",
51761=>"001001001",
51762=>"000010111",
51763=>"101001010",
51764=>"000000101",
51765=>"010010100",
51766=>"000000100",
51767=>"000000111",
51768=>"010111011",
51769=>"000100000",
51770=>"000000011",
51771=>"101111011",
51772=>"000100011",
51773=>"111111111",
51774=>"111010001",
51775=>"100110000",
51776=>"011111000",
51777=>"010000000",
51778=>"010110111",
51779=>"001001100",
51780=>"010111000",
51781=>"000000110",
51782=>"111111101",
51783=>"110010011",
51784=>"100100000",
51785=>"100110011",
51786=>"111111111",
51787=>"000101001",
51788=>"000000111",
51789=>"001001000",
51790=>"100100100",
51791=>"111011000",
51792=>"010000100",
51793=>"111001111",
51794=>"010011010",
51795=>"011011000",
51796=>"010111101",
51797=>"001011101",
51798=>"001011000",
51799=>"001000111",
51800=>"111111000",
51801=>"001111011",
51802=>"011110100",
51803=>"011101100",
51804=>"110111111",
51805=>"000010001",
51806=>"000010110",
51807=>"100000001",
51808=>"101000000",
51809=>"010000000",
51810=>"111001001",
51811=>"110011111",
51812=>"000101010",
51813=>"111001110",
51814=>"000101000",
51815=>"010100000",
51816=>"111110000",
51817=>"110000001",
51818=>"111000111",
51819=>"000000000",
51820=>"001100101",
51821=>"000000000",
51822=>"111011101",
51823=>"010111111",
51824=>"001101000",
51825=>"110000001",
51826=>"000000101",
51827=>"000000000",
51828=>"111111111",
51829=>"000000100",
51830=>"000000000",
51831=>"000000111",
51832=>"110111111",
51833=>"010110111",
51834=>"101010110",
51835=>"000000000",
51836=>"000110110",
51837=>"100110000",
51838=>"010110111",
51839=>"000101000",
51840=>"101100010",
51841=>"110000100",
51842=>"000111111",
51843=>"000111110",
51844=>"001000000",
51845=>"010010000",
51846=>"011001001",
51847=>"101000001",
51848=>"000101000",
51849=>"100000000",
51850=>"110100010",
51851=>"000011100",
51852=>"000110000",
51853=>"000000010",
51854=>"010111101",
51855=>"101001001",
51856=>"001101100",
51857=>"111100000",
51858=>"011101010",
51859=>"111110111",
51860=>"011111011",
51861=>"000000111",
51862=>"111111101",
51863=>"001111011",
51864=>"010010111",
51865=>"000111111",
51866=>"110010000",
51867=>"010010010",
51868=>"000011000",
51869=>"010111011",
51870=>"010010011",
51871=>"111000000",
51872=>"111011000",
51873=>"111111110",
51874=>"000010010",
51875=>"111010111",
51876=>"110011011",
51877=>"111001011",
51878=>"000101011",
51879=>"000110000",
51880=>"011000001",
51881=>"011111111",
51882=>"000010100",
51883=>"001000000",
51884=>"101111011",
51885=>"000101100",
51886=>"111010110",
51887=>"111010000",
51888=>"111111010",
51889=>"001101000",
51890=>"000000000",
51891=>"001000100",
51892=>"000011000",
51893=>"110011111",
51894=>"111011000",
51895=>"000001000",
51896=>"000001100",
51897=>"100110110",
51898=>"001101010",
51899=>"111110111",
51900=>"110111100",
51901=>"011001111",
51902=>"001011011",
51903=>"011000010",
51904=>"010110100",
51905=>"100001000",
51906=>"010000001",
51907=>"101111111",
51908=>"000000001",
51909=>"110111011",
51910=>"100100011",
51911=>"000001111",
51912=>"000101110",
51913=>"111101101",
51914=>"111011111",
51915=>"010010000",
51916=>"000010011",
51917=>"000001011",
51918=>"000100111",
51919=>"000001111",
51920=>"000110010",
51921=>"011100110",
51922=>"001101111",
51923=>"010010110",
51924=>"000011101",
51925=>"110101001",
51926=>"110111111",
51927=>"110101011",
51928=>"000111000",
51929=>"000000010",
51930=>"111110100",
51931=>"000000000",
51932=>"011110111",
51933=>"010111110",
51934=>"111111000",
51935=>"011000011",
51936=>"010111111",
51937=>"100000111",
51938=>"000011101",
51939=>"100000000",
51940=>"110000010",
51941=>"011001011",
51942=>"111111010",
51943=>"101101111",
51944=>"111100100",
51945=>"011010110",
51946=>"001000000",
51947=>"001011111",
51948=>"111110111",
51949=>"001101101",
51950=>"110010010",
51951=>"000000110",
51952=>"111111100",
51953=>"011101110",
51954=>"000000010",
51955=>"100110000",
51956=>"100111001",
51957=>"100101000",
51958=>"000000011",
51959=>"111010001",
51960=>"000010110",
51961=>"110110101",
51962=>"111111101",
51963=>"000111111",
51964=>"000000110",
51965=>"101001100",
51966=>"101011010",
51967=>"111100111",
51968=>"011001001",
51969=>"000000001",
51970=>"110110100",
51971=>"101111110",
51972=>"001001010",
51973=>"000100110",
51974=>"101111101",
51975=>"100110111",
51976=>"011001011",
51977=>"001000111",
51978=>"000000001",
51979=>"000001000",
51980=>"111001001",
51981=>"000010001",
51982=>"100100100",
51983=>"101011000",
51984=>"101000100",
51985=>"000000011",
51986=>"000000000",
51987=>"000000111",
51988=>"100111111",
51989=>"110110110",
51990=>"011001010",
51991=>"000000000",
51992=>"001000000",
51993=>"110100000",
51994=>"101111111",
51995=>"000000001",
51996=>"000000001",
51997=>"000000000",
51998=>"000000000",
51999=>"111110010",
52000=>"000000000",
52001=>"010110110",
52002=>"000001010",
52003=>"001001001",
52004=>"100100000",
52005=>"000011010",
52006=>"010010010",
52007=>"011000111",
52008=>"011110010",
52009=>"010001101",
52010=>"111110000",
52011=>"110100000",
52012=>"110110110",
52013=>"000110111",
52014=>"010011000",
52015=>"101101010",
52016=>"001000000",
52017=>"001100111",
52018=>"001001101",
52019=>"001001111",
52020=>"000000001",
52021=>"000111110",
52022=>"011000000",
52023=>"011010000",
52024=>"000100111",
52025=>"000100000",
52026=>"000000101",
52027=>"000000001",
52028=>"110011011",
52029=>"110111010",
52030=>"000101001",
52031=>"000110110",
52032=>"111111111",
52033=>"001001111",
52034=>"111111000",
52035=>"011111011",
52036=>"000010111",
52037=>"000000100",
52038=>"100101111",
52039=>"000110110",
52040=>"111111111",
52041=>"001110010",
52042=>"010000001",
52043=>"111010111",
52044=>"000110111",
52045=>"011001110",
52046=>"000000001",
52047=>"011101111",
52048=>"111111110",
52049=>"110111000",
52050=>"111101111",
52051=>"001100000",
52052=>"001101000",
52053=>"011011111",
52054=>"011001001",
52055=>"001001111",
52056=>"110111000",
52057=>"011011110",
52058=>"111011010",
52059=>"100100000",
52060=>"000000000",
52061=>"001001001",
52062=>"010010000",
52063=>"110111101",
52064=>"101101000",
52065=>"010010000",
52066=>"001001101",
52067=>"111111110",
52068=>"000000110",
52069=>"100000110",
52070=>"010111110",
52071=>"111111000",
52072=>"011101111",
52073=>"000001101",
52074=>"111101011",
52075=>"000000000",
52076=>"010000000",
52077=>"101101001",
52078=>"111111100",
52079=>"111000110",
52080=>"001001100",
52081=>"010000000",
52082=>"110000000",
52083=>"001000001",
52084=>"111110010",
52085=>"000000000",
52086=>"010000100",
52087=>"001010000",
52088=>"110110000",
52089=>"000101000",
52090=>"000111110",
52091=>"000001001",
52092=>"101010000",
52093=>"100000000",
52094=>"010100000",
52095=>"001001111",
52096=>"100001001",
52097=>"100100100",
52098=>"111000000",
52099=>"111000000",
52100=>"111001000",
52101=>"111111111",
52102=>"100100110",
52103=>"000000100",
52104=>"100110111",
52105=>"000111101",
52106=>"101100111",
52107=>"000000000",
52108=>"011000000",
52109=>"111101111",
52110=>"000000000",
52111=>"000001000",
52112=>"011001010",
52113=>"111110000",
52114=>"111001111",
52115=>"000000010",
52116=>"000000111",
52117=>"000000111",
52118=>"110111111",
52119=>"110110000",
52120=>"000000000",
52121=>"001111100",
52122=>"000010111",
52123=>"000000011",
52124=>"000000011",
52125=>"000000100",
52126=>"111111111",
52127=>"000100101",
52128=>"110111111",
52129=>"001000101",
52130=>"010001101",
52131=>"111111111",
52132=>"010111000",
52133=>"111111111",
52134=>"111111000",
52135=>"100101000",
52136=>"000000000",
52137=>"000001001",
52138=>"001001001",
52139=>"000000110",
52140=>"001101111",
52141=>"011111111",
52142=>"100101111",
52143=>"111111011",
52144=>"000000000",
52145=>"011101001",
52146=>"001001001",
52147=>"011001000",
52148=>"111111011",
52149=>"111111110",
52150=>"111010000",
52151=>"110110000",
52152=>"111111110",
52153=>"110010000",
52154=>"111010000",
52155=>"110000010",
52156=>"000001001",
52157=>"111111101",
52158=>"101011111",
52159=>"000000111",
52160=>"111110111",
52161=>"001111100",
52162=>"111110110",
52163=>"000000110",
52164=>"000000111",
52165=>"000111011",
52166=>"111000111",
52167=>"111100101",
52168=>"100000000",
52169=>"110110111",
52170=>"000000010",
52171=>"001000011",
52172=>"110110000",
52173=>"011101001",
52174=>"101001000",
52175=>"111001000",
52176=>"111110111",
52177=>"111101111",
52178=>"000000110",
52179=>"101101000",
52180=>"001000000",
52181=>"001001001",
52182=>"000001001",
52183=>"001111111",
52184=>"000000000",
52185=>"111111111",
52186=>"110110111",
52187=>"001000101",
52188=>"110100001",
52189=>"000110010",
52190=>"111110110",
52191=>"010000010",
52192=>"011110000",
52193=>"000011011",
52194=>"000000000",
52195=>"001101110",
52196=>"101101001",
52197=>"000001001",
52198=>"000000000",
52199=>"011101110",
52200=>"111101100",
52201=>"011001000",
52202=>"001101001",
52203=>"001001001",
52204=>"010010000",
52205=>"000000001",
52206=>"110100000",
52207=>"001100110",
52208=>"000000010",
52209=>"010100100",
52210=>"110111000",
52211=>"111111110",
52212=>"110100111",
52213=>"101010010",
52214=>"001000010",
52215=>"111000010",
52216=>"000000111",
52217=>"000110111",
52218=>"111111110",
52219=>"000010110",
52220=>"011111000",
52221=>"111101111",
52222=>"100100110",
52223=>"000001000",
52224=>"110000111",
52225=>"110111110",
52226=>"101001100",
52227=>"000000001",
52228=>"111111111",
52229=>"111001101",
52230=>"000110000",
52231=>"100111111",
52232=>"000000111",
52233=>"100001000",
52234=>"011011010",
52235=>"000000001",
52236=>"001001111",
52237=>"101101001",
52238=>"100000000",
52239=>"111111011",
52240=>"111001001",
52241=>"111001111",
52242=>"111101000",
52243=>"000011001",
52244=>"000110110",
52245=>"011010011",
52246=>"111111010",
52247=>"010110001",
52248=>"111000000",
52249=>"000001111",
52250=>"111111111",
52251=>"000000110",
52252=>"101000010",
52253=>"111111111",
52254=>"111010000",
52255=>"000000000",
52256=>"001001001",
52257=>"100111010",
52258=>"000000000",
52259=>"110001101",
52260=>"100110000",
52261=>"000001111",
52262=>"000000100",
52263=>"010000000",
52264=>"111111111",
52265=>"000001000",
52266=>"101001000",
52267=>"110011110",
52268=>"000010100",
52269=>"111111111",
52270=>"111001011",
52271=>"011000001",
52272=>"111111011",
52273=>"000110100",
52274=>"001111000",
52275=>"110111000",
52276=>"010001111",
52277=>"100100000",
52278=>"001000000",
52279=>"000110010",
52280=>"110000001",
52281=>"000010000",
52282=>"010001111",
52283=>"010110000",
52284=>"000001110",
52285=>"111110100",
52286=>"000001001",
52287=>"000001001",
52288=>"000000111",
52289=>"111100001",
52290=>"000101000",
52291=>"001001000",
52292=>"000010000",
52293=>"000111110",
52294=>"101010000",
52295=>"110110101",
52296=>"101111111",
52297=>"000000000",
52298=>"001100101",
52299=>"000010110",
52300=>"001001111",
52301=>"011011001",
52302=>"000110011",
52303=>"000110000",
52304=>"110000001",
52305=>"111111101",
52306=>"011010000",
52307=>"010010001",
52308=>"000000011",
52309=>"110110000",
52310=>"000100110",
52311=>"111100110",
52312=>"110011001",
52313=>"001111000",
52314=>"000100111",
52315=>"000010110",
52316=>"000000000",
52317=>"000000110",
52318=>"011111000",
52319=>"000000101",
52320=>"111000000",
52321=>"000001111",
52322=>"101001111",
52323=>"111001001",
52324=>"000000000",
52325=>"000010011",
52326=>"000101101",
52327=>"000000110",
52328=>"000000000",
52329=>"001001000",
52330=>"100001001",
52331=>"010000000",
52332=>"001000110",
52333=>"001101111",
52334=>"101111000",
52335=>"110111011",
52336=>"001010011",
52337=>"111110000",
52338=>"100000001",
52339=>"000111000",
52340=>"110101111",
52341=>"100111011",
52342=>"000000000",
52343=>"000000000",
52344=>"101111111",
52345=>"000010010",
52346=>"110101001",
52347=>"001111001",
52348=>"010000001",
52349=>"100101100",
52350=>"010011000",
52351=>"000000111",
52352=>"110011011",
52353=>"111001000",
52354=>"000010010",
52355=>"000110100",
52356=>"011000000",
52357=>"000000000",
52358=>"100000110",
52359=>"000001011",
52360=>"100111110",
52361=>"000000000",
52362=>"101101100",
52363=>"001000001",
52364=>"000001011",
52365=>"101111111",
52366=>"000010000",
52367=>"001001100",
52368=>"000001000",
52369=>"001111110",
52370=>"000001000",
52371=>"110110000",
52372=>"000110110",
52373=>"101001000",
52374=>"111111011",
52375=>"100100000",
52376=>"000101110",
52377=>"111110111",
52378=>"000101010",
52379=>"111001000",
52380=>"000001101",
52381=>"001000010",
52382=>"000000011",
52383=>"010100110",
52384=>"011011110",
52385=>"110010111",
52386=>"000001110",
52387=>"000010111",
52388=>"111000011",
52389=>"100100010",
52390=>"000000010",
52391=>"000011000",
52392=>"111110110",
52393=>"000000000",
52394=>"111001111",
52395=>"110011111",
52396=>"001111111",
52397=>"100000110",
52398=>"101010110",
52399=>"000000111",
52400=>"111111110",
52401=>"000010001",
52402=>"111111111",
52403=>"010001000",
52404=>"101100000",
52405=>"110110000",
52406=>"111101101",
52407=>"000000110",
52408=>"000100110",
52409=>"001111010",
52410=>"000000000",
52411=>"000000011",
52412=>"101000110",
52413=>"111001111",
52414=>"111010010",
52415=>"000001001",
52416=>"110110010",
52417=>"000001110",
52418=>"111110001",
52419=>"100100010",
52420=>"000000111",
52421=>"110110111",
52422=>"000001110",
52423=>"001000111",
52424=>"101111000",
52425=>"101001111",
52426=>"111001011",
52427=>"000100001",
52428=>"000000000",
52429=>"100000001",
52430=>"110100111",
52431=>"010001111",
52432=>"101101001",
52433=>"010111111",
52434=>"000000111",
52435=>"001010111",
52436=>"111101111",
52437=>"100100111",
52438=>"001000000",
52439=>"111110000",
52440=>"000110111",
52441=>"111111101",
52442=>"100110110",
52443=>"101001111",
52444=>"110111001",
52445=>"001001001",
52446=>"010111111",
52447=>"000001111",
52448=>"001001111",
52449=>"111000011",
52450=>"011111111",
52451=>"100110111",
52452=>"000000001",
52453=>"000100010",
52454=>"101111000",
52455=>"000100110",
52456=>"011001111",
52457=>"000110111",
52458=>"101110111",
52459=>"111001001",
52460=>"001001101",
52461=>"000001011",
52462=>"111101110",
52463=>"111110100",
52464=>"000111110",
52465=>"011111110",
52466=>"001011010",
52467=>"000000000",
52468=>"000010010",
52469=>"101001000",
52470=>"001001111",
52471=>"010000111",
52472=>"110000000",
52473=>"000000000",
52474=>"010111111",
52475=>"100110100",
52476=>"111111001",
52477=>"101111111",
52478=>"100111111",
52479=>"000000000",
52480=>"000010110",
52481=>"111111001",
52482=>"000000111",
52483=>"111010000",
52484=>"010000011",
52485=>"101101111",
52486=>"111000000",
52487=>"011110000",
52488=>"000000011",
52489=>"000111000",
52490=>"111101000",
52491=>"111111111",
52492=>"000000111",
52493=>"000000111",
52494=>"100000100",
52495=>"010111111",
52496=>"111101000",
52497=>"000000111",
52498=>"000010111",
52499=>"101100000",
52500=>"000000011",
52501=>"111101100",
52502=>"111110001",
52503=>"010111110",
52504=>"000100110",
52505=>"111111101",
52506=>"010001010",
52507=>"111000000",
52508=>"001100000",
52509=>"101111101",
52510=>"000011000",
52511=>"000000101",
52512=>"110000111",
52513=>"111000000",
52514=>"000000111",
52515=>"000010000",
52516=>"011010110",
52517=>"000000000",
52518=>"111100010",
52519=>"010010111",
52520=>"011011100",
52521=>"010000001",
52522=>"111011000",
52523=>"111111010",
52524=>"011000000",
52525=>"111110010",
52526=>"111111101",
52527=>"000000100",
52528=>"111011111",
52529=>"110110011",
52530=>"010111111",
52531=>"111001110",
52532=>"101000000",
52533=>"000000000",
52534=>"101100000",
52535=>"100100000",
52536=>"110000000",
52537=>"000101101",
52538=>"000000111",
52539=>"001010010",
52540=>"011001100",
52541=>"011000000",
52542=>"001001111",
52543=>"101000000",
52544=>"010111111",
52545=>"000111000",
52546=>"110010101",
52547=>"000000000",
52548=>"111111000",
52549=>"001101001",
52550=>"110110000",
52551=>"001000111",
52552=>"110111110",
52553=>"111110010",
52554=>"001101000",
52555=>"111100000",
52556=>"000000111",
52557=>"110000111",
52558=>"110001100",
52559=>"110000100",
52560=>"000101101",
52561=>"111000000",
52562=>"010101111",
52563=>"001010010",
52564=>"000000000",
52565=>"111100001",
52566=>"110010000",
52567=>"111000000",
52568=>"011001111",
52569=>"011010111",
52570=>"100100111",
52571=>"111110111",
52572=>"111000000",
52573=>"001110110",
52574=>"000111111",
52575=>"001010000",
52576=>"110010111",
52577=>"111111000",
52578=>"000111111",
52579=>"011011001",
52580=>"110001011",
52581=>"000000100",
52582=>"000010101",
52583=>"100001001",
52584=>"110000010",
52585=>"000000011",
52586=>"000111111",
52587=>"000101111",
52588=>"111000000",
52589=>"000000111",
52590=>"111000000",
52591=>"010000000",
52592=>"111110110",
52593=>"111010000",
52594=>"000010000",
52595=>"001000111",
52596=>"100000000",
52597=>"000111101",
52598=>"111010011",
52599=>"000001000",
52600=>"101010010",
52601=>"011111111",
52602=>"001110000",
52603=>"000011111",
52604=>"010001000",
52605=>"000010011",
52606=>"100000000",
52607=>"000101100",
52608=>"111000000",
52609=>"101001010",
52610=>"111110000",
52611=>"111111100",
52612=>"000101101",
52613=>"000111001",
52614=>"010000000",
52615=>"111010000",
52616=>"011010000",
52617=>"000111001",
52618=>"011011110",
52619=>"000011111",
52620=>"100101001",
52621=>"111000100",
52622=>"100000000",
52623=>"001001001",
52624=>"000011110",
52625=>"000000000",
52626=>"000000000",
52627=>"101001011",
52628=>"111100000",
52629=>"101011011",
52630=>"110100101",
52631=>"111110110",
52632=>"010111100",
52633=>"111001000",
52634=>"100000111",
52635=>"100000000",
52636=>"011000000",
52637=>"100000000",
52638=>"111010000",
52639=>"110000110",
52640=>"001010110",
52641=>"010011111",
52642=>"111010111",
52643=>"111111000",
52644=>"000011111",
52645=>"110011000",
52646=>"001011111",
52647=>"101000000",
52648=>"111101000",
52649=>"111000000",
52650=>"100010110",
52651=>"000000000",
52652=>"000000111",
52653=>"111110010",
52654=>"000000011",
52655=>"111111000",
52656=>"101111011",
52657=>"110110111",
52658=>"100110000",
52659=>"110000010",
52660=>"110110111",
52661=>"111010011",
52662=>"101011101",
52663=>"010111111",
52664=>"110000100",
52665=>"111011000",
52666=>"011100000",
52667=>"011010000",
52668=>"000101111",
52669=>"000100111",
52670=>"110000000",
52671=>"000000000",
52672=>"011011000",
52673=>"010000000",
52674=>"000000000",
52675=>"000000000",
52676=>"001101111",
52677=>"100100100",
52678=>"111011011",
52679=>"000111111",
52680=>"101110111",
52681=>"001101111",
52682=>"111100000",
52683=>"100100111",
52684=>"101010100",
52685=>"111100000",
52686=>"010001100",
52687=>"000000111",
52688=>"001100111",
52689=>"001000000",
52690=>"111111001",
52691=>"011010110",
52692=>"100110000",
52693=>"111001001",
52694=>"111000110",
52695=>"111000000",
52696=>"111111011",
52697=>"100000000",
52698=>"110010110",
52699=>"000101111",
52700=>"111111000",
52701=>"000000111",
52702=>"111001101",
52703=>"111111000",
52704=>"000000010",
52705=>"001011001",
52706=>"000111111",
52707=>"000100011",
52708=>"101000000",
52709=>"100001100",
52710=>"110000010",
52711=>"110100100",
52712=>"010011010",
52713=>"101101111",
52714=>"000000000",
52715=>"000011011",
52716=>"000001011",
52717=>"000100100",
52718=>"101000000",
52719=>"111000000",
52720=>"000000100",
52721=>"001000011",
52722=>"110010101",
52723=>"010011110",
52724=>"011011011",
52725=>"100111101",
52726=>"000000111",
52727=>"111111111",
52728=>"010010000",
52729=>"010000111",
52730=>"011001100",
52731=>"111110110",
52732=>"111100000",
52733=>"111111011",
52734=>"000000110",
52735=>"110110000",
52736=>"100111011",
52737=>"110011101",
52738=>"001000111",
52739=>"010010001",
52740=>"100010000",
52741=>"000000101",
52742=>"001110000",
52743=>"000101101",
52744=>"100001111",
52745=>"111100111",
52746=>"000000001",
52747=>"101101101",
52748=>"110110010",
52749=>"000100110",
52750=>"010110000",
52751=>"000000111",
52752=>"001110101",
52753=>"100000000",
52754=>"111111010",
52755=>"011111001",
52756=>"111111111",
52757=>"011001101",
52758=>"010111011",
52759=>"000000001",
52760=>"000100111",
52761=>"111100110",
52762=>"000000111",
52763=>"000000010",
52764=>"100111001",
52765=>"101101010",
52766=>"110111101",
52767=>"100000000",
52768=>"100000111",
52769=>"000000011",
52770=>"111011000",
52771=>"101000100",
52772=>"110110100",
52773=>"011000000",
52774=>"100000010",
52775=>"000000000",
52776=>"000111011",
52777=>"101000000",
52778=>"111100111",
52779=>"101111100",
52780=>"111011110",
52781=>"011111011",
52782=>"100111101",
52783=>"000000101",
52784=>"000000000",
52785=>"110110111",
52786=>"011101110",
52787=>"111100000",
52788=>"000000000",
52789=>"111010000",
52790=>"000000010",
52791=>"000110010",
52792=>"000111111",
52793=>"000110000",
52794=>"110101101",
52795=>"000000000",
52796=>"000110000",
52797=>"111010101",
52798=>"100000010",
52799=>"000011111",
52800=>"111111000",
52801=>"000110000",
52802=>"101101101",
52803=>"000110111",
52804=>"111111011",
52805=>"001010101",
52806=>"000011111",
52807=>"111111011",
52808=>"011111111",
52809=>"111111000",
52810=>"000100101",
52811=>"110111101",
52812=>"011100111",
52813=>"111111010",
52814=>"100010001",
52815=>"111111111",
52816=>"100010010",
52817=>"111111110",
52818=>"111111100",
52819=>"111011001",
52820=>"111111010",
52821=>"010011001",
52822=>"100111111",
52823=>"111101111",
52824=>"001000110",
52825=>"010010000",
52826=>"011000000",
52827=>"100110011",
52828=>"000010000",
52829=>"010011000",
52830=>"010111110",
52831=>"011011010",
52832=>"010000001",
52833=>"010110000",
52834=>"011100111",
52835=>"011011000",
52836=>"101110000",
52837=>"011001001",
52838=>"000110111",
52839=>"100101111",
52840=>"111000010",
52841=>"001100000",
52842=>"100111111",
52843=>"101011000",
52844=>"100111101",
52845=>"111000111",
52846=>"000000000",
52847=>"000000111",
52848=>"011011011",
52849=>"000000101",
52850=>"000000000",
52851=>"111101111",
52852=>"100100110",
52853=>"000000101",
52854=>"000000000",
52855=>"010000111",
52856=>"110000111",
52857=>"110000111",
52858=>"111011101",
52859=>"000000000",
52860=>"110011001",
52861=>"111110100",
52862=>"000000111",
52863=>"110000000",
52864=>"000101111",
52865=>"011111100",
52866=>"000010111",
52867=>"001100000",
52868=>"111011010",
52869=>"001001111",
52870=>"100100101",
52871=>"100100100",
52872=>"111111000",
52873=>"000000001",
52874=>"000000010",
52875=>"010101111",
52876=>"001000010",
52877=>"000101011",
52878=>"000011000",
52879=>"001001111",
52880=>"111011111",
52881=>"000000000",
52882=>"000000000",
52883=>"100110000",
52884=>"000011100",
52885=>"000101110",
52886=>"111111100",
52887=>"001110100",
52888=>"100000011",
52889=>"011000001",
52890=>"001100111",
52891=>"111100101",
52892=>"011011111",
52893=>"000100000",
52894=>"111010010",
52895=>"111110110",
52896=>"001010011",
52897=>"011011111",
52898=>"000000101",
52899=>"111111111",
52900=>"111110000",
52901=>"001000010",
52902=>"011011000",
52903=>"110111001",
52904=>"000111101",
52905=>"010011000",
52906=>"101101111",
52907=>"110111011",
52908=>"111101100",
52909=>"010110011",
52910=>"011111000",
52911=>"111000001",
52912=>"110100101",
52913=>"100111000",
52914=>"111011000",
52915=>"110001001",
52916=>"000110000",
52917=>"111111111",
52918=>"111110000",
52919=>"110000111",
52920=>"010011010",
52921=>"100011001",
52922=>"000010011",
52923=>"101111010",
52924=>"000011010",
52925=>"111101111",
52926=>"111111111",
52927=>"100000000",
52928=>"010111010",
52929=>"110011001",
52930=>"111111000",
52931=>"100110011",
52932=>"111001111",
52933=>"111111111",
52934=>"000100111",
52935=>"011000100",
52936=>"100000100",
52937=>"010100010",
52938=>"101000111",
52939=>"000000111",
52940=>"000000000",
52941=>"011110110",
52942=>"010000011",
52943=>"111111110",
52944=>"010111111",
52945=>"110110111",
52946=>"100011101",
52947=>"000010010",
52948=>"000111011",
52949=>"100000000",
52950=>"010111010",
52951=>"011110000",
52952=>"001000000",
52953=>"000011001",
52954=>"111110100",
52955=>"111100101",
52956=>"110110110",
52957=>"010100111",
52958=>"110000010",
52959=>"000010111",
52960=>"000100111",
52961=>"111010010",
52962=>"010000001",
52963=>"111011001",
52964=>"000000000",
52965=>"101100111",
52966=>"000000101",
52967=>"100110010",
52968=>"101100111",
52969=>"101100011",
52970=>"001000000",
52971=>"000000101",
52972=>"000000111",
52973=>"111000000",
52974=>"110111111",
52975=>"000101111",
52976=>"101001111",
52977=>"111111011",
52978=>"010111001",
52979=>"010001000",
52980=>"001011110",
52981=>"100100001",
52982=>"111100001",
52983=>"110100001",
52984=>"010011000",
52985=>"000000111",
52986=>"100011110",
52987=>"100110010",
52988=>"011011111",
52989=>"101000111",
52990=>"110110010",
52991=>"000111100",
52992=>"011001010",
52993=>"000000010",
52994=>"000010000",
52995=>"111000110",
52996=>"000000111",
52997=>"110101100",
52998=>"000000100",
52999=>"111101110",
53000=>"011011000",
53001=>"000000101",
53002=>"000111110",
53003=>"000011010",
53004=>"000111010",
53005=>"111111100",
53006=>"000011011",
53007=>"001101100",
53008=>"111101111",
53009=>"000111111",
53010=>"111000000",
53011=>"000000111",
53012=>"110010100",
53013=>"010010000",
53014=>"011001100",
53015=>"011010010",
53016=>"000000011",
53017=>"000101110",
53018=>"010000000",
53019=>"000111111",
53020=>"111001111",
53021=>"110100111",
53022=>"111101000",
53023=>"100101001",
53024=>"000101111",
53025=>"000111000",
53026=>"000010110",
53027=>"001001011",
53028=>"111101100",
53029=>"001001011",
53030=>"111000001",
53031=>"000000100",
53032=>"110110000",
53033=>"100000001",
53034=>"101000100",
53035=>"000000000",
53036=>"100001011",
53037=>"111010000",
53038=>"111111001",
53039=>"111111001",
53040=>"000000000",
53041=>"001001011",
53042=>"101001101",
53043=>"111000000",
53044=>"000111111",
53045=>"000010001",
53046=>"111111111",
53047=>"111001001",
53048=>"111101011",
53049=>"110110000",
53050=>"000101000",
53051=>"000111100",
53052=>"101011011",
53053=>"111111111",
53054=>"110000000",
53055=>"110011111",
53056=>"010110111",
53057=>"000000111",
53058=>"001001000",
53059=>"011011001",
53060=>"111000011",
53061=>"110010000",
53062=>"000111110",
53063=>"111111000",
53064=>"110111100",
53065=>"111111111",
53066=>"111001101",
53067=>"100111111",
53068=>"001000011",
53069=>"000011011",
53070=>"111111100",
53071=>"000010111",
53072=>"100100111",
53073=>"111000000",
53074=>"111111000",
53075=>"111000111",
53076=>"111111111",
53077=>"111010111",
53078=>"000001001",
53079=>"111111111",
53080=>"000010110",
53081=>"111001001",
53082=>"000100011",
53083=>"000111011",
53084=>"110110111",
53085=>"001001001",
53086=>"000010111",
53087=>"111100100",
53088=>"001010011",
53089=>"010100111",
53090=>"010011110",
53091=>"101001111",
53092=>"110101110",
53093=>"000001001",
53094=>"000111110",
53095=>"111000000",
53096=>"000110111",
53097=>"000000000",
53098=>"111011000",
53099=>"111000010",
53100=>"111000000",
53101=>"000001110",
53102=>"111111110",
53103=>"000000110",
53104=>"100100000",
53105=>"000001001",
53106=>"011111110",
53107=>"000000011",
53108=>"111000000",
53109=>"101000000",
53110=>"000000100",
53111=>"100110110",
53112=>"111010110",
53113=>"010000110",
53114=>"000000000",
53115=>"010111111",
53116=>"011001101",
53117=>"110100000",
53118=>"110111101",
53119=>"110111101",
53120=>"110110001",
53121=>"111101100",
53122=>"001111001",
53123=>"000000010",
53124=>"111111000",
53125=>"001111010",
53126=>"000000111",
53127=>"100100100",
53128=>"111011011",
53129=>"100111111",
53130=>"110111111",
53131=>"010000010",
53132=>"000111111",
53133=>"000111111",
53134=>"110101111",
53135=>"000001001",
53136=>"101100100",
53137=>"000000110",
53138=>"111111101",
53139=>"111000000",
53140=>"111101001",
53141=>"111101101",
53142=>"000010010",
53143=>"110100000",
53144=>"000000010",
53145=>"011000010",
53146=>"000010111",
53147=>"111111111",
53148=>"000001111",
53149=>"000000111",
53150=>"000000111",
53151=>"111000000",
53152=>"000111100",
53153=>"111111000",
53154=>"111101100",
53155=>"000000111",
53156=>"111000000",
53157=>"000010000",
53158=>"111111001",
53159=>"000000111",
53160=>"111111111",
53161=>"100100000",
53162=>"111011000",
53163=>"000000010",
53164=>"101111100",
53165=>"111001000",
53166=>"100101011",
53167=>"110110110",
53168=>"001000010",
53169=>"011011001",
53170=>"101001101",
53171=>"000001100",
53172=>"010110110",
53173=>"111111101",
53174=>"000111111",
53175=>"000000100",
53176=>"100100100",
53177=>"111001101",
53178=>"000000010",
53179=>"001001111",
53180=>"000110110",
53181=>"110000011",
53182=>"111111110",
53183=>"111101101",
53184=>"010110111",
53185=>"000110111",
53186=>"101111111",
53187=>"111111000",
53188=>"100111000",
53189=>"110110010",
53190=>"111110000",
53191=>"011011000",
53192=>"000011010",
53193=>"100110000",
53194=>"111101100",
53195=>"000111111",
53196=>"000000111",
53197=>"110100001",
53198=>"000010000",
53199=>"010001000",
53200=>"000010010",
53201=>"001011011",
53202=>"010111000",
53203=>"101100000",
53204=>"110111110",
53205=>"000000100",
53206=>"111111110",
53207=>"111111010",
53208=>"000000110",
53209=>"110010011",
53210=>"001100100",
53211=>"000000010",
53212=>"111111011",
53213=>"011110111",
53214=>"010111111",
53215=>"111110010",
53216=>"001110111",
53217=>"000000000",
53218=>"010011010",
53219=>"100100111",
53220=>"010111111",
53221=>"000111000",
53222=>"110000000",
53223=>"110101101",
53224=>"010010000",
53225=>"101000110",
53226=>"010110111",
53227=>"001111111",
53228=>"000000101",
53229=>"101001000",
53230=>"011010000",
53231=>"011000000",
53232=>"111111010",
53233=>"011011010",
53234=>"111001001",
53235=>"110101101",
53236=>"110110101",
53237=>"000000000",
53238=>"000000111",
53239=>"000000111",
53240=>"010010000",
53241=>"111101000",
53242=>"111111111",
53243=>"111111010",
53244=>"111111111",
53245=>"010110111",
53246=>"110100111",
53247=>"101001000",
53248=>"110100100",
53249=>"000111111",
53250=>"011000111",
53251=>"000111111",
53252=>"000111000",
53253=>"000000011",
53254=>"111111100",
53255=>"011011111",
53256=>"000100001",
53257=>"010000111",
53258=>"111000100",
53259=>"000000000",
53260=>"101111010",
53261=>"000000011",
53262=>"001011100",
53263=>"101000001",
53264=>"000100000",
53265=>"111000000",
53266=>"110000010",
53267=>"111100001",
53268=>"000001111",
53269=>"111111000",
53270=>"000111001",
53271=>"000111110",
53272=>"000000101",
53273=>"000111111",
53274=>"100100000",
53275=>"110000111",
53276=>"000100000",
53277=>"001000000",
53278=>"101001011",
53279=>"111000000",
53280=>"000000000",
53281=>"000100110",
53282=>"111000100",
53283=>"100111000",
53284=>"010010000",
53285=>"011011011",
53286=>"100110000",
53287=>"101000000",
53288=>"110111111",
53289=>"000010000",
53290=>"000000000",
53291=>"111000000",
53292=>"111111011",
53293=>"111111000",
53294=>"101100111",
53295=>"000000011",
53296=>"100001000",
53297=>"110011010",
53298=>"000000101",
53299=>"000000111",
53300=>"111000101",
53301=>"111001000",
53302=>"011011111",
53303=>"010011000",
53304=>"101010111",
53305=>"000000111",
53306=>"000101010",
53307=>"000101111",
53308=>"011011011",
53309=>"010011011",
53310=>"010000101",
53311=>"011011001",
53312=>"101000111",
53313=>"001001011",
53314=>"101001111",
53315=>"011100010",
53316=>"001000010",
53317=>"101101101",
53318=>"111111000",
53319=>"000000011",
53320=>"010111111",
53321=>"101000110",
53322=>"000000000",
53323=>"111000000",
53324=>"101000111",
53325=>"011111111",
53326=>"000110111",
53327=>"111000000",
53328=>"000001000",
53329=>"011111111",
53330=>"101111001",
53331=>"001100000",
53332=>"000000000",
53333=>"100110100",
53334=>"111010000",
53335=>"000000100",
53336=>"000111111",
53337=>"000011110",
53338=>"011000000",
53339=>"000100011",
53340=>"001000101",
53341=>"000100110",
53342=>"111111000",
53343=>"000001011",
53344=>"000001111",
53345=>"111101100",
53346=>"001000111",
53347=>"100101110",
53348=>"100000011",
53349=>"000000100",
53350=>"001001110",
53351=>"110110001",
53352=>"001110111",
53353=>"111011111",
53354=>"110011000",
53355=>"000101001",
53356=>"001000111",
53357=>"111110010",
53358=>"001001001",
53359=>"010111111",
53360=>"001011010",
53361=>"000110110",
53362=>"100100100",
53363=>"010111001",
53364=>"000011000",
53365=>"100100101",
53366=>"101010111",
53367=>"111001001",
53368=>"010000111",
53369=>"111011010",
53370=>"110111101",
53371=>"100111110",
53372=>"111011001",
53373=>"100011010",
53374=>"111011101",
53375=>"110010001",
53376=>"001001000",
53377=>"000110101",
53378=>"000000111",
53379=>"011110000",
53380=>"111111000",
53381=>"110000000",
53382=>"100101111",
53383=>"000011001",
53384=>"010110000",
53385=>"000001000",
53386=>"111111000",
53387=>"001000111",
53388=>"010110101",
53389=>"001000001",
53390=>"000000000",
53391=>"101000000",
53392=>"000111011",
53393=>"111110000",
53394=>"010000111",
53395=>"000010111",
53396=>"100111000",
53397=>"001000111",
53398=>"101101111",
53399=>"001110110",
53400=>"110010000",
53401=>"000000110",
53402=>"000111000",
53403=>"111000011",
53404=>"111110011",
53405=>"001000111",
53406=>"001111000",
53407=>"111001111",
53408=>"011111011",
53409=>"111010111",
53410=>"111111110",
53411=>"000000000",
53412=>"111110001",
53413=>"110011001",
53414=>"111111111",
53415=>"001111111",
53416=>"011111000",
53417=>"000100001",
53418=>"000000000",
53419=>"000000100",
53420=>"011000011",
53421=>"000000000",
53422=>"110100100",
53423=>"111111000",
53424=>"101000000",
53425=>"000100100",
53426=>"101001111",
53427=>"100111011",
53428=>"111010010",
53429=>"101100111",
53430=>"111010100",
53431=>"001101001",
53432=>"110110100",
53433=>"111111100",
53434=>"100101000",
53435=>"100000000",
53436=>"111000000",
53437=>"000011001",
53438=>"001010100",
53439=>"000101000",
53440=>"101000000",
53441=>"010000000",
53442=>"000000000",
53443=>"111110100",
53444=>"110000000",
53445=>"010000001",
53446=>"111110000",
53447=>"110111000",
53448=>"110000111",
53449=>"110000001",
53450=>"000000100",
53451=>"111001111",
53452=>"001001010",
53453=>"000111101",
53454=>"111000101",
53455=>"110000000",
53456=>"011011000",
53457=>"111011000",
53458=>"111010111",
53459=>"111000000",
53460=>"000000000",
53461=>"000000001",
53462=>"001000000",
53463=>"000001000",
53464=>"111111000",
53465=>"111011100",
53466=>"100001111",
53467=>"011000000",
53468=>"001011111",
53469=>"111111111",
53470=>"101101101",
53471=>"001101010",
53472=>"010000001",
53473=>"001000111",
53474=>"111110000",
53475=>"100100000",
53476=>"101001000",
53477=>"011000000",
53478=>"001011111",
53479=>"111111011",
53480=>"000000110",
53481=>"001000111",
53482=>"011001001",
53483=>"101000001",
53484=>"000000000",
53485=>"000111101",
53486=>"000100000",
53487=>"000010000",
53488=>"111000000",
53489=>"100000110",
53490=>"111101001",
53491=>"100001010",
53492=>"100001011",
53493=>"010000000",
53494=>"000101000",
53495=>"111111100",
53496=>"000111111",
53497=>"111011100",
53498=>"000011000",
53499=>"001000001",
53500=>"110001000",
53501=>"001000000",
53502=>"110000000",
53503=>"000000110",
53504=>"010000000",
53505=>"000000001",
53506=>"000000101",
53507=>"001000000",
53508=>"101001111",
53509=>"000100010",
53510=>"101000011",
53511=>"100001111",
53512=>"101100111",
53513=>"101001001",
53514=>"001001011",
53515=>"010010111",
53516=>"000000010",
53517=>"010000000",
53518=>"001111110",
53519=>"111011010",
53520=>"010110111",
53521=>"000111101",
53522=>"101001010",
53523=>"000011011",
53524=>"111111010",
53525=>"000000010",
53526=>"010110110",
53527=>"001111111",
53528=>"101000000",
53529=>"101100111",
53530=>"001011111",
53531=>"000010110",
53532=>"010100000",
53533=>"000000000",
53534=>"001000000",
53535=>"111111000",
53536=>"010000101",
53537=>"000000111",
53538=>"101100100",
53539=>"101011010",
53540=>"010110011",
53541=>"000000001",
53542=>"001000000",
53543=>"100101100",
53544=>"110110110",
53545=>"110111111",
53546=>"010000000",
53547=>"010000000",
53548=>"001011011",
53549=>"000000000",
53550=>"000100001",
53551=>"110110111",
53552=>"001000000",
53553=>"100110111",
53554=>"000111111",
53555=>"111010111",
53556=>"000000000",
53557=>"111111111",
53558=>"011000000",
53559=>"100000000",
53560=>"000010111",
53561=>"001011001",
53562=>"111101000",
53563=>"000101111",
53564=>"000111111",
53565=>"111110110",
53566=>"000000001",
53567=>"110110110",
53568=>"001001101",
53569=>"101011001",
53570=>"111110000",
53571=>"110111100",
53572=>"111101010",
53573=>"101101010",
53574=>"011101111",
53575=>"001011010",
53576=>"001111111",
53577=>"001000000",
53578=>"101000000",
53579=>"111111111",
53580=>"000000000",
53581=>"001001111",
53582=>"011010111",
53583=>"111011111",
53584=>"110000000",
53585=>"100111110",
53586=>"001000000",
53587=>"001001000",
53588=>"000000000",
53589=>"000111011",
53590=>"011011011",
53591=>"000000001",
53592=>"010110000",
53593=>"110011000",
53594=>"111111000",
53595=>"110100010",
53596=>"000000111",
53597=>"011001100",
53598=>"101110100",
53599=>"011000001",
53600=>"111111000",
53601=>"010011011",
53602=>"100000100",
53603=>"110110000",
53604=>"000111111",
53605=>"111100010",
53606=>"110111110",
53607=>"111100000",
53608=>"011111000",
53609=>"000111010",
53610=>"000010111",
53611=>"010011111",
53612=>"101001111",
53613=>"000010111",
53614=>"101000101",
53615=>"000001111",
53616=>"011011011",
53617=>"000010111",
53618=>"110000000",
53619=>"001000000",
53620=>"111111111",
53621=>"100001000",
53622=>"011111010",
53623=>"101111111",
53624=>"001111100",
53625=>"010111111",
53626=>"110010000",
53627=>"000001111",
53628=>"101100111",
53629=>"101101001",
53630=>"111101101",
53631=>"111100101",
53632=>"001001001",
53633=>"100000010",
53634=>"110000111",
53635=>"111111111",
53636=>"100100000",
53637=>"001000000",
53638=>"001100100",
53639=>"100011110",
53640=>"111111110",
53641=>"000000001",
53642=>"111111000",
53643=>"000000001",
53644=>"001101000",
53645=>"111100111",
53646=>"000101100",
53647=>"101001001",
53648=>"100111000",
53649=>"110111110",
53650=>"000001101",
53651=>"111010111",
53652=>"001111111",
53653=>"000101111",
53654=>"111010110",
53655=>"101100101",
53656=>"110111000",
53657=>"100100000",
53658=>"010110010",
53659=>"100011111",
53660=>"011000000",
53661=>"010000001",
53662=>"001000101",
53663=>"000000110",
53664=>"000111110",
53665=>"111111101",
53666=>"101001000",
53667=>"010111010",
53668=>"000101010",
53669=>"111001010",
53670=>"000001101",
53671=>"001111111",
53672=>"000000000",
53673=>"001011011",
53674=>"000000000",
53675=>"010001101",
53676=>"001010111",
53677=>"000000000",
53678=>"011011001",
53679=>"111010000",
53680=>"000010111",
53681=>"001110111",
53682=>"101101111",
53683=>"110110111",
53684=>"111110010",
53685=>"111101111",
53686=>"000000000",
53687=>"010110001",
53688=>"000011011",
53689=>"001011011",
53690=>"000010000",
53691=>"111111011",
53692=>"001111000",
53693=>"000110111",
53694=>"011011011",
53695=>"001000000",
53696=>"000000101",
53697=>"010110000",
53698=>"010011000",
53699=>"110010000",
53700=>"000001101",
53701=>"000000001",
53702=>"011000100",
53703=>"101000000",
53704=>"000000010",
53705=>"000100000",
53706=>"001000001",
53707=>"000000001",
53708=>"111101000",
53709=>"101011110",
53710=>"111011001",
53711=>"111111100",
53712=>"110010000",
53713=>"111100110",
53714=>"101111111",
53715=>"011110000",
53716=>"000000011",
53717=>"000111001",
53718=>"011111000",
53719=>"000001111",
53720=>"000000011",
53721=>"101011011",
53722=>"100111110",
53723=>"110000000",
53724=>"111101111",
53725=>"111010111",
53726=>"111101010",
53727=>"000000000",
53728=>"101101011",
53729=>"100000010",
53730=>"110101000",
53731=>"110111111",
53732=>"000000001",
53733=>"000000011",
53734=>"111010111",
53735=>"111111001",
53736=>"111000000",
53737=>"011111111",
53738=>"110110100",
53739=>"111111110",
53740=>"000011011",
53741=>"000000000",
53742=>"001111010",
53743=>"000101000",
53744=>"000010010",
53745=>"001000000",
53746=>"000000000",
53747=>"111011000",
53748=>"000110010",
53749=>"111000000",
53750=>"111011000",
53751=>"111111100",
53752=>"000000111",
53753=>"011000111",
53754=>"111111110",
53755=>"000111110",
53756=>"110111110",
53757=>"111111111",
53758=>"101011011",
53759=>"010010000",
53760=>"011001110",
53761=>"010010010",
53762=>"000000111",
53763=>"101101000",
53764=>"111011001",
53765=>"000001011",
53766=>"111110000",
53767=>"111111101",
53768=>"001101110",
53769=>"000010111",
53770=>"111100001",
53771=>"100101101",
53772=>"101101000",
53773=>"010111000",
53774=>"011111100",
53775=>"111111011",
53776=>"111111011",
53777=>"111111000",
53778=>"000111111",
53779=>"000010000",
53780=>"000111010",
53781=>"011111100",
53782=>"111111011",
53783=>"000111001",
53784=>"001110111",
53785=>"011001001",
53786=>"001111011",
53787=>"000000000",
53788=>"110000000",
53789=>"000000000",
53790=>"000110011",
53791=>"110110000",
53792=>"010000000",
53793=>"101101010",
53794=>"101010111",
53795=>"000000111",
53796=>"111111011",
53797=>"000001000",
53798=>"000101101",
53799=>"111011111",
53800=>"100001000",
53801=>"000000111",
53802=>"000100000",
53803=>"101010001",
53804=>"000111000",
53805=>"111000000",
53806=>"100010101",
53807=>"111110000",
53808=>"111101000",
53809=>"111001011",
53810=>"011010111",
53811=>"010011000",
53812=>"000000000",
53813=>"001000000",
53814=>"010010000",
53815=>"111000000",
53816=>"001100111",
53817=>"110100000",
53818=>"101101010",
53819=>"100101101",
53820=>"010000000",
53821=>"011010111",
53822=>"101001000",
53823=>"101110000",
53824=>"000000111",
53825=>"010000110",
53826=>"000010000",
53827=>"011011100",
53828=>"001101111",
53829=>"001000000",
53830=>"100110000",
53831=>"111111111",
53832=>"101100011",
53833=>"001000000",
53834=>"111111000",
53835=>"010111001",
53836=>"001001011",
53837=>"001011010",
53838=>"000100100",
53839=>"100000101",
53840=>"000000000",
53841=>"000111111",
53842=>"101001111",
53843=>"111100010",
53844=>"000010001",
53845=>"000100011",
53846=>"011111000",
53847=>"000001011",
53848=>"000000101",
53849=>"111111110",
53850=>"111000000",
53851=>"111111010",
53852=>"000111111",
53853=>"001100000",
53854=>"010010111",
53855=>"110011000",
53856=>"000011110",
53857=>"010000010",
53858=>"000000111",
53859=>"111001000",
53860=>"111101000",
53861=>"011111000",
53862=>"010001000",
53863=>"000000010",
53864=>"111111010",
53865=>"000000111",
53866=>"011010111",
53867=>"010000001",
53868=>"000000111",
53869=>"001101000",
53870=>"110000000",
53871=>"001011010",
53872=>"111111000",
53873=>"111100110",
53874=>"010010000",
53875=>"000000001",
53876=>"011010000",
53877=>"000100000",
53878=>"010100000",
53879=>"000000111",
53880=>"000010111",
53881=>"010111111",
53882=>"111010000",
53883=>"000111111",
53884=>"111011110",
53885=>"100001001",
53886=>"111111111",
53887=>"000000010",
53888=>"001001111",
53889=>"111000111",
53890=>"000101111",
53891=>"100100111",
53892=>"000000010",
53893=>"111111111",
53894=>"000000000",
53895=>"100001000",
53896=>"100100000",
53897=>"111000111",
53898=>"101000111",
53899=>"000000111",
53900=>"000000011",
53901=>"101000111",
53902=>"111101000",
53903=>"100100000",
53904=>"101101000",
53905=>"111111001",
53906=>"000101000",
53907=>"010011101",
53908=>"001010000",
53909=>"000000010",
53910=>"010000000",
53911=>"011000000",
53912=>"110010000",
53913=>"000110111",
53914=>"000101101",
53915=>"010000101",
53916=>"110011111",
53917=>"000101111",
53918=>"000010000",
53919=>"111011000",
53920=>"101001111",
53921=>"111111111",
53922=>"011110100",
53923=>"101100111",
53924=>"000111000",
53925=>"011001010",
53926=>"000000000",
53927=>"000111010",
53928=>"001100101",
53929=>"111010000",
53930=>"111000000",
53931=>"000110011",
53932=>"101110110",
53933=>"101101111",
53934=>"111111001",
53935=>"111000001",
53936=>"000110000",
53937=>"011001000",
53938=>"110000000",
53939=>"000001111",
53940=>"000111000",
53941=>"111111000",
53942=>"000000000",
53943=>"000000111",
53944=>"110000000",
53945=>"101001001",
53946=>"000000111",
53947=>"110101111",
53948=>"000000000",
53949=>"001000101",
53950=>"000000111",
53951=>"111000000",
53952=>"111101000",
53953=>"010000000",
53954=>"111111000",
53955=>"001100000",
53956=>"100111111",
53957=>"111101001",
53958=>"100011011",
53959=>"000111111",
53960=>"000110110",
53961=>"110010011",
53962=>"111101100",
53963=>"110000000",
53964=>"010011000",
53965=>"111110111",
53966=>"000110000",
53967=>"011001110",
53968=>"111000000",
53969=>"111111100",
53970=>"111000101",
53971=>"111111011",
53972=>"111001001",
53973=>"100011000",
53974=>"111111000",
53975=>"010011000",
53976=>"111111000",
53977=>"101011110",
53978=>"101100111",
53979=>"001000111",
53980=>"111110100",
53981=>"000000000",
53982=>"111010011",
53983=>"001000001",
53984=>"000001111",
53985=>"000000000",
53986=>"111110000",
53987=>"111111001",
53988=>"000001000",
53989=>"111111001",
53990=>"000110110",
53991=>"111111111",
53992=>"111000110",
53993=>"000000000",
53994=>"110001100",
53995=>"000000000",
53996=>"000111000",
53997=>"000000101",
53998=>"000111000",
53999=>"101111110",
54000=>"001100000",
54001=>"011001100",
54002=>"111111000",
54003=>"001011000",
54004=>"111111011",
54005=>"000000000",
54006=>"100000111",
54007=>"010000100",
54008=>"101110111",
54009=>"111111001",
54010=>"101001011",
54011=>"001000000",
54012=>"111111000",
54013=>"111110000",
54014=>"000011110",
54015=>"111111000",
54016=>"011000000",
54017=>"000001000",
54018=>"000000000",
54019=>"000000000",
54020=>"000000001",
54021=>"101100110",
54022=>"010000000",
54023=>"001000010",
54024=>"000001111",
54025=>"101101111",
54026=>"001000000",
54027=>"000000111",
54028=>"111010110",
54029=>"111000110",
54030=>"000001011",
54031=>"000000000",
54032=>"111111111",
54033=>"010000111",
54034=>"000110010",
54035=>"000011111",
54036=>"000010110",
54037=>"111111111",
54038=>"000000000",
54039=>"000000000",
54040=>"010011001",
54041=>"111111111",
54042=>"111111111",
54043=>"111111010",
54044=>"111111111",
54045=>"000001001",
54046=>"000000010",
54047=>"111111111",
54048=>"100001000",
54049=>"000010000",
54050=>"000010000",
54051=>"111111111",
54052=>"000000000",
54053=>"111111110",
54054=>"111101100",
54055=>"111001101",
54056=>"111011001",
54057=>"010000000",
54058=>"001010101",
54059=>"111111111",
54060=>"010010000",
54061=>"000000000",
54062=>"001010000",
54063=>"000000001",
54064=>"000000000",
54065=>"100000000",
54066=>"001000001",
54067=>"000001111",
54068=>"010001000",
54069=>"000001000",
54070=>"111111001",
54071=>"000000111",
54072=>"000000000",
54073=>"000010000",
54074=>"011011001",
54075=>"000000111",
54076=>"000001111",
54077=>"111111110",
54078=>"000000110",
54079=>"000000011",
54080=>"100110110",
54081=>"111111010",
54082=>"111000000",
54083=>"101101110",
54084=>"110110110",
54085=>"000010010",
54086=>"010111100",
54087=>"000000111",
54088=>"001101100",
54089=>"111110100",
54090=>"000010010",
54091=>"000000011",
54092=>"111111111",
54093=>"001000001",
54094=>"001000000",
54095=>"100000000",
54096=>"111101101",
54097=>"110000011",
54098=>"001000111",
54099=>"000000000",
54100=>"010110010",
54101=>"001011100",
54102=>"000000000",
54103=>"111111111",
54104=>"000100000",
54105=>"000000000",
54106=>"101101100",
54107=>"101101011",
54108=>"001000000",
54109=>"000001001",
54110=>"111111111",
54111=>"100011011",
54112=>"101101111",
54113=>"101100101",
54114=>"111111110",
54115=>"010111010",
54116=>"101001100",
54117=>"110011011",
54118=>"011101100",
54119=>"011111111",
54120=>"000100110",
54121=>"000000010",
54122=>"111111111",
54123=>"110111111",
54124=>"111110111",
54125=>"000000010",
54126=>"111111111",
54127=>"000100011",
54128=>"001011011",
54129=>"000000000",
54130=>"111111110",
54131=>"000110111",
54132=>"111000000",
54133=>"000100100",
54134=>"000000100",
54135=>"110100100",
54136=>"111111111",
54137=>"000100111",
54138=>"000000000",
54139=>"000000000",
54140=>"000111111",
54141=>"000000001",
54142=>"001000000",
54143=>"101111111",
54144=>"111011000",
54145=>"100100000",
54146=>"111000000",
54147=>"000000000",
54148=>"000100000",
54149=>"000110010",
54150=>"111111011",
54151=>"111111111",
54152=>"111100011",
54153=>"011010000",
54154=>"000000000",
54155=>"000000011",
54156=>"111111010",
54157=>"011011001",
54158=>"000010111",
54159=>"000001111",
54160=>"001001001",
54161=>"001010000",
54162=>"111111111",
54163=>"111110101",
54164=>"011111111",
54165=>"000000101",
54166=>"110111011",
54167=>"100000000",
54168=>"111000100",
54169=>"111111111",
54170=>"111110111",
54171=>"000001100",
54172=>"011010000",
54173=>"000000000",
54174=>"111000000",
54175=>"000000000",
54176=>"011101000",
54177=>"101101000",
54178=>"111100000",
54179=>"101000110",
54180=>"111000001",
54181=>"110111111",
54182=>"000001011",
54183=>"100000011",
54184=>"010000110",
54185=>"000000000",
54186=>"101101101",
54187=>"001010110",
54188=>"001111011",
54189=>"111110111",
54190=>"000000011",
54191=>"111111111",
54192=>"101100010",
54193=>"000000011",
54194=>"000000011",
54195=>"000000000",
54196=>"000000100",
54197=>"000000011",
54198=>"011110110",
54199=>"010111001",
54200=>"011110111",
54201=>"110111111",
54202=>"111111001",
54203=>"111100111",
54204=>"000110111",
54205=>"111111111",
54206=>"001001111",
54207=>"000000110",
54208=>"111111111",
54209=>"111111011",
54210=>"000000111",
54211=>"100100100",
54212=>"111111000",
54213=>"000000111",
54214=>"100000001",
54215=>"100001010",
54216=>"111011011",
54217=>"111111111",
54218=>"110011001",
54219=>"111110110",
54220=>"000100011",
54221=>"010011111",
54222=>"100110111",
54223=>"000000000",
54224=>"000010000",
54225=>"001001011",
54226=>"111111110",
54227=>"000000000",
54228=>"011100010",
54229=>"000000001",
54230=>"110110010",
54231=>"111000011",
54232=>"111010000",
54233=>"000000111",
54234=>"000000010",
54235=>"010000000",
54236=>"011010101",
54237=>"000001100",
54238=>"110111111",
54239=>"010000000",
54240=>"010111111",
54241=>"010000000",
54242=>"111111111",
54243=>"100000100",
54244=>"110111110",
54245=>"110111111",
54246=>"111111111",
54247=>"001000100",
54248=>"100000000",
54249=>"100000000",
54250=>"000000000",
54251=>"101000111",
54252=>"111111111",
54253=>"000010010",
54254=>"000000000",
54255=>"100000000",
54256=>"101111111",
54257=>"000000011",
54258=>"001000111",
54259=>"000000000",
54260=>"100000000",
54261=>"011011000",
54262=>"010010111",
54263=>"101000100",
54264=>"111110110",
54265=>"000000000",
54266=>"000000000",
54267=>"000000111",
54268=>"000000000",
54269=>"110000110",
54270=>"000011111",
54271=>"010000000",
54272=>"110000000",
54273=>"000111111",
54274=>"101000000",
54275=>"111000010",
54276=>"100000111",
54277=>"000000000",
54278=>"101010100",
54279=>"101110110",
54280=>"101100111",
54281=>"000000100",
54282=>"000011000",
54283=>"111010110",
54284=>"111111011",
54285=>"000000000",
54286=>"000100110",
54287=>"111111010",
54288=>"110010000",
54289=>"111011111",
54290=>"111101111",
54291=>"000000100",
54292=>"101101111",
54293=>"101101101",
54294=>"110011011",
54295=>"101111011",
54296=>"010111001",
54297=>"101111100",
54298=>"000110000",
54299=>"001000111",
54300=>"101101101",
54301=>"001111111",
54302=>"011110000",
54303=>"111000000",
54304=>"111101111",
54305=>"111111111",
54306=>"000010111",
54307=>"000111111",
54308=>"101111111",
54309=>"000000011",
54310=>"000000001",
54311=>"110111111",
54312=>"111001111",
54313=>"011111111",
54314=>"000111000",
54315=>"110111011",
54316=>"000000100",
54317=>"000111111",
54318=>"101100000",
54319=>"110110111",
54320=>"111000111",
54321=>"000000111",
54322=>"111111010",
54323=>"010110101",
54324=>"000010000",
54325=>"111111110",
54326=>"001011110",
54327=>"000100111",
54328=>"110000000",
54329=>"000000011",
54330=>"110000011",
54331=>"000000000",
54332=>"001101001",
54333=>"010110110",
54334=>"000000000",
54335=>"110001110",
54336=>"100000111",
54337=>"000000111",
54338=>"001000000",
54339=>"110110001",
54340=>"111001000",
54341=>"101001001",
54342=>"001000000",
54343=>"011101000",
54344=>"110101011",
54345=>"001101001",
54346=>"111110110",
54347=>"101001100",
54348=>"100000001",
54349=>"101100100",
54350=>"011000111",
54351=>"100100000",
54352=>"101111111",
54353=>"111010000",
54354=>"111011110",
54355=>"111001001",
54356=>"011000101",
54357=>"111111100",
54358=>"111111110",
54359=>"000000000",
54360=>"111000001",
54361=>"100101011",
54362=>"000000011",
54363=>"101111110",
54364=>"001001010",
54365=>"010000110",
54366=>"111101111",
54367=>"011010100",
54368=>"000110000",
54369=>"101011000",
54370=>"101000000",
54371=>"110111111",
54372=>"101000111",
54373=>"111111111",
54374=>"111011010",
54375=>"000000010",
54376=>"101111101",
54377=>"111000000",
54378=>"111100111",
54379=>"111000000",
54380=>"100010111",
54381=>"000000000",
54382=>"000000000",
54383=>"000111000",
54384=>"010001000",
54385=>"000000110",
54386=>"100010001",
54387=>"000000000",
54388=>"011000000",
54389=>"001000100",
54390=>"000000000",
54391=>"000000000",
54392=>"111000010",
54393=>"110001000",
54394=>"001001000",
54395=>"110101110",
54396=>"111010101",
54397=>"111100100",
54398=>"001111111",
54399=>"101000001",
54400=>"101001000",
54401=>"111110010",
54402=>"101100011",
54403=>"101000111",
54404=>"100001111",
54405=>"111101101",
54406=>"001000010",
54407=>"000001001",
54408=>"001100000",
54409=>"001000101",
54410=>"111100111",
54411=>"111001000",
54412=>"100101100",
54413=>"000000100",
54414=>"010001101",
54415=>"000100000",
54416=>"011111011",
54417=>"001000000",
54418=>"000000000",
54419=>"110111000",
54420=>"011010000",
54421=>"101111000",
54422=>"111010110",
54423=>"110101111",
54424=>"111111111",
54425=>"000010101",
54426=>"111000101",
54427=>"100000000",
54428=>"010100111",
54429=>"000001001",
54430=>"111010010",
54431=>"000010001",
54432=>"001001000",
54433=>"001111110",
54434=>"000110000",
54435=>"000111111",
54436=>"010010100",
54437=>"001101110",
54438=>"001001000",
54439=>"000011001",
54440=>"000111111",
54441=>"000101111",
54442=>"111000001",
54443=>"010000011",
54444=>"100000111",
54445=>"101000101",
54446=>"011001111",
54447=>"000101101",
54448=>"110111111",
54449=>"110010100",
54450=>"110000010",
54451=>"000100010",
54452=>"110111111",
54453=>"100111111",
54454=>"110011101",
54455=>"001000000",
54456=>"000101101",
54457=>"110011000",
54458=>"101001010",
54459=>"111111000",
54460=>"000000111",
54461=>"001010100",
54462=>"001000001",
54463=>"111010000",
54464=>"111001000",
54465=>"000000000",
54466=>"101001011",
54467=>"010000111",
54468=>"001001000",
54469=>"111100000",
54470=>"000000010",
54471=>"111101100",
54472=>"000110111",
54473=>"000000001",
54474=>"111111110",
54475=>"111000001",
54476=>"000100111",
54477=>"010010100",
54478=>"000001001",
54479=>"110100100",
54480=>"000000110",
54481=>"011101111",
54482=>"100110111",
54483=>"110111101",
54484=>"101001000",
54485=>"011110010",
54486=>"000010000",
54487=>"000000111",
54488=>"000111111",
54489=>"000001001",
54490=>"110101000",
54491=>"111000100",
54492=>"111100110",
54493=>"101010010",
54494=>"011010000",
54495=>"111101011",
54496=>"001000110",
54497=>"011100010",
54498=>"111000011",
54499=>"111001111",
54500=>"001101101",
54501=>"111000000",
54502=>"000000000",
54503=>"100000101",
54504=>"001001011",
54505=>"000111000",
54506=>"011010000",
54507=>"001000000",
54508=>"000010111",
54509=>"111111000",
54510=>"000000000",
54511=>"001000000",
54512=>"000000110",
54513=>"001001101",
54514=>"101001110",
54515=>"011011111",
54516=>"001100000",
54517=>"000100101",
54518=>"101000000",
54519=>"000000010",
54520=>"000100000",
54521=>"010110110",
54522=>"111110000",
54523=>"010100010",
54524=>"011000101",
54525=>"111000111",
54526=>"011011111",
54527=>"000000100",
54528=>"011001001",
54529=>"110100100",
54530=>"110000110",
54531=>"100000000",
54532=>"100111011",
54533=>"000000010",
54534=>"000000000",
54535=>"110111111",
54536=>"000110100",
54537=>"000011011",
54538=>"010001011",
54539=>"000011011",
54540=>"000100100",
54541=>"100100111",
54542=>"010111001",
54543=>"001000100",
54544=>"011011000",
54545=>"100100010",
54546=>"100000011",
54547=>"000101111",
54548=>"111111010",
54549=>"011000100",
54550=>"011100100",
54551=>"000111111",
54552=>"000011010",
54553=>"111011011",
54554=>"111011010",
54555=>"100000000",
54556=>"000100100",
54557=>"110011111",
54558=>"010011010",
54559=>"100000000",
54560=>"111101000",
54561=>"110100100",
54562=>"111101111",
54563=>"000100101",
54564=>"100011001",
54565=>"011010010",
54566=>"111011010",
54567=>"000000000",
54568=>"111000000",
54569=>"111111100",
54570=>"000100100",
54571=>"000000000",
54572=>"111110111",
54573=>"111111111",
54574=>"011011110",
54575=>"000000111",
54576=>"111000000",
54577=>"111011100",
54578=>"011100000",
54579=>"111110000",
54580=>"101000000",
54581=>"011000111",
54582=>"000110101",
54583=>"000000011",
54584=>"000100001",
54585=>"000100100",
54586=>"011100110",
54587=>"000000000",
54588=>"100111001",
54589=>"011100000",
54590=>"100000000",
54591=>"000011011",
54592=>"111111000",
54593=>"111011000",
54594=>"111110101",
54595=>"000011011",
54596=>"011000100",
54597=>"011000000",
54598=>"000100000",
54599=>"111100111",
54600=>"011111110",
54601=>"001011011",
54602=>"111011000",
54603=>"111100100",
54604=>"011011011",
54605=>"001011000",
54606=>"000110110",
54607=>"011111100",
54608=>"001100000",
54609=>"011101001",
54610=>"111110111",
54611=>"010101100",
54612=>"000111011",
54613=>"000011011",
54614=>"000110010",
54615=>"000011011",
54616=>"111010100",
54617=>"010110110",
54618=>"000001000",
54619=>"011011011",
54620=>"000000000",
54621=>"011100010",
54622=>"111100100",
54623=>"110011011",
54624=>"100100100",
54625=>"001111111",
54626=>"111000100",
54627=>"001110111",
54628=>"000010000",
54629=>"110110000",
54630=>"100011000",
54631=>"001011011",
54632=>"000111111",
54633=>"101110011",
54634=>"011011001",
54635=>"111111101",
54636=>"100000110",
54637=>"101100011",
54638=>"000110000",
54639=>"111100000",
54640=>"101001001",
54641=>"001010111",
54642=>"001001000",
54643=>"111000100",
54644=>"011010000",
54645=>"001000000",
54646=>"000000011",
54647=>"011011011",
54648=>"111000000",
54649=>"100100011",
54650=>"111100100",
54651=>"000000101",
54652=>"000110010",
54653=>"011110000",
54654=>"010000000",
54655=>"000111011",
54656=>"111000101",
54657=>"000011011",
54658=>"011011000",
54659=>"110100001",
54660=>"011011100",
54661=>"110111111",
54662=>"011111001",
54663=>"000010011",
54664=>"110110011",
54665=>"110111100",
54666=>"011000000",
54667=>"100000110",
54668=>"000011010",
54669=>"000000101",
54670=>"000001111",
54671=>"000000000",
54672=>"011101110",
54673=>"000010010",
54674=>"000011000",
54675=>"110100000",
54676=>"010111111",
54677=>"000000000",
54678=>"111111111",
54679=>"010000100",
54680=>"000100000",
54681=>"011111011",
54682=>"001001000",
54683=>"010000100",
54684=>"110100100",
54685=>"001011010",
54686=>"101101110",
54687=>"011000000",
54688=>"100010111",
54689=>"100111111",
54690=>"110000000",
54691=>"000101000",
54692=>"011101000",
54693=>"001111111",
54694=>"101100111",
54695=>"001100100",
54696=>"010000110",
54697=>"000100000",
54698=>"100100110",
54699=>"010000100",
54700=>"111000111",
54701=>"001011000",
54702=>"001100000",
54703=>"000000100",
54704=>"100111110",
54705=>"101000100",
54706=>"001111111",
54707=>"001100000",
54708=>"000111111",
54709=>"110100111",
54710=>"011111101",
54711=>"011100000",
54712=>"011011010",
54713=>"000111011",
54714=>"000011001",
54715=>"011011001",
54716=>"111111100",
54717=>"011000000",
54718=>"010010111",
54719=>"001000010",
54720=>"010011010",
54721=>"100011011",
54722=>"011000011",
54723=>"100010110",
54724=>"000000000",
54725=>"110000000",
54726=>"000000011",
54727=>"101111011",
54728=>"100111110",
54729=>"000011011",
54730=>"111101111",
54731=>"000011000",
54732=>"000011001",
54733=>"000001011",
54734=>"000000011",
54735=>"100111011",
54736=>"000000111",
54737=>"011001001",
54738=>"110111011",
54739=>"000000100",
54740=>"111000100",
54741=>"110100100",
54742=>"000100010",
54743=>"110000000",
54744=>"110100011",
54745=>"100100100",
54746=>"100000100",
54747=>"111100111",
54748=>"110111111",
54749=>"110101011",
54750=>"010000000",
54751=>"010011000",
54752=>"000000000",
54753=>"010100100",
54754=>"000111011",
54755=>"101111111",
54756=>"100011000",
54757=>"111100101",
54758=>"000000000",
54759=>"000110001",
54760=>"001000111",
54761=>"110000000",
54762=>"000010000",
54763=>"010101111",
54764=>"000000100",
54765=>"000000111",
54766=>"000000000",
54767=>"000001001",
54768=>"111111011",
54769=>"001001101",
54770=>"000000011",
54771=>"001001101",
54772=>"101101010",
54773=>"000000100",
54774=>"000000001",
54775=>"000000101",
54776=>"000100000",
54777=>"100110011",
54778=>"010000110",
54779=>"000001111",
54780=>"111100100",
54781=>"010011011",
54782=>"010110000",
54783=>"110000000",
54784=>"000011100",
54785=>"000000010",
54786=>"010010010",
54787=>"001101111",
54788=>"000000011",
54789=>"000000001",
54790=>"011111111",
54791=>"110111011",
54792=>"000000100",
54793=>"111010101",
54794=>"111111111",
54795=>"110111010",
54796=>"000111111",
54797=>"000101000",
54798=>"111111110",
54799=>"111111111",
54800=>"000000111",
54801=>"111110111",
54802=>"111110110",
54803=>"111000111",
54804=>"011111101",
54805=>"000000101",
54806=>"011111101",
54807=>"111111111",
54808=>"000001100",
54809=>"000000111",
54810=>"000000000",
54811=>"010100100",
54812=>"000000000",
54813=>"111101000",
54814=>"001111111",
54815=>"101100000",
54816=>"000111101",
54817=>"110111000",
54818=>"001101100",
54819=>"000010011",
54820=>"001011111",
54821=>"000001001",
54822=>"000111110",
54823=>"110111111",
54824=>"111011110",
54825=>"000000000",
54826=>"111111101",
54827=>"000000100",
54828=>"000001011",
54829=>"000000010",
54830=>"000000110",
54831=>"110011000",
54832=>"000101001",
54833=>"110110111",
54834=>"000101001",
54835=>"001101000",
54836=>"110111111",
54837=>"000110001",
54838=>"111111111",
54839=>"101111100",
54840=>"000101111",
54841=>"111101000",
54842=>"111101000",
54843=>"000101111",
54844=>"000000000",
54845=>"111111111",
54846=>"000101111",
54847=>"100100100",
54848=>"000001111",
54849=>"000000000",
54850=>"101001101",
54851=>"111111111",
54852=>"111111111",
54853=>"000000111",
54854=>"111110111",
54855=>"000001011",
54856=>"000000000",
54857=>"111101000",
54858=>"111101101",
54859=>"110000010",
54860=>"000000000",
54861=>"110100111",
54862=>"001010110",
54863=>"000000111",
54864=>"111111111",
54865=>"100011101",
54866=>"001011001",
54867=>"000001000",
54868=>"000010010",
54869=>"000001000",
54870=>"111011010",
54871=>"110111111",
54872=>"001000101",
54873=>"110100101",
54874=>"111101011",
54875=>"111000111",
54876=>"000000000",
54877=>"100100111",
54878=>"000000111",
54879=>"110111111",
54880=>"000011000",
54881=>"010010000",
54882=>"110111111",
54883=>"111011000",
54884=>"001000101",
54885=>"011100000",
54886=>"000000000",
54887=>"111111100",
54888=>"111111110",
54889=>"111101000",
54890=>"000100000",
54891=>"001000000",
54892=>"000111111",
54893=>"111011011",
54894=>"111111101",
54895=>"111011000",
54896=>"011011011",
54897=>"010101000",
54898=>"111111111",
54899=>"000000000",
54900=>"011110000",
54901=>"000000000",
54902=>"000111100",
54903=>"000111111",
54904=>"010110110",
54905=>"111111000",
54906=>"111110000",
54907=>"001101111",
54908=>"111111111",
54909=>"011000001",
54910=>"111101111",
54911=>"010010011",
54912=>"001001010",
54913=>"011000101",
54914=>"000000000",
54915=>"101111101",
54916=>"010110010",
54917=>"000000000",
54918=>"000000100",
54919=>"101000110",
54920=>"000100111",
54921=>"111011010",
54922=>"000000000",
54923=>"101000010",
54924=>"001000010",
54925=>"000010000",
54926=>"000000000",
54927=>"010110011",
54928=>"111101100",
54929=>"100000000",
54930=>"100011011",
54931=>"111110000",
54932=>"000000000",
54933=>"111111111",
54934=>"000000010",
54935=>"000100000",
54936=>"000010010",
54937=>"101001000",
54938=>"110110010",
54939=>"000010011",
54940=>"000110111",
54941=>"000000111",
54942=>"010001001",
54943=>"011011000",
54944=>"000000100",
54945=>"000111000",
54946=>"000000100",
54947=>"111111111",
54948=>"110111111",
54949=>"001010011",
54950=>"001000000",
54951=>"000000111",
54952=>"111100000",
54953=>"000000000",
54954=>"110100100",
54955=>"011111111",
54956=>"001011000",
54957=>"111010000",
54958=>"111101111",
54959=>"001000000",
54960=>"000000001",
54961=>"111011001",
54962=>"000110010",
54963=>"011111111",
54964=>"111100100",
54965=>"111111010",
54966=>"000111011",
54967=>"000000101",
54968=>"000000000",
54969=>"000010001",
54970=>"000000000",
54971=>"000111111",
54972=>"000000000",
54973=>"111111111",
54974=>"000001000",
54975=>"111011000",
54976=>"000000111",
54977=>"111000111",
54978=>"001000011",
54979=>"110110010",
54980=>"000001111",
54981=>"100001000",
54982=>"111111111",
54983=>"000001000",
54984=>"111101101",
54985=>"000011010",
54986=>"010101111",
54987=>"010010111",
54988=>"100100000",
54989=>"111111011",
54990=>"111111111",
54991=>"111111111",
54992=>"111111111",
54993=>"000010000",
54994=>"101000001",
54995=>"111111010",
54996=>"000000011",
54997=>"011111101",
54998=>"000011000",
54999=>"011101000",
55000=>"000000000",
55001=>"111010000",
55002=>"001001000",
55003=>"111111111",
55004=>"101111000",
55005=>"111000000",
55006=>"111100110",
55007=>"001000000",
55008=>"111111110",
55009=>"011101000",
55010=>"101000001",
55011=>"011011011",
55012=>"111000000",
55013=>"000000000",
55014=>"000000000",
55015=>"111111111",
55016=>"000100110",
55017=>"101111110",
55018=>"111111111",
55019=>"000111111",
55020=>"000111111",
55021=>"010111010",
55022=>"111110000",
55023=>"100000000",
55024=>"000000010",
55025=>"000000000",
55026=>"000011000",
55027=>"011001000",
55028=>"001100101",
55029=>"111111111",
55030=>"000011111",
55031=>"101101111",
55032=>"011111111",
55033=>"111111111",
55034=>"000000001",
55035=>"001000000",
55036=>"000100110",
55037=>"111010110",
55038=>"110001110",
55039=>"000111111",
55040=>"011001100",
55041=>"111100100",
55042=>"111100100",
55043=>"000101111",
55044=>"111110111",
55045=>"111110101",
55046=>"000011011",
55047=>"001100010",
55048=>"000000110",
55049=>"000000000",
55050=>"010110011",
55051=>"101011111",
55052=>"000100010",
55053=>"000010000",
55054=>"110110110",
55055=>"000110010",
55056=>"100111101",
55057=>"000011010",
55058=>"111001010",
55059=>"010000000",
55060=>"001100100",
55061=>"111101101",
55062=>"111101101",
55063=>"101111111",
55064=>"111101000",
55065=>"111111010",
55066=>"011111111",
55067=>"001101110",
55068=>"011111111",
55069=>"000011111",
55070=>"010101101",
55071=>"011111110",
55072=>"111101101",
55073=>"111100100",
55074=>"101100110",
55075=>"111100001",
55076=>"011110110",
55077=>"001100111",
55078=>"110100100",
55079=>"000001010",
55080=>"111101111",
55081=>"101100111",
55082=>"100010011",
55083=>"111011110",
55084=>"000110111",
55085=>"011011000",
55086=>"101111100",
55087=>"110110100",
55088=>"010111101",
55089=>"111111001",
55090=>"001111111",
55091=>"110111111",
55092=>"000000100",
55093=>"110010100",
55094=>"101100000",
55095=>"000000000",
55096=>"011111110",
55097=>"000000000",
55098=>"100100010",
55099=>"110011000",
55100=>"011000110",
55101=>"111111000",
55102=>"111100100",
55103=>"000111011",
55104=>"000101001",
55105=>"000110100",
55106=>"010100100",
55107=>"111111000",
55108=>"000010010",
55109=>"000000000",
55110=>"000000000",
55111=>"001101011",
55112=>"011101000",
55113=>"100101111",
55114=>"110110101",
55115=>"100111011",
55116=>"111101011",
55117=>"100101111",
55118=>"101100110",
55119=>"110110100",
55120=>"111111000",
55121=>"111100100",
55122=>"000010111",
55123=>"000011011",
55124=>"010000101",
55125=>"011000100",
55126=>"000010010",
55127=>"111000100",
55128=>"100111110",
55129=>"000000001",
55130=>"011101011",
55131=>"000000110",
55132=>"000010010",
55133=>"011011000",
55134=>"111111101",
55135=>"111100000",
55136=>"111111111",
55137=>"000000000",
55138=>"100000100",
55139=>"011110000",
55140=>"111000100",
55141=>"111000100",
55142=>"000000000",
55143=>"101001011",
55144=>"011000111",
55145=>"010100111",
55146=>"111111011",
55147=>"100101111",
55148=>"010000100",
55149=>"010010010",
55150=>"000000000",
55151=>"000001010",
55152=>"100111111",
55153=>"000101100",
55154=>"110001000",
55155=>"001111111",
55156=>"000000000",
55157=>"010000100",
55158=>"010111111",
55159=>"100100000",
55160=>"111111000",
55161=>"100110010",
55162=>"000101000",
55163=>"000111100",
55164=>"111111011",
55165=>"011000000",
55166=>"111100101",
55167=>"111111101",
55168=>"100011000",
55169=>"111000000",
55170=>"110110100",
55171=>"000100111",
55172=>"111111111",
55173=>"111000010",
55174=>"100100100",
55175=>"010100000",
55176=>"010111111",
55177=>"010000000",
55178=>"100000000",
55179=>"100000011",
55180=>"011100000",
55181=>"000100000",
55182=>"111111110",
55183=>"010000000",
55184=>"101100001",
55185=>"011001101",
55186=>"000000000",
55187=>"111101101",
55188=>"010111101",
55189=>"001101101",
55190=>"100111111",
55191=>"101011100",
55192=>"000000101",
55193=>"010111110",
55194=>"000001110",
55195=>"101100000",
55196=>"111100100",
55197=>"110101101",
55198=>"000000110",
55199=>"001111110",
55200=>"110111010",
55201=>"111011100",
55202=>"000111010",
55203=>"110111111",
55204=>"111101111",
55205=>"000110010",
55206=>"100100101",
55207=>"000000111",
55208=>"000111011",
55209=>"000001000",
55210=>"111100000",
55211=>"111100000",
55212=>"101010011",
55213=>"010011010",
55214=>"011000000",
55215=>"000010000",
55216=>"100011011",
55217=>"111111111",
55218=>"000010000",
55219=>"110011000",
55220=>"000001011",
55221=>"100111000",
55222=>"000011010",
55223=>"011100000",
55224=>"110110000",
55225=>"000110101",
55226=>"010000000",
55227=>"010110111",
55228=>"010000011",
55229=>"011111111",
55230=>"000011011",
55231=>"010111101",
55232=>"110010000",
55233=>"111111111",
55234=>"111010000",
55235=>"100001011",
55236=>"011010010",
55237=>"110001101",
55238=>"000000011",
55239=>"011100101",
55240=>"011101000",
55241=>"111000100",
55242=>"111111011",
55243=>"111000100",
55244=>"001011000",
55245=>"111100111",
55246=>"101010010",
55247=>"011101100",
55248=>"100000000",
55249=>"010111011",
55250=>"000100111",
55251=>"000011011",
55252=>"000000000",
55253=>"111100001",
55254=>"111101100",
55255=>"100000101",
55256=>"000011001",
55257=>"010111000",
55258=>"011111110",
55259=>"101110000",
55260=>"111100001",
55261=>"001111000",
55262=>"000011011",
55263=>"000010000",
55264=>"001100000",
55265=>"110100000",
55266=>"110111111",
55267=>"000100110",
55268=>"111100111",
55269=>"100100101",
55270=>"000111010",
55271=>"100100000",
55272=>"011011011",
55273=>"000010010",
55274=>"100100010",
55275=>"100000100",
55276=>"011010101",
55277=>"100111111",
55278=>"111000000",
55279=>"000111111",
55280=>"010011011",
55281=>"011100100",
55282=>"000101100",
55283=>"100110110",
55284=>"101000100",
55285=>"111101000",
55286=>"100000010",
55287=>"001010011",
55288=>"111111100",
55289=>"111111011",
55290=>"111111111",
55291=>"000110111",
55292=>"000101011",
55293=>"011011111",
55294=>"011011111",
55295=>"111101001",
55296=>"100001000",
55297=>"101100100",
55298=>"000000000",
55299=>"001000111",
55300=>"000000110",
55301=>"000110010",
55302=>"111011111",
55303=>"110101000",
55304=>"110010000",
55305=>"110010010",
55306=>"000110010",
55307=>"000001011",
55308=>"111101001",
55309=>"100001001",
55310=>"000100101",
55311=>"111101000",
55312=>"111110111",
55313=>"111010010",
55314=>"010000000",
55315=>"001010010",
55316=>"000101111",
55317=>"101001001",
55318=>"100100000",
55319=>"110111110",
55320=>"111000010",
55321=>"110111111",
55322=>"111111111",
55323=>"101000110",
55324=>"111100100",
55325=>"110000000",
55326=>"111111001",
55327=>"010000000",
55328=>"111010000",
55329=>"000010110",
55330=>"010000001",
55331=>"111011010",
55332=>"000110110",
55333=>"000100001",
55334=>"111110010",
55335=>"000110110",
55336=>"000011111",
55337=>"111111110",
55338=>"101111010",
55339=>"010010001",
55340=>"100111100",
55341=>"101111011",
55342=>"010000100",
55343=>"000000100",
55344=>"010010000",
55345=>"010001100",
55346=>"010010111",
55347=>"000000101",
55348=>"100110010",
55349=>"000111111",
55350=>"011011011",
55351=>"000100000",
55352=>"111010001",
55353=>"111001000",
55354=>"000000101",
55355=>"100010010",
55356=>"110000100",
55357=>"111001000",
55358=>"110010000",
55359=>"000001111",
55360=>"111110000",
55361=>"111110010",
55362=>"111000000",
55363=>"110000000",
55364=>"111111000",
55365=>"000101111",
55366=>"000101011",
55367=>"011010111",
55368=>"111110011",
55369=>"111110000",
55370=>"111000000",
55371=>"000011110",
55372=>"000000000",
55373=>"010011000",
55374=>"000101000",
55375=>"000000101",
55376=>"000010010",
55377=>"111111111",
55378=>"101111001",
55379=>"000011000",
55380=>"111000010",
55381=>"100100100",
55382=>"000011111",
55383=>"111010110",
55384=>"010000001",
55385=>"011010011",
55386=>"000100110",
55387=>"010001011",
55388=>"000111101",
55389=>"010000000",
55390=>"111111111",
55391=>"001000000",
55392=>"111111000",
55393=>"000000000",
55394=>"111010000",
55395=>"000010001",
55396=>"100000001",
55397=>"000001011",
55398=>"101000000",
55399=>"000001101",
55400=>"111000111",
55401=>"111101101",
55402=>"000010111",
55403=>"000100000",
55404=>"111000100",
55405=>"000110110",
55406=>"000001001",
55407=>"000000000",
55408=>"000100100",
55409=>"000000000",
55410=>"110110110",
55411=>"000000000",
55412=>"001001001",
55413=>"101000000",
55414=>"111001101",
55415=>"111000000",
55416=>"111001010",
55417=>"000000000",
55418=>"001010111",
55419=>"000001001",
55420=>"110100000",
55421=>"000100000",
55422=>"000010010",
55423=>"000000000",
55424=>"101111111",
55425=>"111111000",
55426=>"000101000",
55427=>"010000010",
55428=>"110011100",
55429=>"000110111",
55430=>"001001100",
55431=>"000101001",
55432=>"001001001",
55433=>"001000011",
55434=>"000101111",
55435=>"010000101",
55436=>"000100000",
55437=>"000001000",
55438=>"101101101",
55439=>"001000100",
55440=>"011000000",
55441=>"111000011",
55442=>"000111110",
55443=>"011011001",
55444=>"101100011",
55445=>"111010000",
55446=>"011111100",
55447=>"000100100",
55448=>"000101110",
55449=>"101101111",
55450=>"111101110",
55451=>"111010000",
55452=>"111000111",
55453=>"111000000",
55454=>"101111011",
55455=>"111000000",
55456=>"000011011",
55457=>"101010000",
55458=>"001000010",
55459=>"101011010",
55460=>"000000010",
55461=>"000100100",
55462=>"000000000",
55463=>"000110110",
55464=>"001100010",
55465=>"000000000",
55466=>"011101000",
55467=>"111010000",
55468=>"110100110",
55469=>"000000000",
55470=>"000000000",
55471=>"000000000",
55472=>"111101000",
55473=>"000111111",
55474=>"010000000",
55475=>"110110110",
55476=>"100110111",
55477=>"111011111",
55478=>"010100101",
55479=>"000110111",
55480=>"111001011",
55481=>"111001100",
55482=>"000101110",
55483=>"111001010",
55484=>"101101101",
55485=>"010111011",
55486=>"110010000",
55487=>"010111000",
55488=>"001000101",
55489=>"000101100",
55490=>"101111011",
55491=>"110100100",
55492=>"001000111",
55493=>"000100000",
55494=>"111101001",
55495=>"111000000",
55496=>"000100101",
55497=>"101101000",
55498=>"000111111",
55499=>"001111111",
55500=>"000000000",
55501=>"111011000",
55502=>"010111000",
55503=>"000001111",
55504=>"000000000",
55505=>"000001001",
55506=>"000100110",
55507=>"111111000",
55508=>"111101001",
55509=>"000011011",
55510=>"101110000",
55511=>"000110111",
55512=>"001101111",
55513=>"001000110",
55514=>"010100100",
55515=>"010110111",
55516=>"110101001",
55517=>"000001100",
55518=>"000001001",
55519=>"010011010",
55520=>"010000001",
55521=>"111000101",
55522=>"000101111",
55523=>"011111111",
55524=>"101011000",
55525=>"010100111",
55526=>"001001001",
55527=>"000001000",
55528=>"111001001",
55529=>"000011010",
55530=>"000010111",
55531=>"111111000",
55532=>"101101111",
55533=>"000111000",
55534=>"010111000",
55535=>"000000000",
55536=>"000010000",
55537=>"000001001",
55538=>"101000000",
55539=>"000111111",
55540=>"000100100",
55541=>"000001001",
55542=>"000100000",
55543=>"111000111",
55544=>"101010111",
55545=>"010111101",
55546=>"011111111",
55547=>"000000001",
55548=>"111111001",
55549=>"000101111",
55550=>"000000011",
55551=>"000000000",
55552=>"001011011",
55553=>"000000000",
55554=>"111000000",
55555=>"100100111",
55556=>"001011011",
55557=>"111101001",
55558=>"100000100",
55559=>"111001010",
55560=>"000100100",
55561=>"000000100",
55562=>"101001111",
55563=>"010000111",
55564=>"110000101",
55565=>"111111100",
55566=>"010011110",
55567=>"101000110",
55568=>"000000010",
55569=>"101011111",
55570=>"111100111",
55571=>"011000000",
55572=>"111011000",
55573=>"100111011",
55574=>"111000011",
55575=>"111001011",
55576=>"111000000",
55577=>"000000000",
55578=>"000100000",
55579=>"110100100",
55580=>"101100000",
55581=>"100100000",
55582=>"010110110",
55583=>"000110110",
55584=>"000000000",
55585=>"000111111",
55586=>"000111111",
55587=>"000011010",
55588=>"011111001",
55589=>"111011000",
55590=>"000010000",
55591=>"100010000",
55592=>"111001111",
55593=>"101001001",
55594=>"000000101",
55595=>"000011010",
55596=>"110100100",
55597=>"000000001",
55598=>"011111100",
55599=>"000111010",
55600=>"111110100",
55601=>"001101011",
55602=>"111011001",
55603=>"111110010",
55604=>"111101111",
55605=>"010111011",
55606=>"110111000",
55607=>"000100110",
55608=>"111110111",
55609=>"111000001",
55610=>"111111000",
55611=>"001001011",
55612=>"111010100",
55613=>"110111011",
55614=>"000000100",
55615=>"011011001",
55616=>"010011001",
55617=>"000010010",
55618=>"111110000",
55619=>"011000100",
55620=>"000011011",
55621=>"101000100",
55622=>"101000011",
55623=>"000000000",
55624=>"100111111",
55625=>"111000000",
55626=>"111000100",
55627=>"101100101",
55628=>"111011010",
55629=>"110111110",
55630=>"001001011",
55631=>"100000011",
55632=>"000000000",
55633=>"110111000",
55634=>"000000001",
55635=>"000011100",
55636=>"111101000",
55637=>"111101100",
55638=>"111111111",
55639=>"100000001",
55640=>"010111111",
55641=>"011001000",
55642=>"101011011",
55643=>"011011000",
55644=>"000010110",
55645=>"101000111",
55646=>"111110111",
55647=>"000001000",
55648=>"011011000",
55649=>"000000010",
55650=>"111000001",
55651=>"111111111",
55652=>"001000011",
55653=>"011111011",
55654=>"010001000",
55655=>"000011011",
55656=>"100000111",
55657=>"101011010",
55658=>"001100000",
55659=>"000111000",
55660=>"000111111",
55661=>"100000011",
55662=>"111111000",
55663=>"101000101",
55664=>"010111110",
55665=>"000011100",
55666=>"001000010",
55667=>"000010001",
55668=>"111100001",
55669=>"101100010",
55670=>"111001000",
55671=>"001011011",
55672=>"111011111",
55673=>"110001111",
55674=>"100101111",
55675=>"000101111",
55676=>"110100000",
55677=>"010100100",
55678=>"110111100",
55679=>"111000000",
55680=>"000010011",
55681=>"111000000",
55682=>"111111101",
55683=>"000001011",
55684=>"100100000",
55685=>"011001001",
55686=>"001010000",
55687=>"101100000",
55688=>"010000001",
55689=>"100111010",
55690=>"000000000",
55691=>"010010000",
55692=>"100110000",
55693=>"101100001",
55694=>"111000101",
55695=>"110000100",
55696=>"111111110",
55697=>"111011011",
55698=>"101000000",
55699=>"100111100",
55700=>"000100000",
55701=>"010000100",
55702=>"011000001",
55703=>"000010001",
55704=>"111011111",
55705=>"111111100",
55706=>"011011000",
55707=>"000100100",
55708=>"111100100",
55709=>"001001111",
55710=>"011110100",
55711=>"010011001",
55712=>"010010001",
55713=>"001000000",
55714=>"110000001",
55715=>"110111110",
55716=>"000111101",
55717=>"110011011",
55718=>"000110110",
55719=>"010011111",
55720=>"101110000",
55721=>"100100000",
55722=>"101100000",
55723=>"101010110",
55724=>"100000011",
55725=>"101100100",
55726=>"001000110",
55727=>"000100111",
55728=>"011101101",
55729=>"010000000",
55730=>"111101010",
55731=>"111010010",
55732=>"000001001",
55733=>"011000000",
55734=>"000011011",
55735=>"000011011",
55736=>"000000100",
55737=>"100101001",
55738=>"010001100",
55739=>"111101101",
55740=>"011010000",
55741=>"111111111",
55742=>"001001000",
55743=>"110111101",
55744=>"100011001",
55745=>"000000010",
55746=>"101111100",
55747=>"001010110",
55748=>"100101110",
55749=>"001001011",
55750=>"000110101",
55751=>"111111101",
55752=>"111000011",
55753=>"000011011",
55754=>"110111111",
55755=>"100100111",
55756=>"011000000",
55757=>"001001100",
55758=>"001000000",
55759=>"100001101",
55760=>"000010111",
55761=>"000000011",
55762=>"111100100",
55763=>"100001111",
55764=>"001010000",
55765=>"101000000",
55766=>"111100100",
55767=>"011111111",
55768=>"000000001",
55769=>"010000011",
55770=>"011001111",
55771=>"111000101",
55772=>"001101001",
55773=>"101111111",
55774=>"011111011",
55775=>"111100101",
55776=>"100010010",
55777=>"111111111",
55778=>"010000011",
55779=>"001000110",
55780=>"010000100",
55781=>"111111100",
55782=>"000111000",
55783=>"100001110",
55784=>"010011000",
55785=>"100110101",
55786=>"100000100",
55787=>"100000101",
55788=>"010011111",
55789=>"010011001",
55790=>"110000000",
55791=>"000011011",
55792=>"010101000",
55793=>"100100110",
55794=>"011010101",
55795=>"100100110",
55796=>"100110110",
55797=>"111000001",
55798=>"000000000",
55799=>"111100000",
55800=>"000101101",
55801=>"111101011",
55802=>"000100111",
55803=>"000000101",
55804=>"000000011",
55805=>"011000011",
55806=>"010110010",
55807=>"110000000",
55808=>"110110110",
55809=>"111111100",
55810=>"111100000",
55811=>"000011110",
55812=>"111111111",
55813=>"111011111",
55814=>"001000010",
55815=>"100111111",
55816=>"000001001",
55817=>"010000000",
55818=>"111111110",
55819=>"100101010",
55820=>"000000000",
55821=>"000000111",
55822=>"001110001",
55823=>"000000000",
55824=>"000100000",
55825=>"111111000",
55826=>"110000000",
55827=>"000011000",
55828=>"011111111",
55829=>"101100000",
55830=>"111111110",
55831=>"111111001",
55832=>"100100001",
55833=>"010001001",
55834=>"101101111",
55835=>"111111111",
55836=>"111111111",
55837=>"011111111",
55838=>"000101011",
55839=>"000101111",
55840=>"111111110",
55841=>"000111111",
55842=>"000000000",
55843=>"011111010",
55844=>"100110100",
55845=>"000000001",
55846=>"111111111",
55847=>"010111010",
55848=>"111111100",
55849=>"111111111",
55850=>"000000000",
55851=>"000000000",
55852=>"100110101",
55853=>"000000000",
55854=>"111111000",
55855=>"001010111",
55856=>"111101111",
55857=>"111111101",
55858=>"100000000",
55859=>"111111111",
55860=>"111111110",
55861=>"000101000",
55862=>"000000110",
55863=>"000000101",
55864=>"010110000",
55865=>"000000000",
55866=>"000100111",
55867=>"111111111",
55868=>"100000000",
55869=>"111011001",
55870=>"111000000",
55871=>"000001100",
55872=>"111111111",
55873=>"000000000",
55874=>"000011110",
55875=>"100111111",
55876=>"000000100",
55877=>"000001011",
55878=>"111111111",
55879=>"000000000",
55880=>"000000000",
55881=>"010110000",
55882=>"001000001",
55883=>"000000001",
55884=>"000000000",
55885=>"011111111",
55886=>"110111111",
55887=>"111111111",
55888=>"000101111",
55889=>"111010111",
55890=>"000011001",
55891=>"110000100",
55892=>"111111110",
55893=>"000001000",
55894=>"111111110",
55895=>"110110010",
55896=>"111101101",
55897=>"001001011",
55898=>"010011011",
55899=>"000000000",
55900=>"000010000",
55901=>"111000100",
55902=>"111111100",
55903=>"111011010",
55904=>"000111111",
55905=>"100001000",
55906=>"110111110",
55907=>"110111110",
55908=>"000000000",
55909=>"111001100",
55910=>"000000010",
55911=>"111111111",
55912=>"110000000",
55913=>"000000111",
55914=>"010001000",
55915=>"000000001",
55916=>"111111110",
55917=>"000000000",
55918=>"000000111",
55919=>"111000110",
55920=>"010010111",
55921=>"000000000",
55922=>"000000111",
55923=>"010000001",
55924=>"000010000",
55925=>"100001111",
55926=>"000110000",
55927=>"000001011",
55928=>"111111101",
55929=>"101100000",
55930=>"000011110",
55931=>"000000001",
55932=>"111011011",
55933=>"001000011",
55934=>"111011101",
55935=>"000000000",
55936=>"011001000",
55937=>"111000000",
55938=>"000011110",
55939=>"010111111",
55940=>"000000000",
55941=>"111101100",
55942=>"000000001",
55943=>"000000000",
55944=>"000101011",
55945=>"111000111",
55946=>"111111111",
55947=>"001011111",
55948=>"001000000",
55949=>"000011001",
55950=>"011011011",
55951=>"000001001",
55952=>"000110110",
55953=>"111000000",
55954=>"000000000",
55955=>"111101101",
55956=>"000001011",
55957=>"000000000",
55958=>"000111001",
55959=>"110010110",
55960=>"000101110",
55961=>"000000110",
55962=>"111101010",
55963=>"111010001",
55964=>"011011001",
55965=>"100100000",
55966=>"010010010",
55967=>"111111010",
55968=>"000000000",
55969=>"111010111",
55970=>"111011001",
55971=>"000000000",
55972=>"010011111",
55973=>"000010011",
55974=>"111011111",
55975=>"000000100",
55976=>"111111100",
55977=>"000100111",
55978=>"000000100",
55979=>"101111101",
55980=>"001000111",
55981=>"000000010",
55982=>"011001011",
55983=>"000000001",
55984=>"000110100",
55985=>"000000000",
55986=>"010011001",
55987=>"100100000",
55988=>"110111110",
55989=>"110011011",
55990=>"111111111",
55991=>"111111000",
55992=>"000000000",
55993=>"000100100",
55994=>"000000011",
55995=>"101101111",
55996=>"111111000",
55997=>"000000000",
55998=>"000001111",
55999=>"111100111",
56000=>"000000000",
56001=>"011000001",
56002=>"000011010",
56003=>"000101100",
56004=>"000000000",
56005=>"000011000",
56006=>"000000000",
56007=>"111101000",
56008=>"111101111",
56009=>"111111111",
56010=>"111111111",
56011=>"010111000",
56012=>"000000000",
56013=>"001011100",
56014=>"011011111",
56015=>"110111011",
56016=>"110000000",
56017=>"010011111",
56018=>"010000001",
56019=>"100111100",
56020=>"000000000",
56021=>"111110011",
56022=>"111111010",
56023=>"110111111",
56024=>"111111000",
56025=>"001111111",
56026=>"000000001",
56027=>"110000110",
56028=>"110101001",
56029=>"000101111",
56030=>"111111111",
56031=>"000000100",
56032=>"010110000",
56033=>"101111110",
56034=>"000000000",
56035=>"111110100",
56036=>"000010000",
56037=>"000001000",
56038=>"110101011",
56039=>"110000000",
56040=>"000111111",
56041=>"111111111",
56042=>"101111000",
56043=>"000001001",
56044=>"001111111",
56045=>"110001000",
56046=>"111000000",
56047=>"111111000",
56048=>"111101001",
56049=>"100000000",
56050=>"111011011",
56051=>"110000000",
56052=>"000001001",
56053=>"111111111",
56054=>"100000000",
56055=>"000000010",
56056=>"000000000",
56057=>"111110000",
56058=>"000000000",
56059=>"111110100",
56060=>"111000000",
56061=>"110000000",
56062=>"000001000",
56063=>"111111110",
56064=>"001100011",
56065=>"111111101",
56066=>"000110111",
56067=>"100111111",
56068=>"000111011",
56069=>"000000000",
56070=>"011101111",
56071=>"010111011",
56072=>"100111111",
56073=>"111111100",
56074=>"111100000",
56075=>"000000000",
56076=>"000000111",
56077=>"010010000",
56078=>"000001101",
56079=>"111111000",
56080=>"111000000",
56081=>"111111111",
56082=>"001010111",
56083=>"001010001",
56084=>"111100111",
56085=>"000101000",
56086=>"110011011",
56087=>"111111101",
56088=>"101000000",
56089=>"111100100",
56090=>"111111101",
56091=>"000111010",
56092=>"111111000",
56093=>"101111000",
56094=>"000000000",
56095=>"000000111",
56096=>"101000000",
56097=>"010000001",
56098=>"011101101",
56099=>"111111000",
56100=>"111110000",
56101=>"100100100",
56102=>"111001000",
56103=>"110111111",
56104=>"111001101",
56105=>"010000000",
56106=>"110000000",
56107=>"101000110",
56108=>"101110101",
56109=>"001010111",
56110=>"101000110",
56111=>"000000011",
56112=>"111000000",
56113=>"001111110",
56114=>"000101101",
56115=>"000001000",
56116=>"010000000",
56117=>"011010110",
56118=>"111100100",
56119=>"000010110",
56120=>"100001000",
56121=>"000100111",
56122=>"001011111",
56123=>"111000001",
56124=>"000100110",
56125=>"111001000",
56126=>"000000010",
56127=>"111011110",
56128=>"001000111",
56129=>"101101001",
56130=>"111100111",
56131=>"000000011",
56132=>"000001111",
56133=>"000111111",
56134=>"111101111",
56135=>"110000111",
56136=>"100111001",
56137=>"010101000",
56138=>"111010111",
56139=>"111111010",
56140=>"000111111",
56141=>"100011010",
56142=>"100111111",
56143=>"000000011",
56144=>"000100111",
56145=>"111101000",
56146=>"101111101",
56147=>"001001001",
56148=>"000000101",
56149=>"100110010",
56150=>"111100011",
56151=>"111101000",
56152=>"000000011",
56153=>"011111100",
56154=>"000110110",
56155=>"111100000",
56156=>"111001000",
56157=>"001110110",
56158=>"111010011",
56159=>"000001100",
56160=>"111101111",
56161=>"000010111",
56162=>"000101111",
56163=>"000001111",
56164=>"000000010",
56165=>"011111001",
56166=>"010001010",
56167=>"000111101",
56168=>"110100111",
56169=>"011000000",
56170=>"111110101",
56171=>"010000101",
56172=>"110111111",
56173=>"101000000",
56174=>"011100000",
56175=>"001111010",
56176=>"110011011",
56177=>"010000101",
56178=>"111001001",
56179=>"000000111",
56180=>"111110111",
56181=>"101111111",
56182=>"111101000",
56183=>"000000110",
56184=>"000000011",
56185=>"000000000",
56186=>"111111000",
56187=>"000000011",
56188=>"000000001",
56189=>"100001110",
56190=>"111000000",
56191=>"000000001",
56192=>"111000000",
56193=>"000001010",
56194=>"111111010",
56195=>"111001011",
56196=>"101111111",
56197=>"100000000",
56198=>"101101111",
56199=>"001000010",
56200=>"011110110",
56201=>"000111011",
56202=>"011000111",
56203=>"000000101",
56204=>"000000111",
56205=>"001010111",
56206=>"101101010",
56207=>"001001101",
56208=>"011111110",
56209=>"111000000",
56210=>"111010000",
56211=>"000000000",
56212=>"000101000",
56213=>"100001000",
56214=>"000111111",
56215=>"101111000",
56216=>"111000000",
56217=>"011001101",
56218=>"111000000",
56219=>"001000000",
56220=>"000000001",
56221=>"000000111",
56222=>"111001101",
56223=>"000001001",
56224=>"001111000",
56225=>"000000111",
56226=>"001000000",
56227=>"011001101",
56228=>"000010000",
56229=>"101001011",
56230=>"110110110",
56231=>"010101000",
56232=>"111110111",
56233=>"000110001",
56234=>"000000000",
56235=>"111110100",
56236=>"010000110",
56237=>"000000111",
56238=>"110100101",
56239=>"000000101",
56240=>"111000111",
56241=>"001001010",
56242=>"000110111",
56243=>"000001001",
56244=>"000100101",
56245=>"111001000",
56246=>"111100100",
56247=>"000000000",
56248=>"000011010",
56249=>"000001100",
56250=>"101000010",
56251=>"000000001",
56252=>"010001001",
56253=>"000101111",
56254=>"101100010",
56255=>"010000110",
56256=>"000000101",
56257=>"111000000",
56258=>"010100101",
56259=>"001011010",
56260=>"000010111",
56261=>"100110011",
56262=>"111101000",
56263=>"010000000",
56264=>"000101000",
56265=>"111100110",
56266=>"111001000",
56267=>"111110111",
56268=>"000100111",
56269=>"011110000",
56270=>"000101000",
56271=>"110000001",
56272=>"000111111",
56273=>"001110111",
56274=>"100000000",
56275=>"110111001",
56276=>"000000100",
56277=>"100001010",
56278=>"000011111",
56279=>"111111101",
56280=>"001000000",
56281=>"000110001",
56282=>"110110010",
56283=>"010101111",
56284=>"001110110",
56285=>"101100111",
56286=>"111101101",
56287=>"000000101",
56288=>"000100111",
56289=>"000101011",
56290=>"001001001",
56291=>"111011011",
56292=>"000000000",
56293=>"101101111",
56294=>"001111111",
56295=>"111101110",
56296=>"000011001",
56297=>"010010000",
56298=>"011011100",
56299=>"110001000",
56300=>"111111100",
56301=>"100010000",
56302=>"010000000",
56303=>"101000000",
56304=>"100000000",
56305=>"011011111",
56306=>"000010101",
56307=>"100011111",
56308=>"111011111",
56309=>"001101000",
56310=>"000000000",
56311=>"011101111",
56312=>"111000000",
56313=>"111000001",
56314=>"111000010",
56315=>"000110111",
56316=>"110110010",
56317=>"001000100",
56318=>"001110110",
56319=>"001110011",
56320=>"111011100",
56321=>"000100111",
56322=>"100000100",
56323=>"000000010",
56324=>"000011011",
56325=>"111000111",
56326=>"011011010",
56327=>"000110111",
56328=>"010010000",
56329=>"010111000",
56330=>"110011111",
56331=>"000000110",
56332=>"100100101",
56333=>"011011010",
56334=>"101011001",
56335=>"000000000",
56336=>"110101111",
56337=>"110011110",
56338=>"000010100",
56339=>"000111111",
56340=>"111011101",
56341=>"010100100",
56342=>"000100011",
56343=>"000010000",
56344=>"000011000",
56345=>"010010000",
56346=>"000100101",
56347=>"111111110",
56348=>"111111000",
56349=>"111011000",
56350=>"101111010",
56351=>"000110100",
56352=>"000000111",
56353=>"000010000",
56354=>"001110101",
56355=>"000101010",
56356=>"000001000",
56357=>"110010000",
56358=>"000100100",
56359=>"000000010",
56360=>"101100111",
56361=>"010011011",
56362=>"111111011",
56363=>"111100100",
56364=>"111111011",
56365=>"001000111",
56366=>"111100111",
56367=>"010011110",
56368=>"001010111",
56369=>"001001001",
56370=>"101001110",
56371=>"011110111",
56372=>"011111010",
56373=>"111111110",
56374=>"111111111",
56375=>"111111110",
56376=>"011111111",
56377=>"000011000",
56378=>"010110111",
56379=>"000111000",
56380=>"100100001",
56381=>"111111001",
56382=>"000000010",
56383=>"101111111",
56384=>"000000000",
56385=>"010000010",
56386=>"101100111",
56387=>"001100110",
56388=>"010011000",
56389=>"000000101",
56390=>"001011000",
56391=>"101001000",
56392=>"000001111",
56393=>"100100111",
56394=>"101100101",
56395=>"100100000",
56396=>"000111010",
56397=>"001101101",
56398=>"100110110",
56399=>"011010010",
56400=>"010011011",
56401=>"000101111",
56402=>"101111000",
56403=>"011000011",
56404=>"111101101",
56405=>"001111011",
56406=>"100110110",
56407=>"001000000",
56408=>"100110111",
56409=>"000001001",
56410=>"001111011",
56411=>"110110100",
56412=>"100000111",
56413=>"001001001",
56414=>"111111000",
56415=>"110100101",
56416=>"000100100",
56417=>"100000101",
56418=>"100100000",
56419=>"110110110",
56420=>"010011001",
56421=>"011011111",
56422=>"111111111",
56423=>"010011000",
56424=>"010010010",
56425=>"000000000",
56426=>"110101100",
56427=>"111000000",
56428=>"000000011",
56429=>"011000000",
56430=>"100100000",
56431=>"111000011",
56432=>"011001001",
56433=>"000000111",
56434=>"111111111",
56435=>"100000000",
56436=>"111000000",
56437=>"100101110",
56438=>"111111111",
56439=>"111000000",
56440=>"000000011",
56441=>"010000000",
56442=>"111101000",
56443=>"010011110",
56444=>"100110001",
56445=>"010000100",
56446=>"111100111",
56447=>"110111111",
56448=>"101000000",
56449=>"111100110",
56450=>"011011010",
56451=>"111011010",
56452=>"011100000",
56453=>"111011010",
56454=>"011001000",
56455=>"100001000",
56456=>"000111110",
56457=>"000000000",
56458=>"000000100",
56459=>"111000100",
56460=>"000000000",
56461=>"000100111",
56462=>"101001001",
56463=>"101000001",
56464=>"111111101",
56465=>"010011101",
56466=>"011010000",
56467=>"000100011",
56468=>"000010011",
56469=>"111000001",
56470=>"101001000",
56471=>"000000001",
56472=>"000010010",
56473=>"000100111",
56474=>"100100100",
56475=>"001100000",
56476=>"000100011",
56477=>"001100000",
56478=>"000000111",
56479=>"101111111",
56480=>"000100000",
56481=>"000000011",
56482=>"110000101",
56483=>"111011010",
56484=>"010010111",
56485=>"000000010",
56486=>"001000011",
56487=>"001011000",
56488=>"111000111",
56489=>"000100000",
56490=>"000000110",
56491=>"111000000",
56492=>"111111001",
56493=>"011111000",
56494=>"110110110",
56495=>"111000111",
56496=>"010000111",
56497=>"001100100",
56498=>"110110000",
56499=>"000110010",
56500=>"101111110",
56501=>"010000000",
56502=>"011000100",
56503=>"111000011",
56504=>"001000100",
56505=>"000110110",
56506=>"111011000",
56507=>"111011010",
56508=>"010000000",
56509=>"110111001",
56510=>"110110100",
56511=>"000000011",
56512=>"000000000",
56513=>"100101100",
56514=>"111000000",
56515=>"001011001",
56516=>"111000001",
56517=>"100111101",
56518=>"000011011",
56519=>"110100100",
56520=>"010100011",
56521=>"000100000",
56522=>"000000000",
56523=>"100100111",
56524=>"010011011",
56525=>"001011010",
56526=>"111111011",
56527=>"101000110",
56528=>"110011010",
56529=>"101000110",
56530=>"000000000",
56531=>"100100101",
56532=>"111101101",
56533=>"000000000",
56534=>"000011011",
56535=>"111010000",
56536=>"100100101",
56537=>"011000100",
56538=>"010000100",
56539=>"101100100",
56540=>"011111111",
56541=>"001010011",
56542=>"100000000",
56543=>"000001111",
56544=>"110000000",
56545=>"101100111",
56546=>"111100100",
56547=>"000000000",
56548=>"000000000",
56549=>"011111000",
56550=>"010000010",
56551=>"010100110",
56552=>"110000111",
56553=>"000000000",
56554=>"111011011",
56555=>"100111000",
56556=>"100100101",
56557=>"101000100",
56558=>"110100000",
56559=>"010101010",
56560=>"000000000",
56561=>"011001110",
56562=>"101100000",
56563=>"011111000",
56564=>"010000011",
56565=>"000011000",
56566=>"000010010",
56567=>"011101100",
56568=>"111100111",
56569=>"000011111",
56570=>"000000000",
56571=>"110100000",
56572=>"000000000",
56573=>"100100000",
56574=>"110110100",
56575=>"100000100",
56576=>"010001000",
56577=>"000101111",
56578=>"111000000",
56579=>"000110110",
56580=>"100110100",
56581=>"101011010",
56582=>"111100000",
56583=>"101010101",
56584=>"010011001",
56585=>"010111010",
56586=>"011111101",
56587=>"000000000",
56588=>"011101101",
56589=>"000000001",
56590=>"000000101",
56591=>"000000000",
56592=>"111111000",
56593=>"101000000",
56594=>"010111010",
56595=>"000111000",
56596=>"111111111",
56597=>"010000100",
56598=>"000000011",
56599=>"111111010",
56600=>"111101001",
56601=>"011000000",
56602=>"100000000",
56603=>"100100101",
56604=>"110000000",
56605=>"111111111",
56606=>"010000000",
56607=>"000000000",
56608=>"111100000",
56609=>"000000101",
56610=>"000000000",
56611=>"000010011",
56612=>"111110110",
56613=>"010010001",
56614=>"000110000",
56615=>"100101001",
56616=>"101001110",
56617=>"111101001",
56618=>"110101100",
56619=>"010111111",
56620=>"111111011",
56621=>"010000101",
56622=>"100010011",
56623=>"010010111",
56624=>"101011000",
56625=>"001010010",
56626=>"111100000",
56627=>"100000101",
56628=>"111000000",
56629=>"010110001",
56630=>"000010011",
56631=>"010110100",
56632=>"101111100",
56633=>"101101111",
56634=>"000010010",
56635=>"111010010",
56636=>"000111001",
56637=>"111111111",
56638=>"100000000",
56639=>"011011011",
56640=>"000000111",
56641=>"000110011",
56642=>"010010100",
56643=>"000111011",
56644=>"110101010",
56645=>"010000000",
56646=>"110010110",
56647=>"111111110",
56648=>"101000000",
56649=>"000010010",
56650=>"111101111",
56651=>"100011011",
56652=>"111100100",
56653=>"111110011",
56654=>"100110001",
56655=>"111111111",
56656=>"111111011",
56657=>"111110111",
56658=>"101010011",
56659=>"110001001",
56660=>"000000000",
56661=>"100100111",
56662=>"101111011",
56663=>"101111000",
56664=>"001000101",
56665=>"001011111",
56666=>"000100100",
56667=>"011011001",
56668=>"000000111",
56669=>"100000000",
56670=>"101000000",
56671=>"001111110",
56672=>"000000001",
56673=>"000011011",
56674=>"000000110",
56675=>"110111001",
56676=>"000100101",
56677=>"110100100",
56678=>"101111111",
56679=>"000111001",
56680=>"110011000",
56681=>"111110111",
56682=>"111111111",
56683=>"100011010",
56684=>"101110111",
56685=>"111000000",
56686=>"000011000",
56687=>"111000000",
56688=>"100111110",
56689=>"100110111",
56690=>"000011011",
56691=>"101000000",
56692=>"111111000",
56693=>"110000000",
56694=>"000000100",
56695=>"111111011",
56696=>"000110000",
56697=>"100100010",
56698=>"111101001",
56699=>"001011111",
56700=>"001110011",
56701=>"100100110",
56702=>"100110000",
56703=>"010011011",
56704=>"001100000",
56705=>"111111111",
56706=>"101011010",
56707=>"000111111",
56708=>"010110101",
56709=>"111111010",
56710=>"000010100",
56711=>"000001000",
56712=>"001011011",
56713=>"101001000",
56714=>"001100000",
56715=>"100000000",
56716=>"111000100",
56717=>"100111001",
56718=>"000010110",
56719=>"100000100",
56720=>"011011001",
56721=>"000001011",
56722=>"011011010",
56723=>"001000010",
56724=>"100001110",
56725=>"011111101",
56726=>"111100100",
56727=>"010110100",
56728=>"111111111",
56729=>"100011010",
56730=>"011111111",
56731=>"111011000",
56732=>"111100000",
56733=>"000000000",
56734=>"110110000",
56735=>"111100101",
56736=>"011011011",
56737=>"011010000",
56738=>"110110000",
56739=>"100000100",
56740=>"100111110",
56741=>"011110110",
56742=>"010000110",
56743=>"000010001",
56744=>"001000000",
56745=>"001100000",
56746=>"101101111",
56747=>"100100101",
56748=>"000000111",
56749=>"000100111",
56750=>"100111000",
56751=>"001111111",
56752=>"100111011",
56753=>"100100000",
56754=>"111010011",
56755=>"000000001",
56756=>"010010111",
56757=>"000000000",
56758=>"011100100",
56759=>"000000000",
56760=>"011111010",
56761=>"001100000",
56762=>"100101111",
56763=>"111001000",
56764=>"001100001",
56765=>"111000000",
56766=>"110110110",
56767=>"000111111",
56768=>"011011010",
56769=>"000111110",
56770=>"011000000",
56771=>"110111101",
56772=>"101100010",
56773=>"111100000",
56774=>"000111111",
56775=>"100000100",
56776=>"001000000",
56777=>"010111010",
56778=>"100000010",
56779=>"000111110",
56780=>"000011000",
56781=>"100100001",
56782=>"011111000",
56783=>"000110111",
56784=>"011111010",
56785=>"011000001",
56786=>"100100000",
56787=>"100111111",
56788=>"110010111",
56789=>"101001000",
56790=>"101100101",
56791=>"000100011",
56792=>"111111111",
56793=>"111011011",
56794=>"110011011",
56795=>"111000100",
56796=>"000000011",
56797=>"001111110",
56798=>"100100110",
56799=>"101101111",
56800=>"010011011",
56801=>"101100001",
56802=>"001111011",
56803=>"000100001",
56804=>"000000000",
56805=>"000000000",
56806=>"111110010",
56807=>"001111101",
56808=>"110111111",
56809=>"101111001",
56810=>"101101010",
56811=>"111000001",
56812=>"111100100",
56813=>"000100011",
56814=>"111001010",
56815=>"010000010",
56816=>"101111000",
56817=>"110100100",
56818=>"001011011",
56819=>"010110110",
56820=>"100001100",
56821=>"000000011",
56822=>"111100010",
56823=>"000011110",
56824=>"110111000",
56825=>"111111100",
56826=>"011011110",
56827=>"110000010",
56828=>"111111111",
56829=>"000110010",
56830=>"001011001",
56831=>"000000101",
56832=>"010000000",
56833=>"000010010",
56834=>"000000001",
56835=>"001001111",
56836=>"000000000",
56837=>"001001101",
56838=>"000000000",
56839=>"101010111",
56840=>"000000000",
56841=>"000000000",
56842=>"111111011",
56843=>"101001101",
56844=>"000000000",
56845=>"101001000",
56846=>"010000001",
56847=>"001111111",
56848=>"000010011",
56849=>"010010010",
56850=>"110110110",
56851=>"000110111",
56852=>"010101111",
56853=>"000011010",
56854=>"111100000",
56855=>"110110010",
56856=>"010000000",
56857=>"011111111",
56858=>"000001111",
56859=>"000000100",
56860=>"000101110",
56861=>"101000010",
56862=>"010011100",
56863=>"000101001",
56864=>"001001111",
56865=>"111100001",
56866=>"011100000",
56867=>"001101111",
56868=>"111101110",
56869=>"001001011",
56870=>"000111010",
56871=>"000000000",
56872=>"010111111",
56873=>"010011011",
56874=>"111110111",
56875=>"011111010",
56876=>"111111111",
56877=>"011001111",
56878=>"111111011",
56879=>"001000000",
56880=>"111101001",
56881=>"100101011",
56882=>"010111110",
56883=>"111111111",
56884=>"011010000",
56885=>"010001000",
56886=>"111110011",
56887=>"000000000",
56888=>"011111111",
56889=>"000000011",
56890=>"000000000",
56891=>"110000111",
56892=>"111100111",
56893=>"111111010",
56894=>"000000001",
56895=>"001000100",
56896=>"111111111",
56897=>"110010010",
56898=>"111111111",
56899=>"000000000",
56900=>"110111111",
56901=>"000000000",
56902=>"000001101",
56903=>"110110111",
56904=>"000100011",
56905=>"101000101",
56906=>"111111111",
56907=>"100110010",
56908=>"101000000",
56909=>"111011011",
56910=>"111101110",
56911=>"010111111",
56912=>"000001000",
56913=>"111010000",
56914=>"101101111",
56915=>"011000000",
56916=>"000000000",
56917=>"000000100",
56918=>"001001000",
56919=>"000010110",
56920=>"000000000",
56921=>"000100111",
56922=>"100100000",
56923=>"001011001",
56924=>"111001101",
56925=>"100100101",
56926=>"010110111",
56927=>"000000001",
56928=>"111000000",
56929=>"001000101",
56930=>"000000001",
56931=>"111111101",
56932=>"101101000",
56933=>"101000000",
56934=>"111101010",
56935=>"000110011",
56936=>"111001000",
56937=>"111111111",
56938=>"000000000",
56939=>"010111001",
56940=>"111110111",
56941=>"010110111",
56942=>"000000000",
56943=>"000100010",
56944=>"100100000",
56945=>"110111010",
56946=>"111010110",
56947=>"000110010",
56948=>"000000111",
56949=>"000101101",
56950=>"011011110",
56951=>"000000001",
56952=>"010011101",
56953=>"000001111",
56954=>"111000010",
56955=>"111101100",
56956=>"111000011",
56957=>"111001101",
56958=>"110000000",
56959=>"000000000",
56960=>"111000000",
56961=>"000110110",
56962=>"010001011",
56963=>"101101100",
56964=>"010000101",
56965=>"101000000",
56966=>"010111010",
56967=>"110001111",
56968=>"011011111",
56969=>"111101000",
56970=>"000000000",
56971=>"010110111",
56972=>"000000000",
56973=>"000101111",
56974=>"010000000",
56975=>"000110100",
56976=>"011011011",
56977=>"000000001",
56978=>"000000010",
56979=>"111001111",
56980=>"100100010",
56981=>"000000111",
56982=>"010110010",
56983=>"100111111",
56984=>"101001000",
56985=>"110110101",
56986=>"000111010",
56987=>"001000000",
56988=>"100100000",
56989=>"101001000",
56990=>"000111110",
56991=>"100000000",
56992=>"010000010",
56993=>"101000111",
56994=>"000111111",
56995=>"111110100",
56996=>"011000000",
56997=>"100110110",
56998=>"000010101",
56999=>"111111111",
57000=>"010000110",
57001=>"111110111",
57002=>"001000000",
57003=>"000000000",
57004=>"110001000",
57005=>"000001011",
57006=>"000001001",
57007=>"111111111",
57008=>"000000010",
57009=>"010110100",
57010=>"000000000",
57011=>"001100100",
57012=>"001111111",
57013=>"111101101",
57014=>"000011111",
57015=>"010111111",
57016=>"110101111",
57017=>"111101011",
57018=>"101001001",
57019=>"110111010",
57020=>"110111111",
57021=>"000010000",
57022=>"000000001",
57023=>"000001101",
57024=>"010110000",
57025=>"000000000",
57026=>"101010010",
57027=>"111100100",
57028=>"100110011",
57029=>"010001010",
57030=>"110000101",
57031=>"101000100",
57032=>"111101111",
57033=>"110111100",
57034=>"010111000",
57035=>"011001000",
57036=>"111010010",
57037=>"111100100",
57038=>"000000100",
57039=>"111100001",
57040=>"000000111",
57041=>"111100110",
57042=>"000111100",
57043=>"000001111",
57044=>"000000000",
57045=>"000010010",
57046=>"000000000",
57047=>"000000010",
57048=>"011111111",
57049=>"010111101",
57050=>"111000111",
57051=>"001001000",
57052=>"100011011",
57053=>"101110111",
57054=>"001111111",
57055=>"000000110",
57056=>"111000101",
57057=>"001011111",
57058=>"000010010",
57059=>"101110110",
57060=>"000000000",
57061=>"001000000",
57062=>"111001111",
57063=>"011000100",
57064=>"011001111",
57065=>"000101111",
57066=>"111110110",
57067=>"000110000",
57068=>"100101101",
57069=>"000111111",
57070=>"000110110",
57071=>"101001110",
57072=>"111101111",
57073=>"001110101",
57074=>"000000000",
57075=>"001000011",
57076=>"111100011",
57077=>"001111000",
57078=>"001101010",
57079=>"111111111",
57080=>"000010111",
57081=>"000111111",
57082=>"010111111",
57083=>"111111001",
57084=>"000010000",
57085=>"001001101",
57086=>"000100100",
57087=>"001011001",
57088=>"101000110",
57089=>"000010111",
57090=>"000011010",
57091=>"111010111",
57092=>"001001000",
57093=>"110110111",
57094=>"101101001",
57095=>"111010111",
57096=>"001101101",
57097=>"011000000",
57098=>"100000000",
57099=>"000000010",
57100=>"000011000",
57101=>"010110000",
57102=>"100011100",
57103=>"111110101",
57104=>"011100000",
57105=>"010010010",
57106=>"100100110",
57107=>"100110001",
57108=>"100011000",
57109=>"000010111",
57110=>"110111111",
57111=>"110100111",
57112=>"010110000",
57113=>"101111111",
57114=>"111011101",
57115=>"111000111",
57116=>"111111111",
57117=>"110000011",
57118=>"111010011",
57119=>"101101111",
57120=>"101111100",
57121=>"000000111",
57122=>"000000001",
57123=>"111111000",
57124=>"000101101",
57125=>"100000011",
57126=>"111111101",
57127=>"111111100",
57128=>"001111111",
57129=>"000010001",
57130=>"010000000",
57131=>"100111111",
57132=>"001001101",
57133=>"000000001",
57134=>"111111000",
57135=>"000100000",
57136=>"000000011",
57137=>"000001000",
57138=>"000010111",
57139=>"111000010",
57140=>"101011010",
57141=>"000000000",
57142=>"000000100",
57143=>"011001000",
57144=>"110010100",
57145=>"000000000",
57146=>"111101111",
57147=>"101011000",
57148=>"101111011",
57149=>"101111101",
57150=>"000000000",
57151=>"011000000",
57152=>"001000111",
57153=>"010110100",
57154=>"010111101",
57155=>"010011001",
57156=>"110000010",
57157=>"000000011",
57158=>"010111000",
57159=>"111111000",
57160=>"000000111",
57161=>"111110000",
57162=>"000100000",
57163=>"111101010",
57164=>"100100101",
57165=>"010101100",
57166=>"100100001",
57167=>"101111000",
57168=>"000111101",
57169=>"000000000",
57170=>"110011010",
57171=>"101001001",
57172=>"000010110",
57173=>"001000101",
57174=>"100001000",
57175=>"011010010",
57176=>"011001001",
57177=>"111001000",
57178=>"000110101",
57179=>"010100000",
57180=>"110010000",
57181=>"001001101",
57182=>"110000111",
57183=>"001000100",
57184=>"001111111",
57185=>"111101110",
57186=>"110100100",
57187=>"100101101",
57188=>"111101000",
57189=>"111101101",
57190=>"110111100",
57191=>"110111000",
57192=>"101000111",
57193=>"111010010",
57194=>"111010110",
57195=>"101111111",
57196=>"001010000",
57197=>"111000000",
57198=>"110100000",
57199=>"001000010",
57200=>"100001000",
57201=>"111010000",
57202=>"000000011",
57203=>"111111011",
57204=>"111010110",
57205=>"000100011",
57206=>"010111111",
57207=>"000110000",
57208=>"110111010",
57209=>"111000011",
57210=>"000000111",
57211=>"111001000",
57212=>"000000011",
57213=>"111100000",
57214=>"111111111",
57215=>"101101101",
57216=>"000010000",
57217=>"100000111",
57218=>"111111000",
57219=>"101001000",
57220=>"111000000",
57221=>"111111110",
57222=>"001001000",
57223=>"101100100",
57224=>"000100000",
57225=>"111111111",
57226=>"111111100",
57227=>"101111010",
57228=>"000101101",
57229=>"110110111",
57230=>"010000100",
57231=>"011011110",
57232=>"001101001",
57233=>"000011111",
57234=>"111000000",
57235=>"011010010",
57236=>"011001100",
57237=>"111010000",
57238=>"111101111",
57239=>"100100100",
57240=>"111000000",
57241=>"000111111",
57242=>"100000100",
57243=>"000000111",
57244=>"000010111",
57245=>"111011111",
57246=>"111010011",
57247=>"001000000",
57248=>"000000001",
57249=>"011000111",
57250=>"011000000",
57251=>"100000111",
57252=>"111110000",
57253=>"100100000",
57254=>"001111000",
57255=>"010011101",
57256=>"111010000",
57257=>"000111111",
57258=>"000100011",
57259=>"010000000",
57260=>"011110011",
57261=>"111111000",
57262=>"110000110",
57263=>"111111000",
57264=>"111000001",
57265=>"000001001",
57266=>"000100111",
57267=>"000000011",
57268=>"110111101",
57269=>"000010101",
57270=>"001000000",
57271=>"000000101",
57272=>"101111110",
57273=>"110111001",
57274=>"111000010",
57275=>"111010001",
57276=>"000011011",
57277=>"000111111",
57278=>"111111001",
57279=>"000010000",
57280=>"000000010",
57281=>"000000000",
57282=>"111111111",
57283=>"000101001",
57284=>"010010111",
57285=>"110110110",
57286=>"000011000",
57287=>"111001111",
57288=>"100000101",
57289=>"000001101",
57290=>"001110000",
57291=>"010110110",
57292=>"111100000",
57293=>"000110110",
57294=>"000011111",
57295=>"001110111",
57296=>"000111000",
57297=>"100100111",
57298=>"101101010",
57299=>"111011011",
57300=>"100111111",
57301=>"100100111",
57302=>"000000101",
57303=>"111000111",
57304=>"001010010",
57305=>"101000010",
57306=>"000100000",
57307=>"111100101",
57308=>"000110110",
57309=>"100111111",
57310=>"000000010",
57311=>"111010000",
57312=>"000101000",
57313=>"010111111",
57314=>"111101000",
57315=>"111101001",
57316=>"111111011",
57317=>"000000101",
57318=>"000011111",
57319=>"011001000",
57320=>"111010111",
57321=>"101111111",
57322=>"011001011",
57323=>"000111111",
57324=>"000000001",
57325=>"000000000",
57326=>"000000000",
57327=>"101101100",
57328=>"100000010",
57329=>"011011001",
57330=>"110111100",
57331=>"111101001",
57332=>"101100000",
57333=>"100101111",
57334=>"000010111",
57335=>"101111111",
57336=>"000000110",
57337=>"000000010",
57338=>"101111111",
57339=>"101111011",
57340=>"111101100",
57341=>"000000000",
57342=>"011000000",
57343=>"111111000",
57344=>"100101011",
57345=>"001000100",
57346=>"000000111",
57347=>"000110110",
57348=>"001000000",
57349=>"111101001",
57350=>"011000000",
57351=>"111111101",
57352=>"001101111",
57353=>"000001101",
57354=>"000000011",
57355=>"010000111",
57356=>"111111010",
57357=>"001111111",
57358=>"000000000",
57359=>"011111111",
57360=>"001101101",
57361=>"000000000",
57362=>"111110111",
57363=>"010000000",
57364=>"101100110",
57365=>"000000101",
57366=>"000000000",
57367=>"011111111",
57368=>"111100111",
57369=>"111111111",
57370=>"101101111",
57371=>"010000100",
57372=>"111000010",
57373=>"001011000",
57374=>"000100100",
57375=>"000000001",
57376=>"111011111",
57377=>"001110111",
57378=>"001011111",
57379=>"001000000",
57380=>"000010000",
57381=>"001001111",
57382=>"100000001",
57383=>"000110111",
57384=>"011010111",
57385=>"010111111",
57386=>"001111000",
57387=>"000000100",
57388=>"001011110",
57389=>"011010111",
57390=>"111101101",
57391=>"011010000",
57392=>"001111110",
57393=>"111101100",
57394=>"000000000",
57395=>"000001100",
57396=>"001000101",
57397=>"000000000",
57398=>"000000000",
57399=>"000100101",
57400=>"111000000",
57401=>"000101101",
57402=>"111010111",
57403=>"000000000",
57404=>"011001011",
57405=>"011011111",
57406=>"000000101",
57407=>"000001001",
57408=>"101111111",
57409=>"011111010",
57410=>"101111111",
57411=>"001000001",
57412=>"000010000",
57413=>"101111010",
57414=>"010101100",
57415=>"001001110",
57416=>"111011111",
57417=>"111111111",
57418=>"000010111",
57419=>"101101101",
57420=>"111111111",
57421=>"000000110",
57422=>"110100010",
57423=>"000000110",
57424=>"000000000",
57425=>"110111110",
57426=>"000000111",
57427=>"111110001",
57428=>"001000001",
57429=>"101101101",
57430=>"010010000",
57431=>"000010111",
57432=>"001101000",
57433=>"111111111",
57434=>"000000000",
57435=>"000100100",
57436=>"000000011",
57437=>"100110000",
57438=>"111111111",
57439=>"101000000",
57440=>"100110111",
57441=>"010000000",
57442=>"111111111",
57443=>"001010000",
57444=>"001000011",
57445=>"010111000",
57446=>"111111100",
57447=>"001101001",
57448=>"000000010",
57449=>"111000001",
57450=>"111001101",
57451=>"111111010",
57452=>"011111001",
57453=>"011000000",
57454=>"010111000",
57455=>"001110111",
57456=>"111100111",
57457=>"101110111",
57458=>"000000001",
57459=>"111111011",
57460=>"111101000",
57461=>"101101000",
57462=>"100000001",
57463=>"001111100",
57464=>"000000000",
57465=>"111001100",
57466=>"000001101",
57467=>"111111110",
57468=>"001001001",
57469=>"111011010",
57470=>"111111111",
57471=>"000100111",
57472=>"001000000",
57473=>"000100000",
57474=>"000111000",
57475=>"101011000",
57476=>"000101111",
57477=>"010001000",
57478=>"000100010",
57479=>"010100111",
57480=>"111000110",
57481=>"000000001",
57482=>"101001111",
57483=>"111011000",
57484=>"001101111",
57485=>"000000100",
57486=>"011111111",
57487=>"000000000",
57488=>"110100010",
57489=>"100001000",
57490=>"110101001",
57491=>"011001101",
57492=>"110100000",
57493=>"000000000",
57494=>"111111110",
57495=>"100111011",
57496=>"101101010",
57497=>"000000001",
57498=>"111111111",
57499=>"000010011",
57500=>"010101000",
57501=>"010111111",
57502=>"000001111",
57503=>"010111001",
57504=>"011110111",
57505=>"000000001",
57506=>"111111111",
57507=>"100111101",
57508=>"000100101",
57509=>"000000100",
57510=>"111110110",
57511=>"111101000",
57512=>"000000000",
57513=>"000000001",
57514=>"111110000",
57515=>"000000000",
57516=>"010111110",
57517=>"000000111",
57518=>"000000000",
57519=>"111111111",
57520=>"000101111",
57521=>"100101001",
57522=>"111000100",
57523=>"111111011",
57524=>"111011011",
57525=>"111110000",
57526=>"010111110",
57527=>"111101101",
57528=>"100100111",
57529=>"110101111",
57530=>"101000001",
57531=>"111111111",
57532=>"111000011",
57533=>"111111110",
57534=>"000101100",
57535=>"000111111",
57536=>"000000111",
57537=>"010000000",
57538=>"001011010",
57539=>"011000001",
57540=>"111111111",
57541=>"001001001",
57542=>"000101000",
57543=>"000100100",
57544=>"010111111",
57545=>"000001000",
57546=>"000000101",
57547=>"100111111",
57548=>"000101101",
57549=>"110000100",
57550=>"101101001",
57551=>"101111111",
57552=>"000000000",
57553=>"111111000",
57554=>"111111111",
57555=>"111111111",
57556=>"000000000",
57557=>"001001111",
57558=>"000111110",
57559=>"101011000",
57560=>"111111001",
57561=>"111111111",
57562=>"011011010",
57563=>"000010011",
57564=>"000000001",
57565=>"010110101",
57566=>"111111010",
57567=>"001101111",
57568=>"100000001",
57569=>"001011111",
57570=>"111011011",
57571=>"011001001",
57572=>"000000001",
57573=>"111111101",
57574=>"111101001",
57575=>"000001001",
57576=>"000000100",
57577=>"111101111",
57578=>"000000001",
57579=>"010010111",
57580=>"111111010",
57581=>"000101111",
57582=>"111111111",
57583=>"000010100",
57584=>"110000111",
57585=>"000000000",
57586=>"110111111",
57587=>"000110111",
57588=>"101101111",
57589=>"000000000",
57590=>"101000110",
57591=>"110111011",
57592=>"000100100",
57593=>"000001100",
57594=>"000110000",
57595=>"001001001",
57596=>"000000011",
57597=>"100011001",
57598=>"010100111",
57599=>"000000010",
57600=>"000101111",
57601=>"000000100",
57602=>"010010010",
57603=>"000001111",
57604=>"100000000",
57605=>"000001111",
57606=>"111111100",
57607=>"101101000",
57608=>"110101101",
57609=>"101101101",
57610=>"100000000",
57611=>"000101111",
57612=>"000001101",
57613=>"101100101",
57614=>"000000110",
57615=>"101111110",
57616=>"011000101",
57617=>"111111010",
57618=>"111111110",
57619=>"000100000",
57620=>"111000000",
57621=>"111000000",
57622=>"100000000",
57623=>"000010111",
57624=>"010010000",
57625=>"111111010",
57626=>"011000101",
57627=>"111000101",
57628=>"111111111",
57629=>"000000001",
57630=>"000101001",
57631=>"101000010",
57632=>"000011111",
57633=>"011000010",
57634=>"111010010",
57635=>"111000000",
57636=>"011000001",
57637=>"000011011",
57638=>"010010011",
57639=>"001000101",
57640=>"111010000",
57641=>"110111101",
57642=>"001001111",
57643=>"001000000",
57644=>"010100111",
57645=>"110010000",
57646=>"000101101",
57647=>"001000011",
57648=>"011111110",
57649=>"101110110",
57650=>"111111110",
57651=>"110000111",
57652=>"000010000",
57653=>"000001010",
57654=>"111001000",
57655=>"111111111",
57656=>"000101000",
57657=>"101000100",
57658=>"110000010",
57659=>"111111101",
57660=>"001001011",
57661=>"111111011",
57662=>"000000000",
57663=>"000001001",
57664=>"101001000",
57665=>"000101110",
57666=>"100001111",
57667=>"000100100",
57668=>"110000010",
57669=>"101100000",
57670=>"111111111",
57671=>"101011000",
57672=>"000000010",
57673=>"000001101",
57674=>"000010000",
57675=>"101101100",
57676=>"111111111",
57677=>"111011000",
57678=>"110000001",
57679=>"010111001",
57680=>"000000010",
57681=>"111000000",
57682=>"000101111",
57683=>"111110110",
57684=>"010000100",
57685=>"001000000",
57686=>"000101110",
57687=>"111001101",
57688=>"111000010",
57689=>"000000100",
57690=>"001101101",
57691=>"111000101",
57692=>"000001000",
57693=>"000000100",
57694=>"111111011",
57695=>"000001000",
57696=>"111111111",
57697=>"000000010",
57698=>"000000010",
57699=>"000111101",
57700=>"001000111",
57701=>"000101000",
57702=>"000101111",
57703=>"100100111",
57704=>"111000110",
57705=>"000000000",
57706=>"111000011",
57707=>"000111111",
57708=>"001011111",
57709=>"111000110",
57710=>"000000100",
57711=>"101111111",
57712=>"000011011",
57713=>"001000000",
57714=>"111001000",
57715=>"101111111",
57716=>"100001000",
57717=>"000000001",
57718=>"000000101",
57719=>"110111111",
57720=>"011110100",
57721=>"111101010",
57722=>"011000110",
57723=>"000000010",
57724=>"011001001",
57725=>"001011011",
57726=>"111001111",
57727=>"100000111",
57728=>"111101101",
57729=>"111011111",
57730=>"101111101",
57731=>"000010000",
57732=>"111000000",
57733=>"001111111",
57734=>"100100111",
57735=>"110110110",
57736=>"010110000",
57737=>"101000010",
57738=>"100010011",
57739=>"111111110",
57740=>"000001000",
57741=>"000000110",
57742=>"001001101",
57743=>"000000000",
57744=>"110101100",
57745=>"000111111",
57746=>"111000101",
57747=>"000000001",
57748=>"101010011",
57749=>"000000101",
57750=>"000000111",
57751=>"111101111",
57752=>"011111111",
57753=>"001000101",
57754=>"010000110",
57755=>"001000001",
57756=>"110001011",
57757=>"111001000",
57758=>"111001000",
57759=>"111001110",
57760=>"100100100",
57761=>"010110100",
57762=>"001100111",
57763=>"110010000",
57764=>"001001101",
57765=>"011011111",
57766=>"111110101",
57767=>"000101101",
57768=>"111111000",
57769=>"000000000",
57770=>"000111100",
57771=>"110111111",
57772=>"111110111",
57773=>"100000000",
57774=>"000001011",
57775=>"111111110",
57776=>"011111101",
57777=>"011001011",
57778=>"101011111",
57779=>"000000000",
57780=>"001111100",
57781=>"001010111",
57782=>"111111011",
57783=>"111001111",
57784=>"100100100",
57785=>"011000000",
57786=>"000111111",
57787=>"100101000",
57788=>"100100010",
57789=>"000000010",
57790=>"000100100",
57791=>"000100101",
57792=>"111010110",
57793=>"111110111",
57794=>"011111111",
57795=>"100100100",
57796=>"000001111",
57797=>"001000100",
57798=>"000100100",
57799=>"101000010",
57800=>"111101001",
57801=>"111110110",
57802=>"111011001",
57803=>"111010111",
57804=>"000000100",
57805=>"110100000",
57806=>"000000000",
57807=>"110001111",
57808=>"110110110",
57809=>"001011011",
57810=>"111101000",
57811=>"001110110",
57812=>"001111101",
57813=>"111100000",
57814=>"000100110",
57815=>"000001000",
57816=>"001001000",
57817=>"000000010",
57818=>"110010011",
57819=>"111110000",
57820=>"000000001",
57821=>"000111111",
57822=>"111001110",
57823=>"110000101",
57824=>"010010010",
57825=>"010000011",
57826=>"111000101",
57827=>"001010011",
57828=>"111110101",
57829=>"100101000",
57830=>"101001101",
57831=>"000000101",
57832=>"000100100",
57833=>"000000000",
57834=>"001001000",
57835=>"000100000",
57836=>"010110111",
57837=>"111000100",
57838=>"101100100",
57839=>"111000000",
57840=>"111101111",
57841=>"110110001",
57842=>"000101111",
57843=>"000011011",
57844=>"011011101",
57845=>"111111001",
57846=>"101111111",
57847=>"111111100",
57848=>"111010000",
57849=>"000000000",
57850=>"111110110",
57851=>"011010000",
57852=>"001001000",
57853=>"000111111",
57854=>"111100111",
57855=>"010011011",
57856=>"000010000",
57857=>"000000000",
57858=>"100000101",
57859=>"000000111",
57860=>"111101101",
57861=>"000000100",
57862=>"001000000",
57863=>"000101011",
57864=>"111011011",
57865=>"000000011",
57866=>"011001111",
57867=>"101000111",
57868=>"000101111",
57869=>"000000000",
57870=>"010111000",
57871=>"111111011",
57872=>"010000001",
57873=>"111111110",
57874=>"110000000",
57875=>"000111111",
57876=>"010111111",
57877=>"000001000",
57878=>"001111000",
57879=>"111111000",
57880=>"000000010",
57881=>"000000111",
57882=>"001000000",
57883=>"110110100",
57884=>"010101011",
57885=>"111001101",
57886=>"111100000",
57887=>"011000110",
57888=>"111111000",
57889=>"011001010",
57890=>"001111111",
57891=>"000000000",
57892=>"000111110",
57893=>"111001000",
57894=>"101000100",
57895=>"011001001",
57896=>"001001111",
57897=>"111101000",
57898=>"010000000",
57899=>"010110110",
57900=>"000100110",
57901=>"000000010",
57902=>"111000111",
57903=>"100111110",
57904=>"110001000",
57905=>"110110100",
57906=>"111111000",
57907=>"011111111",
57908=>"110110111",
57909=>"111111111",
57910=>"011111111",
57911=>"011110000",
57912=>"000011111",
57913=>"110000100",
57914=>"000000100",
57915=>"000111110",
57916=>"001001111",
57917=>"000111111",
57918=>"010000000",
57919=>"001000000",
57920=>"000111111",
57921=>"110110000",
57922=>"011111010",
57923=>"010100000",
57924=>"111111111",
57925=>"000010010",
57926=>"011001010",
57927=>"111000100",
57928=>"000000001",
57929=>"000000001",
57930=>"100111000",
57931=>"010001000",
57932=>"001000111",
57933=>"011011011",
57934=>"011011001",
57935=>"101000001",
57936=>"001010111",
57937=>"110111111",
57938=>"111100000",
57939=>"001110100",
57940=>"000101111",
57941=>"001111101",
57942=>"000110100",
57943=>"000001000",
57944=>"000000111",
57945=>"110110000",
57946=>"000000011",
57947=>"011110111",
57948=>"001001000",
57949=>"000101111",
57950=>"011000100",
57951=>"110000101",
57952=>"111001001",
57953=>"000000110",
57954=>"111111111",
57955=>"000000110",
57956=>"000011010",
57957=>"000011000",
57958=>"011001000",
57959=>"001101111",
57960=>"000000100",
57961=>"111111000",
57962=>"000000101",
57963=>"111100111",
57964=>"111001001",
57965=>"110000000",
57966=>"000010000",
57967=>"111111111",
57968=>"001001000",
57969=>"110111000",
57970=>"110111111",
57971=>"111110011",
57972=>"111001111",
57973=>"000110110",
57974=>"000001000",
57975=>"000100100",
57976=>"010000000",
57977=>"000000000",
57978=>"000010011",
57979=>"001111111",
57980=>"110011001",
57981=>"000001001",
57982=>"010011000",
57983=>"000000000",
57984=>"000111000",
57985=>"000010110",
57986=>"000111111",
57987=>"001011101",
57988=>"111000000",
57989=>"000001111",
57990=>"110010000",
57991=>"100100100",
57992=>"100100110",
57993=>"011000100",
57994=>"001000000",
57995=>"111111111",
57996=>"000000000",
57997=>"000000000",
57998=>"111000000",
57999=>"000001000",
58000=>"100100110",
58001=>"000001101",
58002=>"000001000",
58003=>"000000001",
58004=>"001010000",
58005=>"000101001",
58006=>"111111000",
58007=>"010110110",
58008=>"000001010",
58009=>"000000101",
58010=>"101000101",
58011=>"111111111",
58012=>"011011000",
58013=>"111111111",
58014=>"111000000",
58015=>"010000010",
58016=>"000001001",
58017=>"110111100",
58018=>"000000000",
58019=>"001001111",
58020=>"000011111",
58021=>"001011110",
58022=>"000000000",
58023=>"100000011",
58024=>"000010000",
58025=>"000001000",
58026=>"111000001",
58027=>"100010000",
58028=>"111000010",
58029=>"101101111",
58030=>"011101101",
58031=>"111000000",
58032=>"001000111",
58033=>"000000110",
58034=>"000000000",
58035=>"011011011",
58036=>"110111111",
58037=>"111111101",
58038=>"000101111",
58039=>"001000111",
58040=>"100100110",
58041=>"001001001",
58042=>"000000110",
58043=>"111101000",
58044=>"100111110",
58045=>"001001111",
58046=>"110110000",
58047=>"111111000",
58048=>"000000111",
58049=>"010111010",
58050=>"110001111",
58051=>"011011001",
58052=>"011000000",
58053=>"111100100",
58054=>"111010111",
58055=>"111010000",
58056=>"001000111",
58057=>"110110010",
58058=>"100101110",
58059=>"000001111",
58060=>"000100100",
58061=>"000100100",
58062=>"111111001",
58063=>"000011100",
58064=>"111111111",
58065=>"110011011",
58066=>"001000100",
58067=>"000001001",
58068=>"000000001",
58069=>"011000001",
58070=>"000000010",
58071=>"111110000",
58072=>"000000000",
58073=>"101110000",
58074=>"000100111",
58075=>"111111000",
58076=>"010111010",
58077=>"111101000",
58078=>"010111011",
58079=>"000001111",
58080=>"010000000",
58081=>"011000001",
58082=>"111000100",
58083=>"011011000",
58084=>"111001000",
58085=>"110001111",
58086=>"111000100",
58087=>"110111011",
58088=>"111101001",
58089=>"100000000",
58090=>"110100100",
58091=>"000100000",
58092=>"100101100",
58093=>"111000001",
58094=>"010111010",
58095=>"111000101",
58096=>"101001001",
58097=>"111010000",
58098=>"001100000",
58099=>"000011010",
58100=>"000000000",
58101=>"100000010",
58102=>"000000000",
58103=>"010111000",
58104=>"111111000",
58105=>"100000111",
58106=>"000111010",
58107=>"111110000",
58108=>"111100000",
58109=>"001000000",
58110=>"100110010",
58111=>"000110000",
58112=>"110011001",
58113=>"001000000",
58114=>"111000000",
58115=>"100000000",
58116=>"010000000",
58117=>"111101101",
58118=>"111101010",
58119=>"000000111",
58120=>"001111111",
58121=>"000000001",
58122=>"110100001",
58123=>"010100000",
58124=>"100000000",
58125=>"100101010",
58126=>"111100000",
58127=>"101001000",
58128=>"000000011",
58129=>"011000111",
58130=>"011000000",
58131=>"000001000",
58132=>"111111001",
58133=>"111110000",
58134=>"110111000",
58135=>"111001111",
58136=>"111000000",
58137=>"001001010",
58138=>"010110101",
58139=>"110000000",
58140=>"000000000",
58141=>"111000100",
58142=>"111110100",
58143=>"000100110",
58144=>"001001000",
58145=>"011111111",
58146=>"110001000",
58147=>"000111010",
58148=>"001001100",
58149=>"110100000",
58150=>"010111111",
58151=>"111001101",
58152=>"101000110",
58153=>"010110000",
58154=>"001011011",
58155=>"010000000",
58156=>"001110101",
58157=>"100100010",
58158=>"111101101",
58159=>"110001000",
58160=>"000001111",
58161=>"010101110",
58162=>"000001111",
58163=>"110111111",
58164=>"001000000",
58165=>"001011000",
58166=>"011110010",
58167=>"000011000",
58168=>"110011111",
58169=>"001000000",
58170=>"111000100",
58171=>"000000010",
58172=>"001000111",
58173=>"011111111",
58174=>"000000100",
58175=>"000100011",
58176=>"000000000",
58177=>"110101111",
58178=>"101110110",
58179=>"001011001",
58180=>"000111110",
58181=>"000000000",
58182=>"110000000",
58183=>"101001010",
58184=>"100100110",
58185=>"000001000",
58186=>"000000000",
58187=>"000000011",
58188=>"111111000",
58189=>"100101001",
58190=>"000101011",
58191=>"001000101",
58192=>"001110111",
58193=>"111011111",
58194=>"101000010",
58195=>"111001000",
58196=>"111110000",
58197=>"001000110",
58198=>"100000000",
58199=>"110000000",
58200=>"111100100",
58201=>"110100100",
58202=>"000000001",
58203=>"100110011",
58204=>"000111111",
58205=>"000001001",
58206=>"111111011",
58207=>"110100000",
58208=>"000111111",
58209=>"010000101",
58210=>"001011010",
58211=>"011011001",
58212=>"000101000",
58213=>"100100100",
58214=>"011011101",
58215=>"101000000",
58216=>"100110000",
58217=>"111101000",
58218=>"100000110",
58219=>"101010111",
58220=>"010111111",
58221=>"111000111",
58222=>"111111101",
58223=>"111101111",
58224=>"011001000",
58225=>"111110111",
58226=>"010010000",
58227=>"000000011",
58228=>"111001000",
58229=>"000000101",
58230=>"100000000",
58231=>"000110011",
58232=>"000010110",
58233=>"111111101",
58234=>"111111010",
58235=>"000000010",
58236=>"110000011",
58237=>"110100000",
58238=>"000111011",
58239=>"001001000",
58240=>"000010000",
58241=>"010001100",
58242=>"100110111",
58243=>"011000111",
58244=>"111001000",
58245=>"000001011",
58246=>"011001000",
58247=>"000000100",
58248=>"110101001",
58249=>"110000000",
58250=>"000000101",
58251=>"000000010",
58252=>"101000010",
58253=>"111111100",
58254=>"110000111",
58255=>"000000000",
58256=>"010011100",
58257=>"011000100",
58258=>"001001000",
58259=>"111001111",
58260=>"011010000",
58261=>"111000000",
58262=>"100111111",
58263=>"000011101",
58264=>"111111111",
58265=>"100010101",
58266=>"101101111",
58267=>"000101101",
58268=>"000111111",
58269=>"000110110",
58270=>"010100010",
58271=>"010011000",
58272=>"100000011",
58273=>"110110111",
58274=>"111000111",
58275=>"111001001",
58276=>"010010000",
58277=>"000001001",
58278=>"111110000",
58279=>"001011111",
58280=>"111111111",
58281=>"000110110",
58282=>"001000000",
58283=>"010001000",
58284=>"001000000",
58285=>"000000000",
58286=>"110100110",
58287=>"000111100",
58288=>"001000000",
58289=>"000011111",
58290=>"000000000",
58291=>"001001111",
58292=>"011000001",
58293=>"000111000",
58294=>"000111111",
58295=>"000000000",
58296=>"000000111",
58297=>"100110101",
58298=>"000001000",
58299=>"111111001",
58300=>"001101111",
58301=>"111110111",
58302=>"000111001",
58303=>"000011111",
58304=>"100000000",
58305=>"000000010",
58306=>"111111111",
58307=>"011111101",
58308=>"111111100",
58309=>"111110111",
58310=>"111111000",
58311=>"000001111",
58312=>"000111111",
58313=>"000110111",
58314=>"011111111",
58315=>"001000001",
58316=>"111000111",
58317=>"011100100",
58318=>"001011011",
58319=>"000000111",
58320=>"001111101",
58321=>"000100110",
58322=>"110000000",
58323=>"001000000",
58324=>"000101110",
58325=>"010100010",
58326=>"010111111",
58327=>"001001001",
58328=>"101101111",
58329=>"000100000",
58330=>"011110111",
58331=>"111000000",
58332=>"110110100",
58333=>"100010000",
58334=>"000111011",
58335=>"101000000",
58336=>"101000011",
58337=>"111000000",
58338=>"111101001",
58339=>"010110001",
58340=>"110111111",
58341=>"110111001",
58342=>"000111111",
58343=>"100011111",
58344=>"000010111",
58345=>"000000000",
58346=>"000000100",
58347=>"000000111",
58348=>"000010111",
58349=>"000111111",
58350=>"000000000",
58351=>"000110110",
58352=>"000001000",
58353=>"111011111",
58354=>"111111001",
58355=>"111001001",
58356=>"011110101",
58357=>"111011111",
58358=>"000000010",
58359=>"111111111",
58360=>"000000111",
58361=>"101111110",
58362=>"000000010",
58363=>"000111111",
58364=>"001000000",
58365=>"000000000",
58366=>"000111111",
58367=>"111000000",
58368=>"001001000",
58369=>"101100111",
58370=>"110011101",
58371=>"000110011",
58372=>"101101011",
58373=>"110101011",
58374=>"011011011",
58375=>"111100010",
58376=>"000000101",
58377=>"000000010",
58378=>"100100110",
58379=>"000101000",
58380=>"111010001",
58381=>"010111001",
58382=>"011000111",
58383=>"001101110",
58384=>"101111011",
58385=>"000000000",
58386=>"000000100",
58387=>"101010011",
58388=>"000101111",
58389=>"011110000",
58390=>"001001101",
58391=>"001101100",
58392=>"000010000",
58393=>"000111000",
58394=>"011010000",
58395=>"111100111",
58396=>"110111111",
58397=>"010111101",
58398=>"001001101",
58399=>"000000101",
58400=>"111111111",
58401=>"000000000",
58402=>"100101111",
58403=>"000100010",
58404=>"111101101",
58405=>"111100000",
58406=>"010000001",
58407=>"011001001",
58408=>"110011101",
58409=>"000100011",
58410=>"101100111",
58411=>"001111010",
58412=>"111101110",
58413=>"011100011",
58414=>"111000001",
58415=>"011100101",
58416=>"000000111",
58417=>"001001001",
58418=>"011010110",
58419=>"111110000",
58420=>"000101101",
58421=>"010000000",
58422=>"001100110",
58423=>"001001111",
58424=>"010010010",
58425=>"000100101",
58426=>"100010111",
58427=>"011000000",
58428=>"110110110",
58429=>"101101101",
58430=>"000000100",
58431=>"001001000",
58432=>"011000000",
58433=>"101101111",
58434=>"010001001",
58435=>"100001001",
58436=>"000000010",
58437=>"010000000",
58438=>"000110010",
58439=>"000000111",
58440=>"111111011",
58441=>"000101010",
58442=>"101100111",
58443=>"101000001",
58444=>"010010010",
58445=>"101101100",
58446=>"100101101",
58447=>"010111110",
58448=>"000000111",
58449=>"000001101",
58450=>"101111111",
58451=>"000000001",
58452=>"111110111",
58453=>"011111111",
58454=>"011001100",
58455=>"101011000",
58456=>"110010000",
58457=>"100000101",
58458=>"110000010",
58459=>"111100100",
58460=>"010111011",
58461=>"001000001",
58462=>"111111000",
58463=>"001100100",
58464=>"110010011",
58465=>"111111111",
58466=>"011001101",
58467=>"000000110",
58468=>"110000100",
58469=>"000100101",
58470=>"011111110",
58471=>"100001100",
58472=>"000010000",
58473=>"000111000",
58474=>"000000110",
58475=>"000111010",
58476=>"111111111",
58477=>"010010110",
58478=>"100111111",
58479=>"000101111",
58480=>"101101100",
58481=>"010000111",
58482=>"100001001",
58483=>"010000000",
58484=>"101000111",
58485=>"000001000",
58486=>"110000000",
58487=>"111111011",
58488=>"000000001",
58489=>"000000010",
58490=>"000000101",
58491=>"101001000",
58492=>"110010011",
58493=>"100100100",
58494=>"000111101",
58495=>"001000111",
58496=>"101000000",
58497=>"000000011",
58498=>"111111111",
58499=>"001111111",
58500=>"000000111",
58501=>"110000101",
58502=>"001001101",
58503=>"010000000",
58504=>"111001001",
58505=>"111000000",
58506=>"111101111",
58507=>"010000010",
58508=>"111110000",
58509=>"110101001",
58510=>"111111111",
58511=>"000000000",
58512=>"111101001",
58513=>"111001000",
58514=>"100111010",
58515=>"100000000",
58516=>"101011111",
58517=>"000001001",
58518=>"111101001",
58519=>"001000000",
58520=>"000111000",
58521=>"000010000",
58522=>"110111100",
58523=>"100111110",
58524=>"011010110",
58525=>"110101100",
58526=>"000110010",
58527=>"000000101",
58528=>"110110100",
58529=>"000101101",
58530=>"111001000",
58531=>"011100101",
58532=>"010000110",
58533=>"001000100",
58534=>"110110000",
58535=>"110111011",
58536=>"011111101",
58537=>"111011000",
58538=>"101000001",
58539=>"100000011",
58540=>"001111000",
58541=>"011010111",
58542=>"001100110",
58543=>"011000000",
58544=>"110010000",
58545=>"011000000",
58546=>"101100100",
58547=>"100000111",
58548=>"111100000",
58549=>"000000011",
58550=>"000000000",
58551=>"011100000",
58552=>"011011111",
58553=>"110010101",
58554=>"100111010",
58555=>"000000001",
58556=>"111111000",
58557=>"010011000",
58558=>"000101001",
58559=>"010010110",
58560=>"011000000",
58561=>"000000000",
58562=>"001110111",
58563=>"111101100",
58564=>"010110110",
58565=>"001011011",
58566=>"000000111",
58567=>"101100010",
58568=>"011110000",
58569=>"101001000",
58570=>"010110111",
58571=>"011011101",
58572=>"000000001",
58573=>"011011110",
58574=>"000000000",
58575=>"000000111",
58576=>"000100000",
58577=>"101001101",
58578=>"000101111",
58579=>"101001011",
58580=>"111001001",
58581=>"100100110",
58582=>"000111011",
58583=>"101010011",
58584=>"011011000",
58585=>"000110111",
58586=>"011001000",
58587=>"000000000",
58588=>"100100101",
58589=>"010010111",
58590=>"001111101",
58591=>"010010111",
58592=>"001111000",
58593=>"101100101",
58594=>"011110000",
58595=>"111110100",
58596=>"010010100",
58597=>"111101101",
58598=>"011010010",
58599=>"100000111",
58600=>"000010011",
58601=>"000000110",
58602=>"001000001",
58603=>"110101111",
58604=>"000111011",
58605=>"000100000",
58606=>"000000001",
58607=>"101100111",
58608=>"101111011",
58609=>"000110110",
58610=>"010000111",
58611=>"100100100",
58612=>"100000101",
58613=>"001000111",
58614=>"000000000",
58615=>"000111101",
58616=>"001001011",
58617=>"000011110",
58618=>"101101101",
58619=>"101111111",
58620=>"001101111",
58621=>"111011111",
58622=>"111001000",
58623=>"111000111",
58624=>"011011000",
58625=>"010000000",
58626=>"001000001",
58627=>"010000110",
58628=>"000100001",
58629=>"000000000",
58630=>"011111011",
58631=>"100100011",
58632=>"000110010",
58633=>"000000100",
58634=>"000100111",
58635=>"100000000",
58636=>"111000000",
58637=>"010011110",
58638=>"000011111",
58639=>"100000000",
58640=>"000100100",
58641=>"001001011",
58642=>"100001000",
58643=>"110100000",
58644=>"011110010",
58645=>"000101111",
58646=>"110111111",
58647=>"111101101",
58648=>"000000000",
58649=>"111101001",
58650=>"110101000",
58651=>"111001110",
58652=>"111000110",
58653=>"100000000",
58654=>"100100000",
58655=>"000110000",
58656=>"000100011",
58657=>"001011111",
58658=>"000011111",
58659=>"110110111",
58660=>"101101001",
58661=>"000000000",
58662=>"000100010",
58663=>"101000100",
58664=>"001111011",
58665=>"011001111",
58666=>"001001100",
58667=>"110000110",
58668=>"100100111",
58669=>"000100000",
58670=>"111010000",
58671=>"010000111",
58672=>"000000001",
58673=>"110111111",
58674=>"001100100",
58675=>"001001000",
58676=>"010110000",
58677=>"010100000",
58678=>"000100011",
58679=>"100110000",
58680=>"000100110",
58681=>"100010010",
58682=>"000001101",
58683=>"011111111",
58684=>"000000000",
58685=>"010011000",
58686=>"100100100",
58687=>"000110000",
58688=>"111101111",
58689=>"011011001",
58690=>"111011011",
58691=>"110110000",
58692=>"001111011",
58693=>"001100001",
58694=>"111001111",
58695=>"100110111",
58696=>"110100000",
58697=>"010110110",
58698=>"001000100",
58699=>"000111011",
58700=>"110000000",
58701=>"110101101",
58702=>"011011000",
58703=>"000000100",
58704=>"010111001",
58705=>"111001101",
58706=>"100000000",
58707=>"011101000",
58708=>"111010010",
58709=>"111101111",
58710=>"111111001",
58711=>"111100100",
58712=>"001011101",
58713=>"001101111",
58714=>"001001100",
58715=>"110111100",
58716=>"011110011",
58717=>"100101000",
58718=>"111111111",
58719=>"000000011",
58720=>"110010010",
58721=>"000010000",
58722=>"111010000",
58723=>"000010001",
58724=>"010001000",
58725=>"010011000",
58726=>"010011000",
58727=>"000111111",
58728=>"110000010",
58729=>"111100100",
58730=>"010010111",
58731=>"100100110",
58732=>"000000110",
58733=>"001101101",
58734=>"100100100",
58735=>"001000000",
58736=>"010010001",
58737=>"110100110",
58738=>"011000000",
58739=>"001011011",
58740=>"110100111",
58741=>"001101110",
58742=>"110010010",
58743=>"110010000",
58744=>"110111110",
58745=>"000101011",
58746=>"001101011",
58747=>"000100111",
58748=>"000000000",
58749=>"000000111",
58750=>"000001010",
58751=>"010011010",
58752=>"111000100",
58753=>"011000101",
58754=>"110100110",
58755=>"000000110",
58756=>"000010110",
58757=>"000010000",
58758=>"010110000",
58759=>"101111000",
58760=>"010011001",
58761=>"001001011",
58762=>"001100110",
58763=>"010100101",
58764=>"100100101",
58765=>"110110110",
58766=>"111101011",
58767=>"001000000",
58768=>"111101111",
58769=>"011111000",
58770=>"011010110",
58771=>"100100011",
58772=>"000100110",
58773=>"100000100",
58774=>"110010110",
58775=>"100010011",
58776=>"110000010",
58777=>"101010100",
58778=>"110110111",
58779=>"100100000",
58780=>"000100001",
58781=>"100111110",
58782=>"011000010",
58783=>"011100100",
58784=>"110100110",
58785=>"011111101",
58786=>"000100110",
58787=>"000000010",
58788=>"010000010",
58789=>"000000010",
58790=>"001111001",
58791=>"010110100",
58792=>"000000011",
58793=>"100111011",
58794=>"100000111",
58795=>"011101101",
58796=>"101011011",
58797=>"110010010",
58798=>"000000011",
58799=>"100110110",
58800=>"000010110",
58801=>"000100000",
58802=>"100100000",
58803=>"010100000",
58804=>"110111110",
58805=>"001011001",
58806=>"101100101",
58807=>"000000011",
58808=>"111111101",
58809=>"000001011",
58810=>"111001101",
58811=>"010100110",
58812=>"100000001",
58813=>"110111111",
58814=>"111000111",
58815=>"001101111",
58816=>"000100100",
58817=>"110110100",
58818=>"111100110",
58819=>"011111001",
58820=>"000100111",
58821=>"011111011",
58822=>"000000110",
58823=>"110111111",
58824=>"111110011",
58825=>"011011001",
58826=>"000000000",
58827=>"001000110",
58828=>"100010010",
58829=>"100110110",
58830=>"101100000",
58831=>"001100000",
58832=>"000001011",
58833=>"011101100",
58834=>"001000101",
58835=>"110100100",
58836=>"110110110",
58837=>"110001111",
58838=>"000000010",
58839=>"000000000",
58840=>"011011010",
58841=>"101111110",
58842=>"001100000",
58843=>"000100101",
58844=>"100000000",
58845=>"100110001",
58846=>"011001011",
58847=>"100100000",
58848=>"000110010",
58849=>"011101001",
58850=>"000000001",
58851=>"011001000",
58852=>"001000010",
58853=>"011111111",
58854=>"101001001",
58855=>"011111100",
58856=>"000110111",
58857=>"100001111",
58858=>"011100100",
58859=>"011100111",
58860=>"101100000",
58861=>"111100110",
58862=>"111000011",
58863=>"010000100",
58864=>"000000101",
58865=>"000000100",
58866=>"010010000",
58867=>"000000110",
58868=>"000100011",
58869=>"100011101",
58870=>"000100110",
58871=>"000100110",
58872=>"111100110",
58873=>"100110111",
58874=>"000100110",
58875=>"100111011",
58876=>"111110110",
58877=>"001000101",
58878=>"100100111",
58879=>"110010000",
58880=>"011011000",
58881=>"011100001",
58882=>"101000000",
58883=>"111100111",
58884=>"110111111",
58885=>"111101000",
58886=>"010010000",
58887=>"111111110",
58888=>"011010000",
58889=>"110010011",
58890=>"100111111",
58891=>"111000100",
58892=>"100000011",
58893=>"110110100",
58894=>"000001111",
58895=>"011101001",
58896=>"111111000",
58897=>"101111111",
58898=>"010110011",
58899=>"110010101",
58900=>"011111111",
58901=>"111010111",
58902=>"100101000",
58903=>"111100111",
58904=>"101000010",
58905=>"001110000",
58906=>"111000000",
58907=>"000010111",
58908=>"010000101",
58909=>"101001101",
58910=>"010011111",
58911=>"000101100",
58912=>"111001001",
58913=>"000000010",
58914=>"000000000",
58915=>"110111011",
58916=>"000011000",
58917=>"110110000",
58918=>"101000000",
58919=>"000000111",
58920=>"011011000",
58921=>"011000000",
58922=>"001100110",
58923=>"010000000",
58924=>"100001011",
58925=>"101000100",
58926=>"000001011",
58927=>"000000000",
58928=>"011000111",
58929=>"010110110",
58930=>"000000001",
58931=>"010010111",
58932=>"010111000",
58933=>"000000010",
58934=>"110111110",
58935=>"010000101",
58936=>"111111000",
58937=>"101000101",
58938=>"000110000",
58939=>"111101101",
58940=>"100110100",
58941=>"111101110",
58942=>"000000100",
58943=>"100111111",
58944=>"111111011",
58945=>"111111000",
58946=>"000000111",
58947=>"111011111",
58948=>"001001111",
58949=>"100000101",
58950=>"000000000",
58951=>"111111000",
58952=>"100000000",
58953=>"101000000",
58954=>"101100101",
58955=>"000111111",
58956=>"111010111",
58957=>"100100110",
58958=>"011011011",
58959=>"000000011",
58960=>"010111111",
58961=>"111010011",
58962=>"110111111",
58963=>"011100100",
58964=>"010010000",
58965=>"001111110",
58966=>"011011001",
58967=>"101000000",
58968=>"100100110",
58969=>"100100100",
58970=>"011111110",
58971=>"000100111",
58972=>"010111010",
58973=>"000001000",
58974=>"000000100",
58975=>"001001111",
58976=>"001000100",
58977=>"000100011",
58978=>"000000000",
58979=>"100111001",
58980=>"000110000",
58981=>"001100100",
58982=>"010010000",
58983=>"010100000",
58984=>"000110111",
58985=>"000010001",
58986=>"010000010",
58987=>"111000000",
58988=>"100100000",
58989=>"000101000",
58990=>"000000101",
58991=>"000000110",
58992=>"000100100",
58993=>"001010101",
58994=>"011111011",
58995=>"000000000",
58996=>"000100111",
58997=>"101100101",
58998=>"100100101",
58999=>"111000101",
59000=>"000111010",
59001=>"010000111",
59002=>"000111111",
59003=>"111100011",
59004=>"100110010",
59005=>"110001001",
59006=>"111110110",
59007=>"000100000",
59008=>"000000001",
59009=>"111000000",
59010=>"010011010",
59011=>"111000111",
59012=>"000011111",
59013=>"111100101",
59014=>"011011000",
59015=>"000000100",
59016=>"000011011",
59017=>"000000000",
59018=>"010111110",
59019=>"100111110",
59020=>"001000000",
59021=>"101000111",
59022=>"101001010",
59023=>"101000000",
59024=>"001011001",
59025=>"111111000",
59026=>"011100000",
59027=>"000010011",
59028=>"000010010",
59029=>"111000001",
59030=>"000010111",
59031=>"110100100",
59032=>"000000000",
59033=>"100111111",
59034=>"010011011",
59035=>"111110010",
59036=>"010000000",
59037=>"001000010",
59038=>"010110001",
59039=>"000000000",
59040=>"000100100",
59041=>"111010000",
59042=>"101000100",
59043=>"000000111",
59044=>"000100111",
59045=>"001001011",
59046=>"111001001",
59047=>"010111011",
59048=>"000000111",
59049=>"011000000",
59050=>"000000011",
59051=>"011011011",
59052=>"111111000",
59053=>"111100000",
59054=>"110100011",
59055=>"100100010",
59056=>"111101100",
59057=>"000101000",
59058=>"000111000",
59059=>"000000011",
59060=>"111111111",
59061=>"111111100",
59062=>"111011011",
59063=>"001011000",
59064=>"001011001",
59065=>"000100011",
59066=>"110000000",
59067=>"001111110",
59068=>"010001101",
59069=>"111111111",
59070=>"000111111",
59071=>"011000000",
59072=>"110010000",
59073=>"000000000",
59074=>"011111101",
59075=>"001111110",
59076=>"000001101",
59077=>"101100010",
59078=>"101110111",
59079=>"111110000",
59080=>"000011000",
59081=>"101111000",
59082=>"111010000",
59083=>"001001001",
59084=>"000000010",
59085=>"001011010",
59086=>"111111000",
59087=>"111010000",
59088=>"010000110",
59089=>"101111000",
59090=>"000000010",
59091=>"010111100",
59092=>"101101111",
59093=>"000100000",
59094=>"101101101",
59095=>"010101011",
59096=>"101100100",
59097=>"000000010",
59098=>"000000001",
59099=>"000100100",
59100=>"111101110",
59101=>"001111000",
59102=>"101101000",
59103=>"010011101",
59104=>"000111010",
59105=>"000001000",
59106=>"000000000",
59107=>"001001111",
59108=>"000100011",
59109=>"111101111",
59110=>"111101110",
59111=>"000101101",
59112=>"111000000",
59113=>"000000111",
59114=>"011111000",
59115=>"111111111",
59116=>"000000000",
59117=>"000000000",
59118=>"000000000",
59119=>"111000001",
59120=>"010000101",
59121=>"001111111",
59122=>"000000010",
59123=>"111111011",
59124=>"110111111",
59125=>"000101101",
59126=>"100000000",
59127=>"010000100",
59128=>"000000010",
59129=>"100000010",
59130=>"111000101",
59131=>"000111110",
59132=>"011011000",
59133=>"111000000",
59134=>"010101101",
59135=>"101000101",
59136=>"101011001",
59137=>"101111101",
59138=>"000000101",
59139=>"111101111",
59140=>"000101000",
59141=>"110000000",
59142=>"000000010",
59143=>"111101101",
59144=>"100000011",
59145=>"111000000",
59146=>"100110111",
59147=>"111100111",
59148=>"000011001",
59149=>"000000000",
59150=>"000101001",
59151=>"000101111",
59152=>"010000111",
59153=>"110110111",
59154=>"000001000",
59155=>"111000000",
59156=>"010011101",
59157=>"000000000",
59158=>"111110011",
59159=>"000000111",
59160=>"111111000",
59161=>"011111111",
59162=>"011010101",
59163=>"000000111",
59164=>"101001100",
59165=>"110000100",
59166=>"010010001",
59167=>"111100000",
59168=>"111101000",
59169=>"100000000",
59170=>"000001000",
59171=>"110001101",
59172=>"111000100",
59173=>"100110111",
59174=>"111111010",
59175=>"000101111",
59176=>"111111010",
59177=>"000110010",
59178=>"000000000",
59179=>"110000000",
59180=>"101000000",
59181=>"111100110",
59182=>"100000001",
59183=>"010001111",
59184=>"000110111",
59185=>"000000000",
59186=>"000011111",
59187=>"000111101",
59188=>"100000111",
59189=>"111110000",
59190=>"110010000",
59191=>"101000000",
59192=>"011001111",
59193=>"111100101",
59194=>"000000111",
59195=>"100101101",
59196=>"100100100",
59197=>"000101101",
59198=>"000000000",
59199=>"111111010",
59200=>"100011111",
59201=>"101100001",
59202=>"111111111",
59203=>"011111010",
59204=>"000010010",
59205=>"000000000",
59206=>"010000000",
59207=>"011111011",
59208=>"000000101",
59209=>"000100011",
59210=>"101101111",
59211=>"000010111",
59212=>"101001011",
59213=>"010011000",
59214=>"000111101",
59215=>"000001111",
59216=>"101111000",
59217=>"010010000",
59218=>"000000100",
59219=>"011101000",
59220=>"101101111",
59221=>"001110000",
59222=>"001011010",
59223=>"001001101",
59224=>"000100011",
59225=>"111101000",
59226=>"111100100",
59227=>"000100111",
59228=>"000000111",
59229=>"100001010",
59230=>"010010011",
59231=>"100011010",
59232=>"111111111",
59233=>"000111111",
59234=>"101000111",
59235=>"001001001",
59236=>"000100001",
59237=>"100111011",
59238=>"000110000",
59239=>"111000000",
59240=>"010110000",
59241=>"010111111",
59242=>"111010010",
59243=>"111000101",
59244=>"000000100",
59245=>"010111110",
59246=>"111111111",
59247=>"100010111",
59248=>"100000111",
59249=>"100000111",
59250=>"010000000",
59251=>"000000011",
59252=>"000100111",
59253=>"101000000",
59254=>"000010111",
59255=>"001111010",
59256=>"001000101",
59257=>"000101101",
59258=>"000000110",
59259=>"101000000",
59260=>"101110000",
59261=>"110110000",
59262=>"111100101",
59263=>"101000111",
59264=>"010010000",
59265=>"101000101",
59266=>"000011111",
59267=>"000010111",
59268=>"000101111",
59269=>"111111101",
59270=>"011001001",
59271=>"000000011",
59272=>"111110000",
59273=>"101100100",
59274=>"010111111",
59275=>"101000000",
59276=>"010111000",
59277=>"101101111",
59278=>"000101101",
59279=>"000000100",
59280=>"011100000",
59281=>"100100000",
59282=>"010000101",
59283=>"000000011",
59284=>"001001100",
59285=>"000000000",
59286=>"010011000",
59287=>"100011011",
59288=>"011111111",
59289=>"111000000",
59290=>"001010011",
59291=>"000000000",
59292=>"100100101",
59293=>"111111000",
59294=>"101101000",
59295=>"000100000",
59296=>"100101011",
59297=>"010111010",
59298=>"001101111",
59299=>"101111110",
59300=>"110010100",
59301=>"010110110",
59302=>"100110011",
59303=>"000000110",
59304=>"111111000",
59305=>"000010101",
59306=>"001111111",
59307=>"000000000",
59308=>"000111101",
59309=>"001101111",
59310=>"100100100",
59311=>"111110000",
59312=>"010111111",
59313=>"000101100",
59314=>"000000010",
59315=>"000000100",
59316=>"101011011",
59317=>"111010000",
59318=>"000011011",
59319=>"001101111",
59320=>"000000001",
59321=>"100110100",
59322=>"111000001",
59323=>"010111111",
59324=>"000000100",
59325=>"001011111",
59326=>"001011011",
59327=>"111000001",
59328=>"001000101",
59329=>"010110111",
59330=>"010111011",
59331=>"000100011",
59332=>"000000111",
59333=>"100000001",
59334=>"110001000",
59335=>"000010000",
59336=>"000010101",
59337=>"010010000",
59338=>"111111000",
59339=>"101000101",
59340=>"010000000",
59341=>"111000001",
59342=>"101111100",
59343=>"000000000",
59344=>"111100111",
59345=>"100110110",
59346=>"000000110",
59347=>"000111111",
59348=>"100000001",
59349=>"010100001",
59350=>"101101101",
59351=>"010110101",
59352=>"100000101",
59353=>"100000000",
59354=>"000011000",
59355=>"000110010",
59356=>"001011110",
59357=>"101011111",
59358=>"010111000",
59359=>"010100000",
59360=>"010000001",
59361=>"001100101",
59362=>"111000111",
59363=>"110001001",
59364=>"000111101",
59365=>"110010010",
59366=>"111000010",
59367=>"101011001",
59368=>"010000011",
59369=>"101000101",
59370=>"000001011",
59371=>"000011000",
59372=>"010010111",
59373=>"010111000",
59374=>"000000000",
59375=>"000000010",
59376=>"101000000",
59377=>"001000100",
59378=>"110110001",
59379=>"101000001",
59380=>"111110100",
59381=>"001000101",
59382=>"000000000",
59383=>"001000011",
59384=>"101000111",
59385=>"000000111",
59386=>"110110000",
59387=>"111000001",
59388=>"101000111",
59389=>"011000101",
59390=>"101110001",
59391=>"000000010",
59392=>"010011011",
59393=>"001000110",
59394=>"111000000",
59395=>"100000001",
59396=>"010000011",
59397=>"110110000",
59398=>"000000000",
59399=>"111011110",
59400=>"010001011",
59401=>"000000000",
59402=>"110100000",
59403=>"000000001",
59404=>"111000000",
59405=>"000111111",
59406=>"001001011",
59407=>"111101000",
59408=>"010111101",
59409=>"000001001",
59410=>"110001000",
59411=>"110010000",
59412=>"111111001",
59413=>"101100000",
59414=>"000011111",
59415=>"111000000",
59416=>"010001001",
59417=>"111111111",
59418=>"000111010",
59419=>"000111011",
59420=>"010101001",
59421=>"110000100",
59422=>"100010000",
59423=>"111000000",
59424=>"000000000",
59425=>"000010000",
59426=>"001101111",
59427=>"000100110",
59428=>"000100001",
59429=>"010010001",
59430=>"000000110",
59431=>"000011010",
59432=>"000110010",
59433=>"110111111",
59434=>"111000100",
59435=>"000001000",
59436=>"010111110",
59437=>"000011001",
59438=>"000000000",
59439=>"110001000",
59440=>"000000111",
59441=>"000111101",
59442=>"001000100",
59443=>"110111001",
59444=>"001000000",
59445=>"000000000",
59446=>"000111101",
59447=>"011000000",
59448=>"110011000",
59449=>"111000000",
59450=>"111101000",
59451=>"000110101",
59452=>"000110111",
59453=>"000001000",
59454=>"001000001",
59455=>"011111111",
59456=>"101110110",
59457=>"100110011",
59458=>"000000000",
59459=>"000011000",
59460=>"111111111",
59461=>"010000101",
59462=>"000111000",
59463=>"111111101",
59464=>"110111111",
59465=>"011001011",
59466=>"111101111",
59467=>"111000001",
59468=>"000110110",
59469=>"111011000",
59470=>"000011011",
59471=>"010110110",
59472=>"000000010",
59473=>"000111100",
59474=>"111011111",
59475=>"010011100",
59476=>"110000000",
59477=>"110111110",
59478=>"010011001",
59479=>"010010011",
59480=>"000111110",
59481=>"000101111",
59482=>"000011111",
59483=>"000000000",
59484=>"001000111",
59485=>"111000001",
59486=>"011011010",
59487=>"010100000",
59488=>"000110110",
59489=>"010110111",
59490=>"001000111",
59491=>"000100110",
59492=>"011011001",
59493=>"111000000",
59494=>"100111111",
59495=>"110000000",
59496=>"010111110",
59497=>"111000000",
59498=>"000111010",
59499=>"111011111",
59500=>"111001000",
59501=>"000000000",
59502=>"011101111",
59503=>"110100001",
59504=>"000110111",
59505=>"111001111",
59506=>"000010111",
59507=>"001100011",
59508=>"000111111",
59509=>"000000001",
59510=>"110000000",
59511=>"000111000",
59512=>"111010000",
59513=>"111011011",
59514=>"000000010",
59515=>"110000001",
59516=>"111000110",
59517=>"000100000",
59518=>"111111000",
59519=>"111000100",
59520=>"111010000",
59521=>"111000010",
59522=>"011111110",
59523=>"111001001",
59524=>"000110000",
59525=>"111001001",
59526=>"100110111",
59527=>"100100110",
59528=>"011111111",
59529=>"111100000",
59530=>"000000101",
59531=>"101010000",
59532=>"111000010",
59533=>"111100000",
59534=>"111000000",
59535=>"000000000",
59536=>"000110111",
59537=>"110110111",
59538=>"101111111",
59539=>"111000110",
59540=>"110110111",
59541=>"111000000",
59542=>"001000011",
59543=>"000011001",
59544=>"000000000",
59545=>"111011110",
59546=>"010111111",
59547=>"010001000",
59548=>"101000101",
59549=>"111000000",
59550=>"000000000",
59551=>"111000000",
59552=>"011100011",
59553=>"000111101",
59554=>"111001001",
59555=>"000000001",
59556=>"111010000",
59557=>"011111111",
59558=>"000111100",
59559=>"010000010",
59560=>"000111100",
59561=>"000111111",
59562=>"010011111",
59563=>"000110001",
59564=>"101110000",
59565=>"000000001",
59566=>"010100001",
59567=>"111100000",
59568=>"000000000",
59569=>"001001001",
59570=>"101010000",
59571=>"010000100",
59572=>"010111110",
59573=>"001000100",
59574=>"000110111",
59575=>"000111111",
59576=>"000110111",
59577=>"101011101",
59578=>"011111011",
59579=>"111110010",
59580=>"100000000",
59581=>"111111111",
59582=>"000110111",
59583=>"000000001",
59584=>"111101001",
59585=>"000000000",
59586=>"000000111",
59587=>"010110000",
59588=>"101000000",
59589=>"101101100",
59590=>"110100100",
59591=>"000110000",
59592=>"010001101",
59593=>"101110110",
59594=>"101101111",
59595=>"101000000",
59596=>"111000000",
59597=>"110001000",
59598=>"101010010",
59599=>"000010111",
59600=>"010000000",
59601=>"000110110",
59602=>"110110110",
59603=>"111110001",
59604=>"111000000",
59605=>"111000110",
59606=>"111000011",
59607=>"010011000",
59608=>"111001000",
59609=>"000000101",
59610=>"001001000",
59611=>"111000000",
59612=>"010111101",
59613=>"010111011",
59614=>"001110010",
59615=>"111111100",
59616=>"001001110",
59617=>"000000001",
59618=>"111001000",
59619=>"000001111",
59620=>"111000000",
59621=>"111001111",
59622=>"100001001",
59623=>"111111001",
59624=>"111111111",
59625=>"010010111",
59626=>"011001000",
59627=>"000000110",
59628=>"000110111",
59629=>"000000111",
59630=>"000000000",
59631=>"010001110",
59632=>"011110100",
59633=>"101001111",
59634=>"111000000",
59635=>"111001001",
59636=>"000111111",
59637=>"010011011",
59638=>"101000000",
59639=>"010000101",
59640=>"110010000",
59641=>"111000000",
59642=>"111000001",
59643=>"000110110",
59644=>"111110100",
59645=>"111101001",
59646=>"000100100",
59647=>"110000000",
59648=>"001101111",
59649=>"011000110",
59650=>"000101111",
59651=>"010011000",
59652=>"000100111",
59653=>"110101100",
59654=>"111011111",
59655=>"011010110",
59656=>"111001111",
59657=>"000000000",
59658=>"000110110",
59659=>"000000000",
59660=>"000011000",
59661=>"111100111",
59662=>"101101110",
59663=>"110000011",
59664=>"111111001",
59665=>"000110100",
59666=>"110101100",
59667=>"000010111",
59668=>"111110111",
59669=>"101100100",
59670=>"001110110",
59671=>"111111101",
59672=>"000100110",
59673=>"001100100",
59674=>"111101111",
59675=>"000000111",
59676=>"001000101",
59677=>"111111101",
59678=>"111100000",
59679=>"101001001",
59680=>"000010010",
59681=>"101100000",
59682=>"000101111",
59683=>"000101000",
59684=>"101100000",
59685=>"100000100",
59686=>"000000100",
59687=>"001111111",
59688=>"000111000",
59689=>"001101110",
59690=>"011000111",
59691=>"111010000",
59692=>"011011000",
59693=>"010100101",
59694=>"011100110",
59695=>"000111011",
59696=>"000000000",
59697=>"101111111",
59698=>"100100101",
59699=>"111100111",
59700=>"000010000",
59701=>"111111110",
59702=>"110000010",
59703=>"011001101",
59704=>"111101101",
59705=>"111101101",
59706=>"100000000",
59707=>"100011101",
59708=>"001011000",
59709=>"111111111",
59710=>"011010011",
59711=>"111001001",
59712=>"100001000",
59713=>"100101100",
59714=>"111101011",
59715=>"101100110",
59716=>"000100111",
59717=>"111000010",
59718=>"010000101",
59719=>"000010000",
59720=>"110001000",
59721=>"000111101",
59722=>"010100011",
59723=>"101000100",
59724=>"111101111",
59725=>"101101100",
59726=>"000110011",
59727=>"111001001",
59728=>"001000100",
59729=>"111110010",
59730=>"111011111",
59731=>"001001001",
59732=>"010011111",
59733=>"101100000",
59734=>"100000001",
59735=>"111100111",
59736=>"111100101",
59737=>"101011011",
59738=>"101001001",
59739=>"101100000",
59740=>"100101111",
59741=>"010001011",
59742=>"101101111",
59743=>"101001100",
59744=>"011000000",
59745=>"111010000",
59746=>"001000100",
59747=>"111100000",
59748=>"000000111",
59749=>"100011001",
59750=>"111100100",
59751=>"000010010",
59752=>"100010111",
59753=>"101000100",
59754=>"100101010",
59755=>"001100111",
59756=>"110000100",
59757=>"000011111",
59758=>"100111111",
59759=>"100100111",
59760=>"001110000",
59761=>"100110110",
59762=>"011000110",
59763=>"000000000",
59764=>"000011111",
59765=>"101000000",
59766=>"100000111",
59767=>"000011010",
59768=>"000000000",
59769=>"101110111",
59770=>"100000111",
59771=>"001000101",
59772=>"111111111",
59773=>"000000000",
59774=>"001000110",
59775=>"101000110",
59776=>"010000000",
59777=>"111001001",
59778=>"000000000",
59779=>"011111110",
59780=>"111110111",
59781=>"010110110",
59782=>"011001000",
59783=>"001001000",
59784=>"000101100",
59785=>"101100111",
59786=>"010111011",
59787=>"000000000",
59788=>"100100100",
59789=>"000010000",
59790=>"000011010",
59791=>"000000000",
59792=>"000001000",
59793=>"101001101",
59794=>"101100111",
59795=>"100000000",
59796=>"000111001",
59797=>"100100101",
59798=>"101111100",
59799=>"110100100",
59800=>"001010000",
59801=>"101000000",
59802=>"000010000",
59803=>"000010100",
59804=>"111100100",
59805=>"000000000",
59806=>"111111100",
59807=>"111101111",
59808=>"000000000",
59809=>"111111111",
59810=>"000110111",
59811=>"000100100",
59812=>"000001111",
59813=>"100110000",
59814=>"001101011",
59815=>"100111011",
59816=>"001011111",
59817=>"001101000",
59818=>"100000101",
59819=>"100100100",
59820=>"100100100",
59821=>"111101111",
59822=>"110110101",
59823=>"010010000",
59824=>"101000000",
59825=>"011100111",
59826=>"101101110",
59827=>"000001110",
59828=>"010011101",
59829=>"010010000",
59830=>"000011011",
59831=>"000011000",
59832=>"010100000",
59833=>"110110100",
59834=>"011011011",
59835=>"001000111",
59836=>"000010110",
59837=>"011111111",
59838=>"011100110",
59839=>"000111000",
59840=>"111101101",
59841=>"000000000",
59842=>"110010100",
59843=>"000011011",
59844=>"101110010",
59845=>"101100100",
59846=>"011011100",
59847=>"101100111",
59848=>"100101111",
59849=>"111000111",
59850=>"010111001",
59851=>"001101000",
59852=>"110011010",
59853=>"000111110",
59854=>"000011000",
59855=>"101000100",
59856=>"111101110",
59857=>"011001111",
59858=>"000000111",
59859=>"110111001",
59860=>"101100000",
59861=>"011001000",
59862=>"111101111",
59863=>"010010000",
59864=>"000000001",
59865=>"000000111",
59866=>"000010000",
59867=>"000011000",
59868=>"101011101",
59869=>"011001111",
59870=>"010111111",
59871=>"000000011",
59872=>"101100101",
59873=>"111001100",
59874=>"010011010",
59875=>"101001001",
59876=>"101000001",
59877=>"101011011",
59878=>"111111111",
59879=>"000010000",
59880=>"000000010",
59881=>"111010000",
59882=>"110011011",
59883=>"100111011",
59884=>"000000011",
59885=>"100000000",
59886=>"110000001",
59887=>"100000010",
59888=>"000000001",
59889=>"001000001",
59890=>"000000000",
59891=>"111110011",
59892=>"110000001",
59893=>"101001011",
59894=>"000000000",
59895=>"000011000",
59896=>"110001000",
59897=>"111110001",
59898=>"101100111",
59899=>"011111100",
59900=>"101100001",
59901=>"000001011",
59902=>"001011001",
59903=>"001000000",
59904=>"001101100",
59905=>"100001111",
59906=>"101000101",
59907=>"000101011",
59908=>"001001011",
59909=>"111110100",
59910=>"100000100",
59911=>"111111111",
59912=>"000000000",
59913=>"100000000",
59914=>"101000000",
59915=>"111101111",
59916=>"000001111",
59917=>"010111001",
59918=>"001001011",
59919=>"111111010",
59920=>"011000010",
59921=>"101000111",
59922=>"111100001",
59923=>"011011000",
59924=>"001010000",
59925=>"101000000",
59926=>"111001000",
59927=>"101101110",
59928=>"101000110",
59929=>"111111101",
59930=>"000000100",
59931=>"100000000",
59932=>"010010010",
59933=>"000000000",
59934=>"110110000",
59935=>"000010010",
59936=>"010011100",
59937=>"010111111",
59938=>"100011010",
59939=>"000000000",
59940=>"000011011",
59941=>"110110011",
59942=>"000010010",
59943=>"011010001",
59944=>"011111001",
59945=>"000110110",
59946=>"101001001",
59947=>"101111100",
59948=>"001011011",
59949=>"101000011",
59950=>"111100000",
59951=>"010111111",
59952=>"010110110",
59953=>"001011011",
59954=>"111000010",
59955=>"100101101",
59956=>"010000000",
59957=>"001001000",
59958=>"100000000",
59959=>"000100101",
59960=>"001101101",
59961=>"001000000",
59962=>"111101000",
59963=>"000100111",
59964=>"001110000",
59965=>"111111010",
59966=>"100000000",
59967=>"111010000",
59968=>"111011011",
59969=>"000000101",
59970=>"100000011",
59971=>"111000100",
59972=>"110000011",
59973=>"111010111",
59974=>"101000000",
59975=>"000001000",
59976=>"010010011",
59977=>"001111001",
59978=>"111100001",
59979=>"011111011",
59980=>"000100000",
59981=>"000100100",
59982=>"000110110",
59983=>"100110111",
59984=>"000101111",
59985=>"010110111",
59986=>"011011000",
59987=>"111101000",
59988=>"111000110",
59989=>"111110110",
59990=>"011100101",
59991=>"001000111",
59992=>"111111100",
59993=>"000111000",
59994=>"110110111",
59995=>"010100111",
59996=>"000100000",
59997=>"001001001",
59998=>"100010000",
59999=>"111000000",
60000=>"010111110",
60001=>"000000000",
60002=>"110111000",
60003=>"111101000",
60004=>"010001101",
60005=>"001001101",
60006=>"010010000",
60007=>"001001000",
60008=>"000000101",
60009=>"110000101",
60010=>"111111101",
60011=>"010011110",
60012=>"001000110",
60013=>"001101000",
60014=>"111101111",
60015=>"100000001",
60016=>"110110001",
60017=>"000100101",
60018=>"011000110",
60019=>"011111000",
60020=>"111010010",
60021=>"000000010",
60022=>"100000101",
60023=>"011010000",
60024=>"111000001",
60025=>"111010000",
60026=>"111010010",
60027=>"101111111",
60028=>"000110110",
60029=>"010100000",
60030=>"011000011",
60031=>"101100000",
60032=>"000101110",
60033=>"010111111",
60034=>"111000010",
60035=>"110001001",
60036=>"010000000",
60037=>"111111111",
60038=>"111101110",
60039=>"011000000",
60040=>"000100000",
60041=>"000000000",
60042=>"100100010",
60043=>"011001000",
60044=>"001010000",
60045=>"000010110",
60046=>"101001001",
60047=>"001001000",
60048=>"000100100",
60049=>"000100111",
60050=>"000100000",
60051=>"111001101",
60052=>"000000000",
60053=>"111000101",
60054=>"111101001",
60055=>"010011011",
60056=>"000110111",
60057=>"000111111",
60058=>"111101101",
60059=>"111101011",
60060=>"111101101",
60061=>"111101101",
60062=>"101101001",
60063=>"000000101",
60064=>"000010000",
60065=>"101100000",
60066=>"011001001",
60067=>"101001010",
60068=>"000000010",
60069=>"000000010",
60070=>"010110100",
60071=>"101000100",
60072=>"101100000",
60073=>"010010111",
60074=>"111100000",
60075=>"010101000",
60076=>"010101001",
60077=>"111101111",
60078=>"001001001",
60079=>"101000111",
60080=>"011101000",
60081=>"111010011",
60082=>"000010010",
60083=>"000001000",
60084=>"101000001",
60085=>"000100000",
60086=>"111111111",
60087=>"000111101",
60088=>"100011011",
60089=>"110000110",
60090=>"011000001",
60091=>"111111001",
60092=>"000000000",
60093=>"111111111",
60094=>"000100100",
60095=>"001101010",
60096=>"101001001",
60097=>"111100111",
60098=>"111100110",
60099=>"011101001",
60100=>"000101010",
60101=>"000101111",
60102=>"000000011",
60103=>"000010000",
60104=>"101001101",
60105=>"010000000",
60106=>"101101101",
60107=>"111001101",
60108=>"111000100",
60109=>"000010011",
60110=>"010111101",
60111=>"010111100",
60112=>"111111000",
60113=>"111101110",
60114=>"010011101",
60115=>"111101010",
60116=>"000010110",
60117=>"001101111",
60118=>"000111111",
60119=>"111100101",
60120=>"000110000",
60121=>"001001100",
60122=>"000000000",
60123=>"100000101",
60124=>"111001000",
60125=>"111011000",
60126=>"010111110",
60127=>"010111011",
60128=>"000011010",
60129=>"111100100",
60130=>"011010000",
60131=>"011101000",
60132=>"111000101",
60133=>"000010110",
60134=>"011111111",
60135=>"001111000",
60136=>"000000011",
60137=>"001000000",
60138=>"100000000",
60139=>"000000000",
60140=>"000000011",
60141=>"010001111",
60142=>"000000100",
60143=>"001011010",
60144=>"010111000",
60145=>"001000110",
60146=>"111000000",
60147=>"010000000",
60148=>"110101110",
60149=>"111101101",
60150=>"000000000",
60151=>"101101001",
60152=>"111001001",
60153=>"111001010",
60154=>"110000000",
60155=>"101101000",
60156=>"001101101",
60157=>"101000000",
60158=>"110110111",
60159=>"101000000",
60160=>"010100100",
60161=>"010000001",
60162=>"111001001",
60163=>"101001110",
60164=>"011011010",
60165=>"111110000",
60166=>"000110111",
60167=>"101000010",
60168=>"100101100",
60169=>"001001111",
60170=>"010111001",
60171=>"000001111",
60172=>"101000001",
60173=>"111001001",
60174=>"100110111",
60175=>"001000001",
60176=>"100000100",
60177=>"111110110",
60178=>"111111100",
60179=>"011000000",
60180=>"011110000",
60181=>"111110010",
60182=>"010101101",
60183=>"100000110",
60184=>"111110000",
60185=>"010111011",
60186=>"010011100",
60187=>"000000111",
60188=>"001010111",
60189=>"000000000",
60190=>"111010100",
60191=>"000011101",
60192=>"101101111",
60193=>"010000001",
60194=>"000000011",
60195=>"111111111",
60196=>"000101100",
60197=>"000010011",
60198=>"111110010",
60199=>"010001001",
60200=>"000111111",
60201=>"001111111",
60202=>"110000000",
60203=>"001101111",
60204=>"111111100",
60205=>"101111010",
60206=>"010000110",
60207=>"000010000",
60208=>"010010000",
60209=>"000100100",
60210=>"110111001",
60211=>"000111111",
60212=>"111111111",
60213=>"001001000",
60214=>"110100011",
60215=>"001101110",
60216=>"110100010",
60217=>"000010011",
60218=>"000111100",
60219=>"100111111",
60220=>"100000011",
60221=>"011111101",
60222=>"000000101",
60223=>"110010001",
60224=>"110111111",
60225=>"000000100",
60226=>"000000111",
60227=>"001100000",
60228=>"111001011",
60229=>"111100101",
60230=>"000110010",
60231=>"010111111",
60232=>"011000111",
60233=>"011110111",
60234=>"100100111",
60235=>"110000100",
60236=>"111001000",
60237=>"001011111",
60238=>"100110100",
60239=>"010111111",
60240=>"001111000",
60241=>"110111000",
60242=>"011010100",
60243=>"000000100",
60244=>"000100000",
60245=>"100100110",
60246=>"000101101",
60247=>"000110101",
60248=>"000011010",
60249=>"001001000",
60250=>"001111000",
60251=>"010011010",
60252=>"010000100",
60253=>"000000000",
60254=>"111111000",
60255=>"100000000",
60256=>"111001101",
60257=>"000111110",
60258=>"101000111",
60259=>"101100000",
60260=>"001000000",
60261=>"001100100",
60262=>"111111000",
60263=>"000000100",
60264=>"111000110",
60265=>"000111111",
60266=>"111000000",
60267=>"111010010",
60268=>"000101111",
60269=>"010111011",
60270=>"010111010",
60271=>"010010010",
60272=>"001001111",
60273=>"000000111",
60274=>"011001110",
60275=>"000111000",
60276=>"111000011",
60277=>"101000011",
60278=>"000000101",
60279=>"011000101",
60280=>"111000101",
60281=>"111000111",
60282=>"101000001",
60283=>"000000001",
60284=>"000101001",
60285=>"010000001",
60286=>"000100000",
60287=>"100111101",
60288=>"010011010",
60289=>"100010010",
60290=>"111000010",
60291=>"011000010",
60292=>"111101101",
60293=>"000000010",
60294=>"011011110",
60295=>"000001011",
60296=>"100100100",
60297=>"000000111",
60298=>"000010101",
60299=>"000000111",
60300=>"000000000",
60301=>"111111010",
60302=>"001100110",
60303=>"001000011",
60304=>"011011001",
60305=>"000010111",
60306=>"010000010",
60307=>"000010111",
60308=>"000000001",
60309=>"111000111",
60310=>"000111000",
60311=>"100110000",
60312=>"111000101",
60313=>"110010010",
60314=>"110010010",
60315=>"000000000",
60316=>"000111010",
60317=>"111100000",
60318=>"010000000",
60319=>"000101111",
60320=>"011011011",
60321=>"001000011",
60322=>"000000001",
60323=>"001110111",
60324=>"010000011",
60325=>"110110100",
60326=>"101111000",
60327=>"101000000",
60328=>"110111110",
60329=>"111000000",
60330=>"111001111",
60331=>"111111111",
60332=>"000010111",
60333=>"100000100",
60334=>"001011011",
60335=>"001101111",
60336=>"101000000",
60337=>"000110110",
60338=>"000100100",
60339=>"000010110",
60340=>"000000000",
60341=>"101100000",
60342=>"111100100",
60343=>"000000101",
60344=>"001000111",
60345=>"000000110",
60346=>"110010000",
60347=>"111011011",
60348=>"000000011",
60349=>"011011011",
60350=>"001001011",
60351=>"100100000",
60352=>"000111110",
60353=>"010111010",
60354=>"111010010",
60355=>"000001000",
60356=>"000000001",
60357=>"110110001",
60358=>"000000111",
60359=>"000111000",
60360=>"110000000",
60361=>"011111010",
60362=>"111110000",
60363=>"010110111",
60364=>"011000001",
60365=>"000101111",
60366=>"001111000",
60367=>"111011110",
60368=>"111011000",
60369=>"001100010",
60370=>"010010011",
60371=>"111101011",
60372=>"111000000",
60373=>"001011000",
60374=>"111111111",
60375=>"110001001",
60376=>"000010010",
60377=>"101000001",
60378=>"100110110",
60379=>"000101001",
60380=>"000001001",
60381=>"111101001",
60382=>"111101101",
60383=>"010000010",
60384=>"010111111",
60385=>"110111111",
60386=>"101001101",
60387=>"001011001",
60388=>"000010000",
60389=>"000000000",
60390=>"111101111",
60391=>"001101100",
60392=>"110000100",
60393=>"000000111",
60394=>"111111110",
60395=>"001101111",
60396=>"000110111",
60397=>"101000001",
60398=>"000000000",
60399=>"000000010",
60400=>"111101001",
60401=>"011011100",
60402=>"000000010",
60403=>"000000001",
60404=>"000001001",
60405=>"010111000",
60406=>"000100000",
60407=>"111100111",
60408=>"111000001",
60409=>"000000111",
60410=>"111010111",
60411=>"111010010",
60412=>"010010000",
60413=>"111111111",
60414=>"000100000",
60415=>"111001000",
60416=>"111110110",
60417=>"000000000",
60418=>"000000100",
60419=>"111111111",
60420=>"110111101",
60421=>"001001111",
60422=>"111110000",
60423=>"111111111",
60424=>"000001001",
60425=>"000100010",
60426=>"110110110",
60427=>"010000000",
60428=>"000000000",
60429=>"000000111",
60430=>"111110111",
60431=>"000000111",
60432=>"111011000",
60433=>"110111111",
60434=>"111110111",
60435=>"000000000",
60436=>"100110111",
60437=>"000000000",
60438=>"111111010",
60439=>"010111011",
60440=>"101001111",
60441=>"000000000",
60442=>"100000111",
60443=>"000001011",
60444=>"111111000",
60445=>"110010101",
60446=>"101111111",
60447=>"010010000",
60448=>"011111111",
60449=>"110000000",
60450=>"111111111",
60451=>"000000000",
60452=>"000000000",
60453=>"100110000",
60454=>"000000001",
60455=>"100100100",
60456=>"100100001",
60457=>"001001100",
60458=>"011011001",
60459=>"011101000",
60460=>"111110100",
60461=>"110000000",
60462=>"111111111",
60463=>"111011111",
60464=>"000010111",
60465=>"000000111",
60466=>"101001000",
60467=>"110110110",
60468=>"111111011",
60469=>"000001000",
60470=>"111000100",
60471=>"000001101",
60472=>"111111111",
60473=>"000000111",
60474=>"011001101",
60475=>"000000000",
60476=>"101101001",
60477=>"111111111",
60478=>"000000000",
60479=>"000010001",
60480=>"101111011",
60481=>"101111000",
60482=>"001000001",
60483=>"001000110",
60484=>"110111111",
60485=>"111111101",
60486=>"000000001",
60487=>"001111111",
60488=>"010000100",
60489=>"110110000",
60490=>"101000000",
60491=>"111101110",
60492=>"000000000",
60493=>"000000011",
60494=>"000110110",
60495=>"010111111",
60496=>"111110111",
60497=>"110110000",
60498=>"000000000",
60499=>"011011111",
60500=>"000000000",
60501=>"100100100",
60502=>"110110110",
60503=>"011111111",
60504=>"100000000",
60505=>"100100010",
60506=>"011001000",
60507=>"100000000",
60508=>"001111011",
60509=>"001011110",
60510=>"000000111",
60511=>"000000110",
60512=>"101000101",
60513=>"010110110",
60514=>"101111111",
60515=>"110110000",
60516=>"100010010",
60517=>"111111111",
60518=>"011000001",
60519=>"100000001",
60520=>"110111111",
60521=>"011110010",
60522=>"001001000",
60523=>"110000000",
60524=>"100111111",
60525=>"000011001",
60526=>"010000000",
60527=>"000000000",
60528=>"110110110",
60529=>"111111000",
60530=>"110011011",
60531=>"000000000",
60532=>"000000100",
60533=>"000000100",
60534=>"111111101",
60535=>"100000011",
60536=>"000000000",
60537=>"000001000",
60538=>"000000000",
60539=>"011111111",
60540=>"100111111",
60541=>"001000001",
60542=>"000000000",
60543=>"000010111",
60544=>"000111101",
60545=>"111111000",
60546=>"000000100",
60547=>"111101111",
60548=>"001000000",
60549=>"000000111",
60550=>"011111110",
60551=>"010010011",
60552=>"011011111",
60553=>"110110100",
60554=>"010111010",
60555=>"000000111",
60556=>"000000000",
60557=>"000000000",
60558=>"111011011",
60559=>"101100100",
60560=>"001011001",
60561=>"011011000",
60562=>"000000000",
60563=>"000000001",
60564=>"010010010",
60565=>"000000000",
60566=>"111011111",
60567=>"110100100",
60568=>"010000000",
60569=>"111000000",
60570=>"000000000",
60571=>"111111111",
60572=>"001100100",
60573=>"000001111",
60574=>"000111000",
60575=>"101000100",
60576=>"011101010",
60577=>"111111001",
60578=>"111111111",
60579=>"010000010",
60580=>"010111100",
60581=>"111111101",
60582=>"100000010",
60583=>"101000001",
60584=>"000000100",
60585=>"011001101",
60586=>"001000101",
60587=>"111000100",
60588=>"001001111",
60589=>"111101111",
60590=>"111111111",
60591=>"010111001",
60592=>"000000001",
60593=>"011111100",
60594=>"011111011",
60595=>"000011001",
60596=>"111001000",
60597=>"011111110",
60598=>"000000100",
60599=>"001111111",
60600=>"111111000",
60601=>"010000100",
60602=>"010000000",
60603=>"000000000",
60604=>"000000000",
60605=>"110111001",
60606=>"000000100",
60607=>"111111010",
60608=>"010010000",
60609=>"000000111",
60610=>"100111110",
60611=>"111001101",
60612=>"000000111",
60613=>"111111100",
60614=>"010111111",
60615=>"001101111",
60616=>"000000101",
60617=>"111001001",
60618=>"101001000",
60619=>"110000000",
60620=>"010000000",
60621=>"000110111",
60622=>"111111110",
60623=>"111111001",
60624=>"000000000",
60625=>"111011111",
60626=>"010010101",
60627=>"111110101",
60628=>"000000111",
60629=>"111111001",
60630=>"110000111",
60631=>"010111111",
60632=>"000110110",
60633=>"000000001",
60634=>"000101000",
60635=>"001001111",
60636=>"111110110",
60637=>"011011000",
60638=>"000000001",
60639=>"011101111",
60640=>"111000000",
60641=>"111111000",
60642=>"000111100",
60643=>"101111011",
60644=>"000000000",
60645=>"000010000",
60646=>"000101101",
60647=>"110110111",
60648=>"000000000",
60649=>"111001000",
60650=>"110111000",
60651=>"111111111",
60652=>"011000001",
60653=>"000000000",
60654=>"000000000",
60655=>"001101111",
60656=>"000000100",
60657=>"010111010",
60658=>"000111111",
60659=>"110010001",
60660=>"001111111",
60661=>"111111101",
60662=>"111000000",
60663=>"100000000",
60664=>"001001000",
60665=>"111110000",
60666=>"111111110",
60667=>"110101000",
60668=>"000000100",
60669=>"111111000",
60670=>"000000110",
60671=>"111111111",
60672=>"100000100",
60673=>"111111111",
60674=>"010010101",
60675=>"000000000",
60676=>"001110010",
60677=>"000000001",
60678=>"100101100",
60679=>"101010111",
60680=>"000001011",
60681=>"011010111",
60682=>"110111001",
60683=>"000000000",
60684=>"000000110",
60685=>"101000100",
60686=>"011010010",
60687=>"111000000",
60688=>"111111111",
60689=>"111111000",
60690=>"101111111",
60691=>"111110111",
60692=>"000111010",
60693=>"000000111",
60694=>"111111111",
60695=>"010111111",
60696=>"111000000",
60697=>"111111111",
60698=>"111000111",
60699=>"010010000",
60700=>"110000010",
60701=>"000000000",
60702=>"000110111",
60703=>"111111111",
60704=>"111001001",
60705=>"011000010",
60706=>"100111100",
60707=>"011000000",
60708=>"110110100",
60709=>"000000000",
60710=>"000000111",
60711=>"111111110",
60712=>"000111000",
60713=>"000100111",
60714=>"000110110",
60715=>"000000100",
60716=>"000110111",
60717=>"111100000",
60718=>"111000000",
60719=>"000011011",
60720=>"111110001",
60721=>"000100101",
60722=>"111001000",
60723=>"111111001",
60724=>"010110010",
60725=>"000011111",
60726=>"111111110",
60727=>"101001101",
60728=>"001101110",
60729=>"000000000",
60730=>"000000111",
60731=>"111111111",
60732=>"000000001",
60733=>"000010111",
60734=>"001000111",
60735=>"100000011",
60736=>"111111101",
60737=>"000000000",
60738=>"101101101",
60739=>"110100010",
60740=>"101101111",
60741=>"100100000",
60742=>"000000000",
60743=>"101001101",
60744=>"001000000",
60745=>"000000110",
60746=>"101100000",
60747=>"000000000",
60748=>"000000110",
60749=>"001111001",
60750=>"000000000",
60751=>"111111000",
60752=>"000110000",
60753=>"111110000",
60754=>"111111111",
60755=>"001110110",
60756=>"001010000",
60757=>"000000010",
60758=>"011111011",
60759=>"000001000",
60760=>"101101111",
60761=>"011110111",
60762=>"010100100",
60763=>"000100110",
60764=>"111111101",
60765=>"111100100",
60766=>"000111111",
60767=>"011001011",
60768=>"000000111",
60769=>"000100000",
60770=>"001000111",
60771=>"010011001",
60772=>"101001001",
60773=>"001111100",
60774=>"111111111",
60775=>"111111111",
60776=>"000000001",
60777=>"011111111",
60778=>"111010111",
60779=>"010101100",
60780=>"000000000",
60781=>"000000000",
60782=>"001000000",
60783=>"000101111",
60784=>"001011011",
60785=>"001000000",
60786=>"111111011",
60787=>"000000010",
60788=>"111111100",
60789=>"111000010",
60790=>"000000011",
60791=>"001001100",
60792=>"110000000",
60793=>"111111101",
60794=>"010010000",
60795=>"111100111",
60796=>"000000001",
60797=>"100001011",
60798=>"000000010",
60799=>"001000111",
60800=>"000111111",
60801=>"000000000",
60802=>"000000000",
60803=>"100000111",
60804=>"100110111",
60805=>"111111010",
60806=>"000000000",
60807=>"001000000",
60808=>"111100010",
60809=>"111111111",
60810=>"111111100",
60811=>"101111111",
60812=>"001000111",
60813=>"111111111",
60814=>"000011011",
60815=>"001000111",
60816=>"001011100",
60817=>"111001000",
60818=>"000000010",
60819=>"001000000",
60820=>"001000000",
60821=>"010111000",
60822=>"110000110",
60823=>"000000001",
60824=>"001101000",
60825=>"101101111",
60826=>"111000110",
60827=>"110010000",
60828=>"000000000",
60829=>"000000000",
60830=>"000100000",
60831=>"000000110",
60832=>"000000000",
60833=>"001000000",
60834=>"101100010",
60835=>"111001100",
60836=>"000001111",
60837=>"001011011",
60838=>"110111111",
60839=>"000000111",
60840=>"010111111",
60841=>"000000110",
60842=>"100100111",
60843=>"000110000",
60844=>"110111111",
60845=>"101101111",
60846=>"000000000",
60847=>"110000110",
60848=>"111100000",
60849=>"001000100",
60850=>"110111100",
60851=>"100110111",
60852=>"110100100",
60853=>"111000111",
60854=>"110111111",
60855=>"100010011",
60856=>"000000000",
60857=>"000000000",
60858=>"111111000",
60859=>"111000000",
60860=>"001000010",
60861=>"011111001",
60862=>"111001110",
60863=>"000100100",
60864=>"001000111",
60865=>"111000000",
60866=>"010010000",
60867=>"000000110",
60868=>"000000101",
60869=>"100110111",
60870=>"000111101",
60871=>"001010011",
60872=>"101101111",
60873=>"000000000",
60874=>"110111111",
60875=>"011000111",
60876=>"111000000",
60877=>"000010110",
60878=>"000010101",
60879=>"111100111",
60880=>"000000110",
60881=>"000000000",
60882=>"000000111",
60883=>"110110010",
60884=>"101101111",
60885=>"001000000",
60886=>"011101111",
60887=>"111101001",
60888=>"001001111",
60889=>"000000000",
60890=>"000000010",
60891=>"000000111",
60892=>"100111111",
60893=>"000000000",
60894=>"000111000",
60895=>"101111111",
60896=>"000000000",
60897=>"111111111",
60898=>"100101000",
60899=>"011001010",
60900=>"101000000",
60901=>"111110101",
60902=>"000000010",
60903=>"000000001",
60904=>"011000011",
60905=>"111011101",
60906=>"011110000",
60907=>"111111111",
60908=>"001001111",
60909=>"000000111",
60910=>"110000000",
60911=>"100000111",
60912=>"000000111",
60913=>"010001001",
60914=>"000110101",
60915=>"011011010",
60916=>"000000010",
60917=>"101101000",
60918=>"101000010",
60919=>"110111111",
60920=>"110010011",
60921=>"001000011",
60922=>"111111111",
60923=>"001000000",
60924=>"111111000",
60925=>"111000000",
60926=>"101010101",
60927=>"000000010",
60928=>"111011111",
60929=>"110000000",
60930=>"000111111",
60931=>"000111000",
60932=>"011000101",
60933=>"100111100",
60934=>"000000111",
60935=>"111010100",
60936=>"000000111",
60937=>"000101000",
60938=>"011011001",
60939=>"101101111",
60940=>"000000111",
60941=>"000000000",
60942=>"110010000",
60943=>"100111101",
60944=>"111010000",
60945=>"111000000",
60946=>"111000000",
60947=>"000000000",
60948=>"101011111",
60949=>"111101000",
60950=>"000000000",
60951=>"111001101",
60952=>"010000000",
60953=>"111011000",
60954=>"000000000",
60955=>"011111000",
60956=>"111110000",
60957=>"010111000",
60958=>"000011111",
60959=>"000111111",
60960=>"111000000",
60961=>"111010000",
60962=>"100110111",
60963=>"000000111",
60964=>"100000100",
60965=>"111111000",
60966=>"111000000",
60967=>"000000011",
60968=>"000000000",
60969=>"111000111",
60970=>"010000000",
60971=>"000100111",
60972=>"111011000",
60973=>"010000000",
60974=>"111000100",
60975=>"001000100",
60976=>"000001000",
60977=>"111110100",
60978=>"111011111",
60979=>"111010000",
60980=>"001000100",
60981=>"000000000",
60982=>"000101111",
60983=>"111101000",
60984=>"000010011",
60985=>"111000000",
60986=>"100000000",
60987=>"000000000",
60988=>"010110001",
60989=>"010100100",
60990=>"000000000",
60991=>"011011000",
60992=>"011110111",
60993=>"111010001",
60994=>"000100000",
60995=>"001001111",
60996=>"000111010",
60997=>"111101101",
60998=>"000000000",
60999=>"000111111",
61000=>"111100000",
61001=>"111000000",
61002=>"101000000",
61003=>"111000000",
61004=>"101000000",
61005=>"011001001",
61006=>"111001100",
61007=>"111101010",
61008=>"100000000",
61009=>"111000111",
61010=>"010111111",
61011=>"001101000",
61012=>"110001000",
61013=>"101000000",
61014=>"000000000",
61015=>"100111000",
61016=>"011110111",
61017=>"111000011",
61018=>"011100100",
61019=>"111010000",
61020=>"111010000",
61021=>"010000000",
61022=>"000000111",
61023=>"100100111",
61024=>"000000010",
61025=>"011000000",
61026=>"000111111",
61027=>"110001001",
61028=>"111001001",
61029=>"000011000",
61030=>"010000000",
61031=>"111000000",
61032=>"000111110",
61033=>"111010000",
61034=>"010011000",
61035=>"111110111",
61036=>"111111111",
61037=>"111000100",
61038=>"000000000",
61039=>"111010000",
61040=>"011000100",
61041=>"111000010",
61042=>"000111110",
61043=>"010000000",
61044=>"111001000",
61045=>"101000000",
61046=>"100111100",
61047=>"000000001",
61048=>"000000011",
61049=>"010010000",
61050=>"101101000",
61051=>"101100110",
61052=>"101011110",
61053=>"110001000",
61054=>"000110010",
61055=>"001111111",
61056=>"000010000",
61057=>"000001111",
61058=>"000000111",
61059=>"111000000",
61060=>"111000000",
61061=>"011000100",
61062=>"110011001",
61063=>"111000000",
61064=>"110100000",
61065=>"100110110",
61066=>"111000000",
61067=>"010011000",
61068=>"000000010",
61069=>"100110110",
61070=>"000000000",
61071=>"111001000",
61072=>"011000001",
61073=>"010111111",
61074=>"001000000",
61075=>"111101101",
61076=>"111100011",
61077=>"100000000",
61078=>"111011111",
61079=>"100100101",
61080=>"100000000",
61081=>"000000111",
61082=>"010100000",
61083=>"000001111",
61084=>"000000011",
61085=>"100000000",
61086=>"010101100",
61087=>"101101111",
61088=>"000001011",
61089=>"011000111",
61090=>"011011000",
61091=>"111001111",
61092=>"000000100",
61093=>"111000000",
61094=>"000101111",
61095=>"111001100",
61096=>"101101000",
61097=>"000000000",
61098=>"101111111",
61099=>"000101010",
61100=>"100001000",
61101=>"001100010",
61102=>"111001011",
61103=>"001010001",
61104=>"100001111",
61105=>"111001101",
61106=>"000011111",
61107=>"000000011",
61108=>"111000000",
61109=>"010110001",
61110=>"101000000",
61111=>"111110100",
61112=>"110011010",
61113=>"111111010",
61114=>"010001000",
61115=>"000101111",
61116=>"111000000",
61117=>"000111111",
61118=>"100101101",
61119=>"111000000",
61120=>"010001011",
61121=>"110000000",
61122=>"110111000",
61123=>"111000000",
61124=>"000000000",
61125=>"011001000",
61126=>"111010111",
61127=>"100111111",
61128=>"000000000",
61129=>"100000000",
61130=>"111100000",
61131=>"001001111",
61132=>"011000000",
61133=>"001000001",
61134=>"010100100",
61135=>"000110010",
61136=>"010000110",
61137=>"110001011",
61138=>"001100000",
61139=>"000001000",
61140=>"101000111",
61141=>"011001000",
61142=>"001001011",
61143=>"111111001",
61144=>"011000111",
61145=>"000010000",
61146=>"000010111",
61147=>"100000010",
61148=>"010000000",
61149=>"111111100",
61150=>"111000100",
61151=>"111111001",
61152=>"000000000",
61153=>"101101010",
61154=>"000101111",
61155=>"011011111",
61156=>"010000000",
61157=>"010111111",
61158=>"000000111",
61159=>"010011110",
61160=>"010111101",
61161=>"000000000",
61162=>"111110100",
61163=>"100101010",
61164=>"100111111",
61165=>"111111000",
61166=>"001000000",
61167=>"100000000",
61168=>"001111111",
61169=>"101101000",
61170=>"111000010",
61171=>"111000000",
61172=>"111000010",
61173=>"011001100",
61174=>"111100000",
61175=>"111000000",
61176=>"000010111",
61177=>"010111111",
61178=>"111000100",
61179=>"111111000",
61180=>"011000100",
61181=>"100000000",
61182=>"011001000",
61183=>"111011011",
61184=>"001101010",
61185=>"110000000",
61186=>"111010010",
61187=>"101101111",
61188=>"000111110",
61189=>"001001100",
61190=>"111110000",
61191=>"110001111",
61192=>"110011000",
61193=>"110110011",
61194=>"001101010",
61195=>"000001000",
61196=>"101000000",
61197=>"100111000",
61198=>"011000010",
61199=>"010110111",
61200=>"000001101",
61201=>"000010111",
61202=>"000000001",
61203=>"001001000",
61204=>"100000000",
61205=>"110110000",
61206=>"111011001",
61207=>"000000110",
61208=>"111101101",
61209=>"001011011",
61210=>"111111000",
61211=>"111111000",
61212=>"000000111",
61213=>"111111000",
61214=>"111111111",
61215=>"111010000",
61216=>"111101111",
61217=>"100100000",
61218=>"000111111",
61219=>"010010111",
61220=>"010110000",
61221=>"000000010",
61222=>"111111000",
61223=>"000010111",
61224=>"001000000",
61225=>"000111100",
61226=>"000000111",
61227=>"011111001",
61228=>"111100110",
61229=>"101001101",
61230=>"000010111",
61231=>"111010000",
61232=>"000111010",
61233=>"111111000",
61234=>"000010111",
61235=>"001111111",
61236=>"111111010",
61237=>"000000000",
61238=>"111000000",
61239=>"010011010",
61240=>"000000111",
61241=>"111100000",
61242=>"100100101",
61243=>"000001000",
61244=>"100000000",
61245=>"101111111",
61246=>"110000000",
61247=>"000000000",
61248=>"111111111",
61249=>"110111111",
61250=>"100100110",
61251=>"001000000",
61252=>"010100010",
61253=>"001011101",
61254=>"000000000",
61255=>"111111101",
61256=>"000000000",
61257=>"111111000",
61258=>"111111111",
61259=>"000000100",
61260=>"011110010",
61261=>"111000000",
61262=>"110101100",
61263=>"011010000",
61264=>"111111010",
61265=>"000111111",
61266=>"111111111",
61267=>"111010010",
61268=>"111000000",
61269=>"000000001",
61270=>"011111000",
61271=>"000010010",
61272=>"111111111",
61273=>"001011001",
61274=>"111111000",
61275=>"011111111",
61276=>"111000111",
61277=>"001001001",
61278=>"010010000",
61279=>"111000000",
61280=>"111111011",
61281=>"000111000",
61282=>"001000000",
61283=>"111111000",
61284=>"110100000",
61285=>"111000001",
61286=>"111101111",
61287=>"111111000",
61288=>"101000001",
61289=>"000000111",
61290=>"101111111",
61291=>"000010000",
61292=>"110101000",
61293=>"000000000",
61294=>"000010010",
61295=>"111111000",
61296=>"111111000",
61297=>"000101111",
61298=>"111001000",
61299=>"000010010",
61300=>"001000111",
61301=>"001000111",
61302=>"111101000",
61303=>"000111011",
61304=>"000010000",
61305=>"100000110",
61306=>"000111000",
61307=>"111111111",
61308=>"000000000",
61309=>"100100000",
61310=>"001000010",
61311=>"110001000",
61312=>"111111010",
61313=>"011111110",
61314=>"010001000",
61315=>"011101111",
61316=>"010111110",
61317=>"000000100",
61318=>"001000000",
61319=>"110000000",
61320=>"111011001",
61321=>"000111000",
61322=>"000000000",
61323=>"100111011",
61324=>"111011110",
61325=>"010000000",
61326=>"111001101",
61327=>"011001011",
61328=>"110111101",
61329=>"111011000",
61330=>"000000111",
61331=>"110000000",
61332=>"111111000",
61333=>"000000010",
61334=>"111001000",
61335=>"001111001",
61336=>"111111111",
61337=>"000000111",
61338=>"110110000",
61339=>"111111001",
61340=>"010111111",
61341=>"001000111",
61342=>"100111111",
61343=>"001100110",
61344=>"001000000",
61345=>"110111111",
61346=>"111001000",
61347=>"111111110",
61348=>"001000000",
61349=>"111011000",
61350=>"000111011",
61351=>"001000000",
61352=>"000000111",
61353=>"110111101",
61354=>"111111000",
61355=>"001000000",
61356=>"110000000",
61357=>"010111110",
61358=>"110100100",
61359=>"110010000",
61360=>"111111100",
61361=>"011000000",
61362=>"101001100",
61363=>"101101110",
61364=>"110100100",
61365=>"001000000",
61366=>"011000001",
61367=>"001111111",
61368=>"011000000",
61369=>"010001000",
61370=>"110111111",
61371=>"010011010",
61372=>"001101110",
61373=>"100000000",
61374=>"011101000",
61375=>"001011111",
61376=>"111010010",
61377=>"101111010",
61378=>"111000001",
61379=>"110000100",
61380=>"000000111",
61381=>"100101001",
61382=>"110110111",
61383=>"111111000",
61384=>"000000000",
61385=>"111111000",
61386=>"111111001",
61387=>"111001111",
61388=>"111010000",
61389=>"111000000",
61390=>"111000000",
61391=>"111011000",
61392=>"111111111",
61393=>"100011001",
61394=>"111111001",
61395=>"111111000",
61396=>"111110000",
61397=>"111000000",
61398=>"010111000",
61399=>"000000000",
61400=>"011000000",
61401=>"110111010",
61402=>"110111110",
61403=>"000000111",
61404=>"111100000",
61405=>"010110111",
61406=>"010011111",
61407=>"000000000",
61408=>"010010000",
61409=>"111111111",
61410=>"100000000",
61411=>"100111000",
61412=>"000000000",
61413=>"001001000",
61414=>"000000001",
61415=>"011111010",
61416=>"111111111",
61417=>"011000100",
61418=>"101100000",
61419=>"111111000",
61420=>"110111111",
61421=>"000000000",
61422=>"000111111",
61423=>"011001011",
61424=>"000000000",
61425=>"001110100",
61426=>"000010010",
61427=>"111111100",
61428=>"101111001",
61429=>"111111001",
61430=>"110000000",
61431=>"100111000",
61432=>"000000110",
61433=>"001000000",
61434=>"101111000",
61435=>"111010000",
61436=>"001000000",
61437=>"000000000",
61438=>"111110000",
61439=>"000000000",
61440=>"011011011",
61441=>"000011110",
61442=>"010000111",
61443=>"000001000",
61444=>"000000100",
61445=>"110011000",
61446=>"000100000",
61447=>"100110110",
61448=>"111111000",
61449=>"110000000",
61450=>"100000000",
61451=>"111010011",
61452=>"000000000",
61453=>"000101111",
61454=>"111001000",
61455=>"000001101",
61456=>"000110010",
61457=>"110000000",
61458=>"000001101",
61459=>"010110111",
61460=>"110110100",
61461=>"111010110",
61462=>"001100100",
61463=>"000011011",
61464=>"010000000",
61465=>"110001000",
61466=>"111110000",
61467=>"101010000",
61468=>"110111010",
61469=>"000111111",
61470=>"010101000",
61471=>"001000111",
61472=>"011001001",
61473=>"110111000",
61474=>"000010111",
61475=>"111111001",
61476=>"000000000",
61477=>"111110110",
61478=>"101010000",
61479=>"111111101",
61480=>"011010111",
61481=>"110111111",
61482=>"010110000",
61483=>"010000111",
61484=>"111011110",
61485=>"000111111",
61486=>"000011101",
61487=>"000100110",
61488=>"000010010",
61489=>"100011111",
61490=>"101000001",
61491=>"111111000",
61492=>"000000010",
61493=>"111010000",
61494=>"110010000",
61495=>"001011000",
61496=>"000111101",
61497=>"101001000",
61498=>"000101101",
61499=>"000000110",
61500=>"000011111",
61501=>"101111111",
61502=>"000000000",
61503=>"000100111",
61504=>"111001000",
61505=>"111000100",
61506=>"111111111",
61507=>"001000011",
61508=>"010011011",
61509=>"000010010",
61510=>"110110001",
61511=>"110000111",
61512=>"000011111",
61513=>"010011000",
61514=>"000110111",
61515=>"011101000",
61516=>"000000000",
61517=>"011000000",
61518=>"001111111",
61519=>"110111000",
61520=>"111000110",
61521=>"010010011",
61522=>"111111110",
61523=>"001100001",
61524=>"110110110",
61525=>"001101100",
61526=>"000000011",
61527=>"111010001",
61528=>"000111110",
61529=>"000111111",
61530=>"101000011",
61531=>"100100101",
61532=>"010101000",
61533=>"000001111",
61534=>"000010011",
61535=>"000100100",
61536=>"111110000",
61537=>"101101011",
61538=>"110000001",
61539=>"000110110",
61540=>"101000001",
61541=>"001001101",
61542=>"110100000",
61543=>"111110110",
61544=>"000111110",
61545=>"000101101",
61546=>"010110111",
61547=>"110000000",
61548=>"000111110",
61549=>"110010000",
61550=>"010110000",
61551=>"010111000",
61552=>"001010101",
61553=>"000101001",
61554=>"011000000",
61555=>"010010001",
61556=>"111111000",
61557=>"000010111",
61558=>"111111101",
61559=>"111000001",
61560=>"010110001",
61561=>"010000111",
61562=>"101110000",
61563=>"000111111",
61564=>"001001010",
61565=>"100000100",
61566=>"100000000",
61567=>"101000111",
61568=>"000111000",
61569=>"001000011",
61570=>"110000101",
61571=>"000100111",
61572=>"111110010",
61573=>"101001000",
61574=>"011000111",
61575=>"011001001",
61576=>"000001110",
61577=>"111111110",
61578=>"000010010",
61579=>"010000100",
61580=>"111000111",
61581=>"100001001",
61582=>"000000000",
61583=>"000000001",
61584=>"000000100",
61585=>"101101001",
61586=>"100001110",
61587=>"001000000",
61588=>"000101100",
61589=>"111111000",
61590=>"111111000",
61591=>"100001000",
61592=>"011000111",
61593=>"010110000",
61594=>"110000111",
61595=>"000000000",
61596=>"110010000",
61597=>"000011010",
61598=>"111101001",
61599=>"010000001",
61600=>"001101011",
61601=>"111111000",
61602=>"000000001",
61603=>"111110101",
61604=>"010011000",
61605=>"000001110",
61606=>"100111011",
61607=>"111111000",
61608=>"000110110",
61609=>"000111110",
61610=>"000000111",
61611=>"110010110",
61612=>"110110110",
61613=>"111000101",
61614=>"111100110",
61615=>"110111001",
61616=>"000000001",
61617=>"100100010",
61618=>"001101111",
61619=>"011100101",
61620=>"100101011",
61621=>"010110011",
61622=>"010010111",
61623=>"011111101",
61624=>"001100111",
61625=>"000100001",
61626=>"010000011",
61627=>"010111111",
61628=>"010010111",
61629=>"100000111",
61630=>"001001110",
61631=>"000000010",
61632=>"010000000",
61633=>"111001000",
61634=>"110111110",
61635=>"001100111",
61636=>"101000000",
61637=>"011001111",
61638=>"111111010",
61639=>"111001000",
61640=>"000000100",
61641=>"000000010",
61642=>"000010111",
61643=>"000000000",
61644=>"111111000",
61645=>"101101000",
61646=>"111000111",
61647=>"000111000",
61648=>"010010111",
61649=>"001001110",
61650=>"010101011",
61651=>"000000001",
61652=>"001100000",
61653=>"000000110",
61654=>"000110110",
61655=>"111111110",
61656=>"000000000",
61657=>"011111110",
61658=>"000101101",
61659=>"000000001",
61660=>"000111110",
61661=>"110111110",
61662=>"000110111",
61663=>"010101000",
61664=>"111000000",
61665=>"111111010",
61666=>"000000010",
61667=>"100101011",
61668=>"000000001",
61669=>"000000010",
61670=>"111001000",
61671=>"111110111",
61672=>"111111000",
61673=>"000110101",
61674=>"000000000",
61675=>"000000011",
61676=>"000001001",
61677=>"001000111",
61678=>"000000001",
61679=>"000000000",
61680=>"010010111",
61681=>"110000100",
61682=>"100011011",
61683=>"001011110",
61684=>"100101001",
61685=>"001000110",
61686=>"000000111",
61687=>"000000110",
61688=>"110001001",
61689=>"111111000",
61690=>"000111111",
61691=>"111001110",
61692=>"001001101",
61693=>"000010111",
61694=>"000001010",
61695=>"011110111",
61696=>"001001100",
61697=>"000000000",
61698=>"001001001",
61699=>"001000001",
61700=>"100000100",
61701=>"111111111",
61702=>"101001101",
61703=>"001101000",
61704=>"000100000",
61705=>"000110110",
61706=>"100110010",
61707=>"110011000",
61708=>"001001111",
61709=>"011111100",
61710=>"101111010",
61711=>"101111000",
61712=>"110010000",
61713=>"000010000",
61714=>"000110110",
61715=>"101001011",
61716=>"000011111",
61717=>"000111110",
61718=>"001001111",
61719=>"001001111",
61720=>"000000001",
61721=>"110001010",
61722=>"110100111",
61723=>"110110010",
61724=>"001000000",
61725=>"001001111",
61726=>"111001010",
61727=>"000000111",
61728=>"011110111",
61729=>"001001111",
61730=>"111101001",
61731=>"001101111",
61732=>"011001000",
61733=>"111111011",
61734=>"000011010",
61735=>"001111001",
61736=>"110011011",
61737=>"100110000",
61738=>"110111000",
61739=>"001000110",
61740=>"110111110",
61741=>"000000111",
61742=>"111111111",
61743=>"010000000",
61744=>"000000111",
61745=>"101000000",
61746=>"110001000",
61747=>"101110111",
61748=>"110110001",
61749=>"011110000",
61750=>"010110001",
61751=>"110000000",
61752=>"110001111",
61753=>"100000000",
61754=>"000000000",
61755=>"000101111",
61756=>"111111100",
61757=>"001001011",
61758=>"000001111",
61759=>"110110000",
61760=>"100100101",
61761=>"001000000",
61762=>"000111011",
61763=>"110110000",
61764=>"001001111",
61765=>"100110000",
61766=>"000111000",
61767=>"001001111",
61768=>"110111111",
61769=>"110010111",
61770=>"101000000",
61771=>"000000110",
61772=>"111111000",
61773=>"111000000",
61774=>"011001000",
61775=>"111000001",
61776=>"001001000",
61777=>"110111111",
61778=>"001110110",
61779=>"111001000",
61780=>"001001000",
61781=>"111111110",
61782=>"001001110",
61783=>"110111111",
61784=>"000000010",
61785=>"100101000",
61786=>"001110011",
61787=>"101101100",
61788=>"110000111",
61789=>"100000100",
61790=>"110110000",
61791=>"110110000",
61792=>"010000000",
61793=>"110110111",
61794=>"000000111",
61795=>"010100110",
61796=>"111001011",
61797=>"111101110",
61798=>"110110011",
61799=>"110010000",
61800=>"000110100",
61801=>"111111010",
61802=>"110110000",
61803=>"100100010",
61804=>"010010011",
61805=>"110110000",
61806=>"000011011",
61807=>"111011111",
61808=>"100000000",
61809=>"110110111",
61810=>"101011000",
61811=>"001000111",
61812=>"111000010",
61813=>"000000000",
61814=>"100010110",
61815=>"110111001",
61816=>"001111000",
61817=>"001001110",
61818=>"000001111",
61819=>"111111111",
61820=>"000110011",
61821=>"000000000",
61822=>"000000101",
61823=>"110000000",
61824=>"101010000",
61825=>"111000001",
61826=>"110011000",
61827=>"001000111",
61828=>"111000000",
61829=>"000110111",
61830=>"110111010",
61831=>"100110100",
61832=>"000001000",
61833=>"001000100",
61834=>"110010011",
61835=>"000110111",
61836=>"110110000",
61837=>"001111011",
61838=>"000111110",
61839=>"000000000",
61840=>"011001001",
61841=>"001101010",
61842=>"000001111",
61843=>"010000000",
61844=>"001111111",
61845=>"110110001",
61846=>"110111111",
61847=>"000011100",
61848=>"110111001",
61849=>"110110111",
61850=>"000000110",
61851=>"000000001",
61852=>"000000101",
61853=>"010110000",
61854=>"000110111",
61855=>"000000111",
61856=>"111100110",
61857=>"110110100",
61858=>"111111111",
61859=>"011001100",
61860=>"111011010",
61861=>"000011001",
61862=>"001111110",
61863=>"001111000",
61864=>"110100010",
61865=>"100111111",
61866=>"001001001",
61867=>"000000000",
61868=>"101000111",
61869=>"000000000",
61870=>"011001101",
61871=>"000011111",
61872=>"000000000",
61873=>"111001111",
61874=>"111000001",
61875=>"100100000",
61876=>"111111000",
61877=>"000100110",
61878=>"100001001",
61879=>"101111100",
61880=>"111110111",
61881=>"010110111",
61882=>"110110101",
61883=>"110010010",
61884=>"111010010",
61885=>"110111111",
61886=>"011001000",
61887=>"001000000",
61888=>"000000111",
61889=>"001000000",
61890=>"000111111",
61891=>"011001000",
61892=>"001100000",
61893=>"111000111",
61894=>"110111111",
61895=>"010010110",
61896=>"010111101",
61897=>"010011000",
61898=>"000000001",
61899=>"010011001",
61900=>"010111000",
61901=>"100111011",
61902=>"000000001",
61903=>"111011110",
61904=>"101101111",
61905=>"100100011",
61906=>"000011000",
61907=>"000000000",
61908=>"001000001",
61909=>"000000111",
61910=>"000100010",
61911=>"001000111",
61912=>"001111111",
61913=>"000000110",
61914=>"111001011",
61915=>"001000111",
61916=>"001001110",
61917=>"111111100",
61918=>"000000011",
61919=>"110111001",
61920=>"111001010",
61921=>"001000111",
61922=>"101111000",
61923=>"111100011",
61924=>"000000111",
61925=>"111001111",
61926=>"111011111",
61927=>"001001111",
61928=>"100110111",
61929=>"101111111",
61930=>"011110000",
61931=>"001001111",
61932=>"000000010",
61933=>"010110000",
61934=>"000000001",
61935=>"111010110",
61936=>"001111111",
61937=>"100000110",
61938=>"111011010",
61939=>"011011000",
61940=>"101001111",
61941=>"001001111",
61942=>"100000001",
61943=>"001001111",
61944=>"000001000",
61945=>"001000111",
61946=>"110000101",
61947=>"000111111",
61948=>"000110000",
61949=>"111000010",
61950=>"000000000",
61951=>"000000001",
61952=>"110111011",
61953=>"011010001",
61954=>"001000111",
61955=>"000000000",
61956=>"110100100",
61957=>"111111101",
61958=>"111101111",
61959=>"000111111",
61960=>"000010000",
61961=>"101101010",
61962=>"001001101",
61963=>"000000101",
61964=>"010000111",
61965=>"000000010",
61966=>"110100000",
61967=>"001111111",
61968=>"111100110",
61969=>"000000010",
61970=>"111010101",
61971=>"111101000",
61972=>"001101010",
61973=>"000111111",
61974=>"111111100",
61975=>"111101100",
61976=>"000001000",
61977=>"001000111",
61978=>"101101110",
61979=>"000000110",
61980=>"100110111",
61981=>"000001010",
61982=>"111111100",
61983=>"011000100",
61984=>"111111010",
61985=>"111111010",
61986=>"011111001",
61987=>"010111100",
61988=>"011101100",
61989=>"000010111",
61990=>"010000110",
61991=>"111001110",
61992=>"000000110",
61993=>"000100010",
61994=>"000000100",
61995=>"001000000",
61996=>"010010001",
61997=>"100101000",
61998=>"001111111",
61999=>"011001000",
62000=>"110101000",
62001=>"100110110",
62002=>"000111111",
62003=>"111111011",
62004=>"000000111",
62005=>"000001010",
62006=>"001000101",
62007=>"000111111",
62008=>"000001100",
62009=>"000000101",
62010=>"001101111",
62011=>"001001011",
62012=>"100001011",
62013=>"110111000",
62014=>"111111111",
62015=>"000100100",
62016=>"000111111",
62017=>"001111111",
62018=>"111111111",
62019=>"101101100",
62020=>"010110111",
62021=>"101000101",
62022=>"000111111",
62023=>"110100111",
62024=>"100110101",
62025=>"111001110",
62026=>"111001000",
62027=>"010100000",
62028=>"110111111",
62029=>"010000110",
62030=>"111011011",
62031=>"100010000",
62032=>"111111000",
62033=>"010110010",
62034=>"001111111",
62035=>"000001100",
62036=>"101001111",
62037=>"011111111",
62038=>"111011011",
62039=>"100100111",
62040=>"000000000",
62041=>"100110100",
62042=>"011000000",
62043=>"100100100",
62044=>"000001001",
62045=>"000000000",
62046=>"110111111",
62047=>"001000001",
62048=>"010111000",
62049=>"111001000",
62050=>"111101100",
62051=>"011001000",
62052=>"000000000",
62053=>"110110010",
62054=>"111001111",
62055=>"110100111",
62056=>"000101111",
62057=>"111101001",
62058=>"000000000",
62059=>"111111111",
62060=>"010001000",
62061=>"000111111",
62062=>"000000001",
62063=>"000000111",
62064=>"111011001",
62065=>"000000100",
62066=>"100000011",
62067=>"000001000",
62068=>"101010110",
62069=>"001001111",
62070=>"000000001",
62071=>"100010000",
62072=>"000000111",
62073=>"111111000",
62074=>"000000000",
62075=>"101101111",
62076=>"000001001",
62077=>"110100010",
62078=>"000000110",
62079=>"111000000",
62080=>"000111111",
62081=>"011011010",
62082=>"101101101",
62083=>"000010111",
62084=>"101101000",
62085=>"000000001",
62086=>"000000111",
62087=>"111100100",
62088=>"110100100",
62089=>"111111111",
62090=>"101101011",
62091=>"011000000",
62092=>"000000000",
62093=>"010110010",
62094=>"000000000",
62095=>"000000000",
62096=>"110100000",
62097=>"111111000",
62098=>"110011000",
62099=>"111100100",
62100=>"000000000",
62101=>"000001000",
62102=>"010111111",
62103=>"001011011",
62104=>"000110111",
62105=>"111111001",
62106=>"100111111",
62107=>"101100010",
62108=>"000010110",
62109=>"110111111",
62110=>"000000000",
62111=>"000000010",
62112=>"010110101",
62113=>"001110110",
62114=>"010000100",
62115=>"000001001",
62116=>"000000001",
62117=>"011111011",
62118=>"000110000",
62119=>"000000000",
62120=>"000001011",
62121=>"000010000",
62122=>"001101010",
62123=>"010000000",
62124=>"111000110",
62125=>"101111111",
62126=>"110110000",
62127=>"111111011",
62128=>"001100000",
62129=>"000000001",
62130=>"111000101",
62131=>"110000000",
62132=>"011100000",
62133=>"000000000",
62134=>"100000000",
62135=>"000000000",
62136=>"000000100",
62137=>"000011011",
62138=>"000100111",
62139=>"110111000",
62140=>"010111111",
62141=>"010110010",
62142=>"001011001",
62143=>"001111111",
62144=>"101000001",
62145=>"101000111",
62146=>"000111111",
62147=>"010000110",
62148=>"011101011",
62149=>"111000100",
62150=>"110111100",
62151=>"001000110",
62152=>"111011110",
62153=>"010000000",
62154=>"001000000",
62155=>"011111000",
62156=>"101101000",
62157=>"000100101",
62158=>"000000001",
62159=>"111111110",
62160=>"001000111",
62161=>"110110010",
62162=>"001000000",
62163=>"011111111",
62164=>"011010110",
62165=>"110110000",
62166=>"000000111",
62167=>"000000101",
62168=>"111000000",
62169=>"010101000",
62170=>"000011111",
62171=>"001001111",
62172=>"111011001",
62173=>"110010000",
62174=>"000000001",
62175=>"000000101",
62176=>"000000101",
62177=>"001000000",
62178=>"101000000",
62179=>"011011000",
62180=>"000000000",
62181=>"101000000",
62182=>"000000111",
62183=>"010111010",
62184=>"001100101",
62185=>"010011111",
62186=>"101101110",
62187=>"000000000",
62188=>"000001000",
62189=>"111010010",
62190=>"000000100",
62191=>"111111001",
62192=>"111000011",
62193=>"110100011",
62194=>"001111110",
62195=>"010111001",
62196=>"000110010",
62197=>"101000000",
62198=>"101111111",
62199=>"110100110",
62200=>"000000010",
62201=>"001010110",
62202=>"010000101",
62203=>"000000000",
62204=>"111111010",
62205=>"010101101",
62206=>"000011011",
62207=>"000010000",
62208=>"100111100",
62209=>"111000000",
62210=>"101101100",
62211=>"000001000",
62212=>"100111111",
62213=>"001000101",
62214=>"000111011",
62215=>"000000000",
62216=>"010111000",
62217=>"101101000",
62218=>"101000000",
62219=>"000000000",
62220=>"111100000",
62221=>"110111111",
62222=>"000100000",
62223=>"011000111",
62224=>"101000000",
62225=>"100101101",
62226=>"100001101",
62227=>"111100000",
62228=>"110010000",
62229=>"111101111",
62230=>"100111110",
62231=>"101101101",
62232=>"111001100",
62233=>"111010100",
62234=>"111101000",
62235=>"101101001",
62236=>"101100111",
62237=>"100000111",
62238=>"101101111",
62239=>"000111111",
62240=>"010100000",
62241=>"010010000",
62242=>"100101011",
62243=>"000000010",
62244=>"000001111",
62245=>"001100111",
62246=>"101101000",
62247=>"001000101",
62248=>"001001100",
62249=>"011010000",
62250=>"111000001",
62251=>"100100101",
62252=>"110110111",
62253=>"000100011",
62254=>"111110101",
62255=>"101001001",
62256=>"111111110",
62257=>"001000111",
62258=>"101100110",
62259=>"101001010",
62260=>"111000101",
62261=>"000111111",
62262=>"111100001",
62263=>"001111111",
62264=>"010010111",
62265=>"000010011",
62266=>"001101101",
62267=>"101101011",
62268=>"000011111",
62269=>"111111000",
62270=>"000000000",
62271=>"000100110",
62272=>"001000000",
62273=>"000000110",
62274=>"011111111",
62275=>"000000100",
62276=>"101100010",
62277=>"111010100",
62278=>"101101111",
62279=>"000010000",
62280=>"000011101",
62281=>"111101111",
62282=>"000000101",
62283=>"000111101",
62284=>"110100111",
62285=>"000100101",
62286=>"000000101",
62287=>"000101110",
62288=>"000100100",
62289=>"111111111",
62290=>"010111010",
62291=>"000101101",
62292=>"111110000",
62293=>"000110100",
62294=>"000001111",
62295=>"000101000",
62296=>"001001110",
62297=>"000001000",
62298=>"000100011",
62299=>"000001100",
62300=>"101000010",
62301=>"100110101",
62302=>"010010110",
62303=>"000000001",
62304=>"001000100",
62305=>"100101000",
62306=>"101000000",
62307=>"001011101",
62308=>"000000001",
62309=>"000111001",
62310=>"110011010",
62311=>"000010010",
62312=>"000000010",
62313=>"111100101",
62314=>"001001011",
62315=>"110111001",
62316=>"000000000",
62317=>"111001010",
62318=>"000000000",
62319=>"010110100",
62320=>"000001111",
62321=>"000000000",
62322=>"101001100",
62323=>"000101110",
62324=>"110000000",
62325=>"101001101",
62326=>"001010101",
62327=>"010010111",
62328=>"101000000",
62329=>"011000100",
62330=>"000001101",
62331=>"110110111",
62332=>"001001000",
62333=>"000101011",
62334=>"001100110",
62335=>"100000000",
62336=>"111000000",
62337=>"010010010",
62338=>"100000100",
62339=>"000110000",
62340=>"000000011",
62341=>"011110010",
62342=>"000000111",
62343=>"100100000",
62344=>"100110101",
62345=>"101011010",
62346=>"000100111",
62347=>"110111001",
62348=>"000011010",
62349=>"001100101",
62350=>"000010101",
62351=>"001001101",
62352=>"010111110",
62353=>"001010101",
62354=>"111101110",
62355=>"000000111",
62356=>"001100010",
62357=>"101000010",
62358=>"110010110",
62359=>"100100101",
62360=>"110000000",
62361=>"000000110",
62362=>"101100001",
62363=>"101101111",
62364=>"111101010",
62365=>"111000111",
62366=>"001000010",
62367=>"010000111",
62368=>"000000111",
62369=>"101111111",
62370=>"111111111",
62371=>"101100000",
62372=>"100001000",
62373=>"010101111",
62374=>"011111000",
62375=>"111011111",
62376=>"111001110",
62377=>"000001010",
62378=>"111001001",
62379=>"101000000",
62380=>"001000000",
62381=>"000000010",
62382=>"001110110",
62383=>"101110110",
62384=>"000000000",
62385=>"100000010",
62386=>"000110101",
62387=>"001001001",
62388=>"111111000",
62389=>"000000001",
62390=>"100000100",
62391=>"011000000",
62392=>"100110111",
62393=>"001000000",
62394=>"111110101",
62395=>"101101111",
62396=>"010010000",
62397=>"001010000",
62398=>"000000010",
62399=>"001111011",
62400=>"000000011",
62401=>"101100100",
62402=>"111101101",
62403=>"100001011",
62404=>"010010000",
62405=>"100000100",
62406=>"000100110",
62407=>"000100100",
62408=>"011010111",
62409=>"000011110",
62410=>"011110000",
62411=>"000010010",
62412=>"100111111",
62413=>"110100000",
62414=>"111111000",
62415=>"010010001",
62416=>"100101011",
62417=>"011111111",
62418=>"101110001",
62419=>"010111111",
62420=>"001000000",
62421=>"010011001",
62422=>"110000010",
62423=>"010000000",
62424=>"000101111",
62425=>"111000010",
62426=>"011010001",
62427=>"111101101",
62428=>"100010000",
62429=>"011000110",
62430=>"111111101",
62431=>"111111010",
62432=>"000010110",
62433=>"101101111",
62434=>"101110110",
62435=>"100001111",
62436=>"111101100",
62437=>"111111111",
62438=>"110111111",
62439=>"000011011",
62440=>"110111101",
62441=>"110111101",
62442=>"111000000",
62443=>"011011000",
62444=>"010010000",
62445=>"000000010",
62446=>"000000100",
62447=>"100101101",
62448=>"010110000",
62449=>"001001000",
62450=>"000000111",
62451=>"110110100",
62452=>"010010001",
62453=>"111100010",
62454=>"100101000",
62455=>"101100101",
62456=>"000000000",
62457=>"010101101",
62458=>"111110100",
62459=>"000011000",
62460=>"001111111",
62461=>"000000011",
62462=>"001001011",
62463=>"111001000",
62464=>"011011001",
62465=>"010001001",
62466=>"001000001",
62467=>"000000001",
62468=>"011011011",
62469=>"110110101",
62470=>"000000000",
62471=>"011000001",
62472=>"011011110",
62473=>"000000000",
62474=>"100000000",
62475=>"000111011",
62476=>"101000111",
62477=>"000000110",
62478=>"001111001",
62479=>"000111110",
62480=>"000000111",
62481=>"011000011",
62482=>"000010110",
62483=>"000100110",
62484=>"111110011",
62485=>"100000000",
62486=>"110100100",
62487=>"111000111",
62488=>"001101100",
62489=>"100000000",
62490=>"101000100",
62491=>"111111000",
62492=>"101000000",
62493=>"000100111",
62494=>"111111100",
62495=>"000000011",
62496=>"000000000",
62497=>"110111100",
62498=>"001001000",
62499=>"000000000",
62500=>"011001100",
62501=>"110110010",
62502=>"011010010",
62503=>"010011000",
62504=>"111011000",
62505=>"001111111",
62506=>"101000011",
62507=>"110110000",
62508=>"001011011",
62509=>"100111111",
62510=>"000100111",
62511=>"000000111",
62512=>"000000111",
62513=>"000001111",
62514=>"101101011",
62515=>"111000000",
62516=>"000000000",
62517=>"010110111",
62518=>"110000001",
62519=>"000000000",
62520=>"011111111",
62521=>"001000000",
62522=>"100000101",
62523=>"000000100",
62524=>"110111011",
62525=>"111111100",
62526=>"000000000",
62527=>"001111000",
62528=>"000000001",
62529=>"111110111",
62530=>"000111101",
62531=>"011010000",
62532=>"011111100",
62533=>"000001101",
62534=>"111000110",
62535=>"101111010",
62536=>"000011010",
62537=>"111111010",
62538=>"111001101",
62539=>"111000101",
62540=>"000000000",
62541=>"111011001",
62542=>"010011110",
62543=>"101000111",
62544=>"000101111",
62545=>"110010001",
62546=>"111111101",
62547=>"111001100",
62548=>"000111000",
62549=>"010011110",
62550=>"111001101",
62551=>"101101111",
62552=>"001001110",
62553=>"100110111",
62554=>"110001101",
62555=>"111110111",
62556=>"100110001",
62557=>"010000000",
62558=>"101010111",
62559=>"000001001",
62560=>"010111010",
62561=>"000101100",
62562=>"110010000",
62563=>"001000101",
62564=>"110010011",
62565=>"000000001",
62566=>"111111000",
62567=>"111000000",
62568=>"111111100",
62569=>"111111010",
62570=>"110111111",
62571=>"100000000",
62572=>"000000011",
62573=>"000000111",
62574=>"001000101",
62575=>"111101111",
62576=>"100110011",
62577=>"000111111",
62578=>"010000100",
62579=>"101111111",
62580=>"011001011",
62581=>"000000000",
62582=>"111110111",
62583=>"111111000",
62584=>"011001101",
62585=>"111111101",
62586=>"001001000",
62587=>"000000110",
62588=>"000111011",
62589=>"011100000",
62590=>"010000010",
62591=>"111010000",
62592=>"111110101",
62593=>"010000000",
62594=>"110111011",
62595=>"100000000",
62596=>"111111101",
62597=>"001000010",
62598=>"011111110",
62599=>"000100000",
62600=>"010111100",
62601=>"101000010",
62602=>"100000111",
62603=>"000000000",
62604=>"000000000",
62605=>"111001000",
62606=>"000000101",
62607=>"000000000",
62608=>"001111110",
62609=>"000110000",
62610=>"111000111",
62611=>"111101000",
62612=>"111111000",
62613=>"111010000",
62614=>"000101001",
62615=>"011111101",
62616=>"011110100",
62617=>"000010001",
62618=>"000010010",
62619=>"000000000",
62620=>"000001010",
62621=>"010111000",
62622=>"111110110",
62623=>"000000100",
62624=>"000100000",
62625=>"111111111",
62626=>"110110001",
62627=>"010000101",
62628=>"111011100",
62629=>"111001001",
62630=>"000001000",
62631=>"000110111",
62632=>"111111000",
62633=>"001101101",
62634=>"000000100",
62635=>"111101111",
62636=>"001001100",
62637=>"111111000",
62638=>"100111111",
62639=>"001100111",
62640=>"000000000",
62641=>"100101001",
62642=>"010000000",
62643=>"011000000",
62644=>"010100100",
62645=>"101000111",
62646=>"000000000",
62647=>"101110010",
62648=>"011111110",
62649=>"101101001",
62650=>"010011111",
62651=>"111111010",
62652=>"000111100",
62653=>"111111111",
62654=>"100111011",
62655=>"000101111",
62656=>"101000000",
62657=>"101000000",
62658=>"111110111",
62659=>"010000011",
62660=>"111111010",
62661=>"000000000",
62662=>"111000000",
62663=>"011110000",
62664=>"000001000",
62665=>"000000000",
62666=>"010011100",
62667=>"000000001",
62668=>"000010010",
62669=>"001101010",
62670=>"000001001",
62671=>"000101000",
62672=>"001111110",
62673=>"100100011",
62674=>"011101000",
62675=>"010111111",
62676=>"101000101",
62677=>"011000111",
62678=>"001111011",
62679=>"000111111",
62680=>"100000001",
62681=>"111000000",
62682=>"000000101",
62683=>"000000111",
62684=>"000001011",
62685=>"000111110",
62686=>"100000010",
62687=>"011010001",
62688=>"000000001",
62689=>"111101101",
62690=>"101111001",
62691=>"101101111",
62692=>"101000111",
62693=>"000011011",
62694=>"000101111",
62695=>"011001111",
62696=>"010010011",
62697=>"110101111",
62698=>"001000001",
62699=>"000000001",
62700=>"110111000",
62701=>"100101001",
62702=>"010000000",
62703=>"000001000",
62704=>"000000111",
62705=>"000000100",
62706=>"100000000",
62707=>"011001001",
62708=>"010110100",
62709=>"001000000",
62710=>"000000001",
62711=>"110000000",
62712=>"111111111",
62713=>"000001011",
62714=>"111001111",
62715=>"001001010",
62716=>"110000111",
62717=>"100101111",
62718=>"111110000",
62719=>"001000100",
62720=>"000001000",
62721=>"000100000",
62722=>"100010011",
62723=>"101111111",
62724=>"110111010",
62725=>"000001011",
62726=>"000011111",
62727=>"000111110",
62728=>"011011010",
62729=>"011010100",
62730=>"110110010",
62731=>"100111111",
62732=>"110100100",
62733=>"010000001",
62734=>"000000000",
62735=>"100001000",
62736=>"110111101",
62737=>"111111001",
62738=>"111100110",
62739=>"100000110",
62740=>"100000011",
62741=>"011011101",
62742=>"110100100",
62743=>"110111111",
62744=>"100000111",
62745=>"100111101",
62746=>"000000111",
62747=>"011011011",
62748=>"111011101",
62749=>"000000100",
62750=>"110111011",
62751=>"000100001",
62752=>"110100000",
62753=>"000101111",
62754=>"000001010",
62755=>"011101000",
62756=>"100110011",
62757=>"111111111",
62758=>"100010100",
62759=>"111010000",
62760=>"000001001",
62761=>"111111011",
62762=>"110110000",
62763=>"100100100",
62764=>"000100100",
62765=>"101100000",
62766=>"111110111",
62767=>"000000110",
62768=>"111110010",
62769=>"110100100",
62770=>"011111000",
62771=>"000011001",
62772=>"100100100",
62773=>"110110000",
62774=>"011000001",
62775=>"000000001",
62776=>"101111010",
62777=>"000000011",
62778=>"000000001",
62779=>"111110110",
62780=>"010000111",
62781=>"000100001",
62782=>"010000000",
62783=>"100000000",
62784=>"100111110",
62785=>"110000000",
62786=>"100100001",
62787=>"000110100",
62788=>"111000001",
62789=>"100111011",
62790=>"001001010",
62791=>"100000000",
62792=>"011011000",
62793=>"011101111",
62794=>"100000111",
62795=>"111101111",
62796=>"000001101",
62797=>"010110111",
62798=>"000100100",
62799=>"111111101",
62800=>"100000101",
62801=>"100110111",
62802=>"111011011",
62803=>"101100100",
62804=>"100110010",
62805=>"110110111",
62806=>"000100100",
62807=>"101011011",
62808=>"001001111",
62809=>"000100100",
62810=>"001001000",
62811=>"000111100",
62812=>"111111000",
62813=>"001000000",
62814=>"011111111",
62815=>"100100001",
62816=>"111000000",
62817=>"111011000",
62818=>"111011111",
62819=>"111110101",
62820=>"000100011",
62821=>"001101000",
62822=>"000000000",
62823=>"000000100",
62824=>"000001001",
62825=>"000110010",
62826=>"011111111",
62827=>"001011111",
62828=>"011110010",
62829=>"011011011",
62830=>"001100000",
62831=>"011111011",
62832=>"100100111",
62833=>"100100010",
62834=>"101110000",
62835=>"001000000",
62836=>"100111011",
62837=>"001111111",
62838=>"111011100",
62839=>"111011011",
62840=>"000010000",
62841=>"001111011",
62842=>"111000111",
62843=>"011100110",
62844=>"001100100",
62845=>"111000011",
62846=>"111011101",
62847=>"100100000",
62848=>"100011011",
62849=>"011000100",
62850=>"110011001",
62851=>"011000000",
62852=>"010000100",
62853=>"010101000",
62854=>"000000000",
62855=>"010100000",
62856=>"000100100",
62857=>"110110010",
62858=>"001001000",
62859=>"001000011",
62860=>"011011001",
62861=>"110001010",
62862=>"011001000",
62863=>"000001100",
62864=>"110110100",
62865=>"111001100",
62866=>"111000001",
62867=>"100100100",
62868=>"000101100",
62869=>"100111011",
62870=>"100100000",
62871=>"000000000",
62872=>"000001011",
62873=>"011011010",
62874=>"000101000",
62875=>"001100000",
62876=>"010010111",
62877=>"110000111",
62878=>"010010000",
62879=>"111100100",
62880=>"100100000",
62881=>"111011001",
62882=>"111100010",
62883=>"110010101",
62884=>"011011011",
62885=>"001001000",
62886=>"011111000",
62887=>"111100000",
62888=>"111111011",
62889=>"000111111",
62890=>"111000000",
62891=>"111100110",
62892=>"001111110",
62893=>"100000111",
62894=>"001000010",
62895=>"111001100",
62896=>"011100101",
62897=>"001001000",
62898=>"111100011",
62899=>"011100110",
62900=>"101101000",
62901=>"011001000",
62902=>"111011110",
62903=>"000000100",
62904=>"001011000",
62905=>"101111011",
62906=>"111001011",
62907=>"110110000",
62908=>"001101011",
62909=>"110111111",
62910=>"010000001",
62911=>"001000101",
62912=>"111011001",
62913=>"110100000",
62914=>"111101010",
62915=>"100100101",
62916=>"000000000",
62917=>"000101111",
62918=>"100111011",
62919=>"111000000",
62920=>"101000100",
62921=>"000011011",
62922=>"100010011",
62923=>"010111010",
62924=>"000111000",
62925=>"000000001",
62926=>"000011001",
62927=>"110010000",
62928=>"100001000",
62929=>"000111110",
62930=>"011000001",
62931=>"110100000",
62932=>"110111001",
62933=>"110111111",
62934=>"000100000",
62935=>"000100010",
62936=>"110100100",
62937=>"111100000",
62938=>"010100110",
62939=>"011011001",
62940=>"000100110",
62941=>"111001010",
62942=>"001110000",
62943=>"111111011",
62944=>"000111000",
62945=>"010010000",
62946=>"011001000",
62947=>"100111110",
62948=>"101001000",
62949=>"100001111",
62950=>"100110010",
62951=>"001111110",
62952=>"011101101",
62953=>"111000000",
62954=>"111001000",
62955=>"111111101",
62956=>"000011000",
62957=>"000100011",
62958=>"000011011",
62959=>"111000000",
62960=>"000111001",
62961=>"000100110",
62962=>"110000011",
62963=>"110000001",
62964=>"000110100",
62965=>"001000000",
62966=>"001011110",
62967=>"010001100",
62968=>"000111111",
62969=>"001001001",
62970=>"111111100",
62971=>"000100101",
62972=>"000101101",
62973=>"010111110",
62974=>"000111000",
62975=>"000010111",
62976=>"001001000",
62977=>"010100011",
62978=>"001001111",
62979=>"001001111",
62980=>"000000110",
62981=>"111001001",
62982=>"001001001",
62983=>"010000000",
62984=>"001001111",
62985=>"000000110",
62986=>"100101101",
62987=>"111011011",
62988=>"001001011",
62989=>"011111110",
62990=>"011001011",
62991=>"010111111",
62992=>"011011110",
62993=>"011001011",
62994=>"001000111",
62995=>"110100000",
62996=>"011001110",
62997=>"110110100",
62998=>"101111011",
62999=>"001110101",
63000=>"011001111",
63001=>"100100100",
63002=>"110011111",
63003=>"011001111",
63004=>"100100110",
63005=>"100010110",
63006=>"111111111",
63007=>"100011000",
63008=>"100111101",
63009=>"001011111",
63010=>"000110000",
63011=>"110000000",
63012=>"000100000",
63013=>"111011000",
63014=>"000000110",
63015=>"001101111",
63016=>"110110110",
63017=>"111011111",
63018=>"001100000",
63019=>"000000000",
63020=>"010000100",
63021=>"111010011",
63022=>"110110110",
63023=>"111001110",
63024=>"110111000",
63025=>"000000000",
63026=>"000110111",
63027=>"100000100",
63028=>"100110110",
63029=>"010000001",
63030=>"111001000",
63031=>"100100110",
63032=>"101000000",
63033=>"001001111",
63034=>"000000101",
63035=>"000100000",
63036=>"100110000",
63037=>"001100001",
63038=>"000000011",
63039=>"000000001",
63040=>"111011001",
63041=>"111111000",
63042=>"011001001",
63043=>"011011001",
63044=>"011011000",
63045=>"001001011",
63046=>"100110000",
63047=>"101000101",
63048=>"111011100",
63049=>"010000100",
63050=>"011011011",
63051=>"100100000",
63052=>"100001000",
63053=>"100010110",
63054=>"000001001",
63055=>"000000100",
63056=>"011000111",
63057=>"100111110",
63058=>"101011111",
63059=>"100111100",
63060=>"011000010",
63061=>"111110111",
63062=>"110110100",
63063=>"001001011",
63064=>"010000000",
63065=>"110100100",
63066=>"110111100",
63067=>"100110000",
63068=>"110110100",
63069=>"100100100",
63070=>"111111011",
63071=>"001010011",
63072=>"000100001",
63073=>"001001111",
63074=>"001001011",
63075=>"100100100",
63076=>"011011001",
63077=>"000110110",
63078=>"111110100",
63079=>"111110110",
63080=>"101101001",
63081=>"100001001",
63082=>"000111111",
63083=>"001111111",
63084=>"110010110",
63085=>"010011001",
63086=>"110110000",
63087=>"111101001",
63088=>"000100000",
63089=>"111100100",
63090=>"001000000",
63091=>"001001000",
63092=>"001001000",
63093=>"000001100",
63094=>"100001110",
63095=>"110110111",
63096=>"110111111",
63097=>"010100000",
63098=>"001100100",
63099=>"001001001",
63100=>"100100101",
63101=>"111001000",
63102=>"101111110",
63103=>"011001111",
63104=>"110111000",
63105=>"000000001",
63106=>"100100100",
63107=>"100100111",
63108=>"111011111",
63109=>"101111000",
63110=>"100100000",
63111=>"000001000",
63112=>"110010000",
63113=>"111000010",
63114=>"111111000",
63115=>"011000110",
63116=>"001111001",
63117=>"001000001",
63118=>"001001110",
63119=>"100000100",
63120=>"111100101",
63121=>"110011001",
63122=>"100111000",
63123=>"011001001",
63124=>"100000110",
63125=>"001001111",
63126=>"000100100",
63127=>"001001000",
63128=>"101101010",
63129=>"000001110",
63130=>"100110100",
63131=>"100001000",
63132=>"111000000",
63133=>"111100000",
63134=>"011100000",
63135=>"010011111",
63136=>"100001011",
63137=>"111010001",
63138=>"001001110",
63139=>"111111011",
63140=>"001011000",
63141=>"110000100",
63142=>"001000111",
63143=>"000100100",
63144=>"110000100",
63145=>"011001010",
63146=>"110010110",
63147=>"011001111",
63148=>"110111001",
63149=>"001001111",
63150=>"010011110",
63151=>"001000111",
63152=>"001111010",
63153=>"001001010",
63154=>"111001111",
63155=>"111001001",
63156=>"111111100",
63157=>"110110000",
63158=>"111110110",
63159=>"000111000",
63160=>"110100111",
63161=>"001100000",
63162=>"110010000",
63163=>"111111000",
63164=>"100010010",
63165=>"101001000",
63166=>"011011111",
63167=>"101000000",
63168=>"111100111",
63169=>"110110100",
63170=>"100101101",
63171=>"001110100",
63172=>"000110000",
63173=>"110011001",
63174=>"111001001",
63175=>"000110110",
63176=>"110100111",
63177=>"100001001",
63178=>"110110110",
63179=>"000100100",
63180=>"110100000",
63181=>"001100101",
63182=>"100110100",
63183=>"100100111",
63184=>"001011011",
63185=>"001110010",
63186=>"101000001",
63187=>"011110101",
63188=>"111100110",
63189=>"100111100",
63190=>"011001011",
63191=>"110110110",
63192=>"100110000",
63193=>"011011010",
63194=>"000000001",
63195=>"110001011",
63196=>"000101001",
63197=>"111011010",
63198=>"110110000",
63199=>"111111000",
63200=>"011001011",
63201=>"011001011",
63202=>"111011001",
63203=>"001001101",
63204=>"111001001",
63205=>"011001011",
63206=>"001001001",
63207=>"100110000",
63208=>"111011011",
63209=>"010110100",
63210=>"111111100",
63211=>"001000000",
63212=>"011001001",
63213=>"110111111",
63214=>"110100110",
63215=>"110110010",
63216=>"100000000",
63217=>"001000011",
63218=>"010001110",
63219=>"100100110",
63220=>"100111111",
63221=>"000111110",
63222=>"000100100",
63223=>"100000100",
63224=>"001110100",
63225=>"000111100",
63226=>"110001011",
63227=>"001011100",
63228=>"110110100",
63229=>"010000000",
63230=>"100111101",
63231=>"111101101",
63232=>"000000110",
63233=>"101000000",
63234=>"001000000",
63235=>"000111010",
63236=>"000000000",
63237=>"110000111",
63238=>"000011010",
63239=>"000000000",
63240=>"110010111",
63241=>"000000001",
63242=>"001011110",
63243=>"000000000",
63244=>"000111110",
63245=>"101000110",
63246=>"000010010",
63247=>"011111001",
63248=>"000000101",
63249=>"111010011",
63250=>"111111011",
63251=>"000100111",
63252=>"000000000",
63253=>"000000000",
63254=>"111111100",
63255=>"110110010",
63256=>"011000010",
63257=>"100111111",
63258=>"011000111",
63259=>"000000000",
63260=>"000000101",
63261=>"001101001",
63262=>"000000000",
63263=>"111111111",
63264=>"111000111",
63265=>"000101000",
63266=>"001100000",
63267=>"101001111",
63268=>"000100110",
63269=>"001000111",
63270=>"000010010",
63271=>"111001010",
63272=>"000000001",
63273=>"111001001",
63274=>"010111110",
63275=>"111111111",
63276=>"010101011",
63277=>"101010000",
63278=>"111111010",
63279=>"000001001",
63280=>"110111111",
63281=>"110110110",
63282=>"000101101",
63283=>"010000010",
63284=>"101000000",
63285=>"001010011",
63286=>"001110010",
63287=>"000000000",
63288=>"010111001",
63289=>"000000000",
63290=>"100111000",
63291=>"010010000",
63292=>"011000010",
63293=>"111111101",
63294=>"101001101",
63295=>"100111001",
63296=>"111010111",
63297=>"000000001",
63298=>"000111000",
63299=>"001000100",
63300=>"110110000",
63301=>"111110010",
63302=>"000000000",
63303=>"000000111",
63304=>"110010101",
63305=>"010000000",
63306=>"100001011",
63307=>"111110110",
63308=>"100101101",
63309=>"011011011",
63310=>"000001011",
63311=>"111111111",
63312=>"000000000",
63313=>"111110110",
63314=>"101000010",
63315=>"101110000",
63316=>"000000001",
63317=>"110000000",
63318=>"000001001",
63319=>"000000000",
63320=>"111111011",
63321=>"101111111",
63322=>"000010100",
63323=>"011111100",
63324=>"111111010",
63325=>"000100100",
63326=>"111000000",
63327=>"000000001",
63328=>"010000001",
63329=>"110110000",
63330=>"000000100",
63331=>"000001001",
63332=>"000111110",
63333=>"111001111",
63334=>"110010000",
63335=>"000000000",
63336=>"000011000",
63337=>"000010010",
63338=>"111000000",
63339=>"101000110",
63340=>"100100000",
63341=>"010010011",
63342=>"000000000",
63343=>"000000000",
63344=>"101111111",
63345=>"111111000",
63346=>"011110011",
63347=>"000101000",
63348=>"000000000",
63349=>"000110000",
63350=>"000111000",
63351=>"111010111",
63352=>"011111101",
63353=>"111111000",
63354=>"111100100",
63355=>"111111011",
63356=>"100010100",
63357=>"000110111",
63358=>"000000010",
63359=>"111000000",
63360=>"110111001",
63361=>"111100000",
63362=>"011011010",
63363=>"011110110",
63364=>"001101001",
63365=>"000111111",
63366=>"010010110",
63367=>"100110011",
63368=>"111111101",
63369=>"101101000",
63370=>"001111001",
63371=>"001000000",
63372=>"000000000",
63373=>"011111101",
63374=>"110110110",
63375=>"001001000",
63376=>"111111111",
63377=>"100011111",
63378=>"111001101",
63379=>"101000110",
63380=>"000110010",
63381=>"111101100",
63382=>"100010000",
63383=>"110110010",
63384=>"100101101",
63385=>"110110111",
63386=>"000110110",
63387=>"000000111",
63388=>"111000110",
63389=>"010111000",
63390=>"111000000",
63391=>"000000000",
63392=>"001011011",
63393=>"111111011",
63394=>"000000111",
63395=>"101011111",
63396=>"000110110",
63397=>"110111010",
63398=>"111001000",
63399=>"000000001",
63400=>"011010010",
63401=>"000000000",
63402=>"111111111",
63403=>"001101000",
63404=>"111111110",
63405=>"101101111",
63406=>"000101011",
63407=>"001111110",
63408=>"000000010",
63409=>"001110110",
63410=>"111111010",
63411=>"000001011",
63412=>"111111111",
63413=>"010011001",
63414=>"101011111",
63415=>"101000110",
63416=>"010010000",
63417=>"001011011",
63418=>"101000010",
63419=>"110111111",
63420=>"000100000",
63421=>"000000111",
63422=>"110110101",
63423=>"010000101",
63424=>"111111010",
63425=>"011011010",
63426=>"111111000",
63427=>"110110100",
63428=>"000001111",
63429=>"110110001",
63430=>"000000100",
63431=>"000000111",
63432=>"000000111",
63433=>"101111111",
63434=>"101000111",
63435=>"010110000",
63436=>"111010010",
63437=>"000000010",
63438=>"001101110",
63439=>"111011000",
63440=>"001000000",
63441=>"101111110",
63442=>"000001100",
63443=>"111101101",
63444=>"001111111",
63445=>"001100001",
63446=>"000000000",
63447=>"110000111",
63448=>"000000000",
63449=>"000001101",
63450=>"100110111",
63451=>"000111111",
63452=>"111001111",
63453=>"111111111",
63454=>"000000000",
63455=>"000000101",
63456=>"111111001",
63457=>"111000000",
63458=>"111010000",
63459=>"001011011",
63460=>"000000000",
63461=>"000000010",
63462=>"000000010",
63463=>"010111100",
63464=>"111000111",
63465=>"000100100",
63466=>"110010000",
63467=>"010000111",
63468=>"000001101",
63469=>"000000001",
63470=>"000111010",
63471=>"000000010",
63472=>"101101111",
63473=>"011010110",
63474=>"101111000",
63475=>"010111011",
63476=>"000001011",
63477=>"000101001",
63478=>"000100110",
63479=>"000001000",
63480=>"000110100",
63481=>"000000000",
63482=>"111111110",
63483=>"111111001",
63484=>"000010010",
63485=>"000000010",
63486=>"100111011",
63487=>"000111111",
63488=>"111110111",
63489=>"010010000",
63490=>"100000000",
63491=>"000010111",
63492=>"011111011",
63493=>"111111010",
63494=>"011110100",
63495=>"010000000",
63496=>"000111010",
63497=>"100111000",
63498=>"101111011",
63499=>"000000100",
63500=>"100000101",
63501=>"111111111",
63502=>"111101000",
63503=>"101001010",
63504=>"001001100",
63505=>"110000110",
63506=>"001000000",
63507=>"011100000",
63508=>"000100100",
63509=>"000010000",
63510=>"010110011",
63511=>"110110001",
63512=>"000001111",
63513=>"000000100",
63514=>"011011000",
63515=>"000111100",
63516=>"101100010",
63517=>"000000111",
63518=>"111010001",
63519=>"000000010",
63520=>"111111111",
63521=>"111111111",
63522=>"101000110",
63523=>"011111111",
63524=>"001011010",
63525=>"101001010",
63526=>"110110000",
63527=>"000000000",
63528=>"011111010",
63529=>"000010000",
63530=>"101111000",
63531=>"010010000",
63532=>"000011011",
63533=>"101111001",
63534=>"111111011",
63535=>"011000010",
63536=>"000000110",
63537=>"001011011",
63538=>"111011110",
63539=>"111111111",
63540=>"101110111",
63541=>"100000000",
63542=>"100000000",
63543=>"000000000",
63544=>"111010000",
63545=>"100000100",
63546=>"111111111",
63547=>"010111110",
63548=>"100000001",
63549=>"111111111",
63550=>"000000001",
63551=>"001111110",
63552=>"111000101",
63553=>"000110111",
63554=>"111111000",
63555=>"110111011",
63556=>"100111111",
63557=>"001100110",
63558=>"011000011",
63559=>"111101011",
63560=>"110001000",
63561=>"000000000",
63562=>"100000101",
63563=>"000000100",
63564=>"011111110",
63565=>"101110011",
63566=>"100111111",
63567=>"010000010",
63568=>"010000000",
63569=>"111111111",
63570=>"000000011",
63571=>"001001001",
63572=>"111000001",
63573=>"111111111",
63574=>"011011011",
63575=>"011000100",
63576=>"111111101",
63577=>"101111111",
63578=>"000001001",
63579=>"110110010",
63580=>"111111100",
63581=>"000011000",
63582=>"000000000",
63583=>"001101111",
63584=>"000011010",
63585=>"110100010",
63586=>"100100100",
63587=>"000110111",
63588=>"100110000",
63589=>"110110111",
63590=>"011110000",
63591=>"111111000",
63592=>"111111111",
63593=>"111111000",
63594=>"110010111",
63595=>"101111000",
63596=>"000000111",
63597=>"011111000",
63598=>"100000000",
63599=>"011001111",
63600=>"100110111",
63601=>"000010111",
63602=>"101000100",
63603=>"000000001",
63604=>"000111000",
63605=>"000000000",
63606=>"001110110",
63607=>"110000000",
63608=>"100101111",
63609=>"111100000",
63610=>"000001000",
63611=>"000111011",
63612=>"011011001",
63613=>"010110100",
63614=>"110111010",
63615=>"000100000",
63616=>"000111011",
63617=>"111101100",
63618=>"010010110",
63619=>"011010011",
63620=>"000111000",
63621=>"000000000",
63622=>"001101111",
63623=>"011000100",
63624=>"001001011",
63625=>"000000111",
63626=>"111000000",
63627=>"101000110",
63628=>"000111000",
63629=>"110011000",
63630=>"100000000",
63631=>"001000001",
63632=>"001001100",
63633=>"011011111",
63634=>"111111011",
63635=>"011000001",
63636=>"011000000",
63637=>"101111110",
63638=>"001000000",
63639=>"000001011",
63640=>"011101110",
63641=>"101000101",
63642=>"111111110",
63643=>"010100000",
63644=>"000011111",
63645=>"111111110",
63646=>"010100111",
63647=>"000000100",
63648=>"010001111",
63649=>"000000111",
63650=>"000000000",
63651=>"111001000",
63652=>"011110010",
63653=>"000000010",
63654=>"001000001",
63655=>"100011010",
63656=>"111111000",
63657=>"000011010",
63658=>"111110111",
63659=>"000111111",
63660=>"011001111",
63661=>"111111111",
63662=>"111011010",
63663=>"000001000",
63664=>"000000010",
63665=>"010000000",
63666=>"000100100",
63667=>"011111011",
63668=>"100110000",
63669=>"000100110",
63670=>"011001010",
63671=>"000000100",
63672=>"001001110",
63673=>"111001000",
63674=>"000000010",
63675=>"100111111",
63676=>"011010000",
63677=>"101101101",
63678=>"010111111",
63679=>"111010001",
63680=>"100000000",
63681=>"000000101",
63682=>"010010010",
63683=>"111010101",
63684=>"111000100",
63685=>"010011111",
63686=>"010010111",
63687=>"101110111",
63688=>"110001100",
63689=>"111110100",
63690=>"010101111",
63691=>"101000100",
63692=>"000011111",
63693=>"010110100",
63694=>"000000100",
63695=>"000111111",
63696=>"000111111",
63697=>"000110110",
63698=>"000000100",
63699=>"000111111",
63700=>"000000000",
63701=>"010000001",
63702=>"010011000",
63703=>"101011111",
63704=>"000000100",
63705=>"101001010",
63706=>"000010111",
63707=>"000000000",
63708=>"100111110",
63709=>"111111111",
63710=>"001000001",
63711=>"011110000",
63712=>"111111010",
63713=>"000000000",
63714=>"000000000",
63715=>"101111100",
63716=>"000000100",
63717=>"111110000",
63718=>"000100111",
63719=>"111101010",
63720=>"000111111",
63721=>"000000100",
63722=>"111011011",
63723=>"101111110",
63724=>"100000000",
63725=>"110000111",
63726=>"010111010",
63727=>"010011001",
63728=>"000100000",
63729=>"010111101",
63730=>"000000010",
63731=>"000111110",
63732=>"101001111",
63733=>"010101010",
63734=>"001000000",
63735=>"001111010",
63736=>"000000100",
63737=>"010111111",
63738=>"000000000",
63739=>"001010010",
63740=>"101000000",
63741=>"111000010",
63742=>"110110110",
63743=>"111100001",
63744=>"011010010",
63745=>"010010010",
63746=>"000011110",
63747=>"111110010",
63748=>"001011001",
63749=>"010000010",
63750=>"111111111",
63751=>"111111100",
63752=>"000000000",
63753=>"001001101",
63754=>"110110010",
63755=>"101001101",
63756=>"101000000",
63757=>"111111000",
63758=>"111111011",
63759=>"001001101",
63760=>"000101110",
63761=>"010111000",
63762=>"001001001",
63763=>"000111111",
63764=>"010010010",
63765=>"001101100",
63766=>"000001000",
63767=>"010110111",
63768=>"000000000",
63769=>"111111111",
63770=>"100100111",
63771=>"111000000",
63772=>"000001111",
63773=>"101000111",
63774=>"010010111",
63775=>"001001001",
63776=>"000011011",
63777=>"000000001",
63778=>"001000000",
63779=>"000000000",
63780=>"011001011",
63781=>"110111100",
63782=>"000000000",
63783=>"000000000",
63784=>"000001101",
63785=>"000001000",
63786=>"110110010",
63787=>"111111101",
63788=>"011111111",
63789=>"101110110",
63790=>"111110100",
63791=>"000100000",
63792=>"010011110",
63793=>"101101101",
63794=>"000000001",
63795=>"110110111",
63796=>"111111111",
63797=>"111111110",
63798=>"001111010",
63799=>"110111010",
63800=>"010000010",
63801=>"111110010",
63802=>"000000001",
63803=>"000000100",
63804=>"000000000",
63805=>"111111111",
63806=>"111101010",
63807=>"100110010",
63808=>"010000100",
63809=>"111100110",
63810=>"101000000",
63811=>"011001101",
63812=>"000000000",
63813=>"010000101",
63814=>"110110110",
63815=>"001001011",
63816=>"101011000",
63817=>"001001111",
63818=>"111111000",
63819=>"010111111",
63820=>"001001010",
63821=>"111111111",
63822=>"100111111",
63823=>"110100000",
63824=>"111000100",
63825=>"110111010",
63826=>"000010010",
63827=>"001001011",
63828=>"001000000",
63829=>"100111001",
63830=>"100100100",
63831=>"000000111",
63832=>"000000111",
63833=>"110100000",
63834=>"111100100",
63835=>"110110110",
63836=>"000001111",
63837=>"001011011",
63838=>"110111111",
63839=>"100000111",
63840=>"111001101",
63841=>"000000000",
63842=>"001000001",
63843=>"001011111",
63844=>"100110100",
63845=>"000001001",
63846=>"100110111",
63847=>"111101101",
63848=>"000010001",
63849=>"000011111",
63850=>"111000100",
63851=>"001101010",
63852=>"000000101",
63853=>"110111010",
63854=>"010010000",
63855=>"100011111",
63856=>"001011001",
63857=>"110110000",
63858=>"110110011",
63859=>"001110110",
63860=>"111001000",
63861=>"000001000",
63862=>"000001000",
63863=>"100000100",
63864=>"010000000",
63865=>"110000000",
63866=>"011001010",
63867=>"001010111",
63868=>"100110110",
63869=>"100000100",
63870=>"111111100",
63871=>"000001111",
63872=>"000000000",
63873=>"111001111",
63874=>"010010000",
63875=>"001000101",
63876=>"000101111",
63877=>"101000000",
63878=>"110101011",
63879=>"111111010",
63880=>"101111111",
63881=>"100110000",
63882=>"100100000",
63883=>"000011101",
63884=>"011101101",
63885=>"000000101",
63886=>"111111110",
63887=>"100001000",
63888=>"101101100",
63889=>"111001001",
63890=>"110111111",
63891=>"011000000",
63892=>"000111101",
63893=>"000000000",
63894=>"001000000",
63895=>"100000000",
63896=>"000000000",
63897=>"111101100",
63898=>"101000001",
63899=>"000000100",
63900=>"000011110",
63901=>"111111001",
63902=>"111111000",
63903=>"111001001",
63904=>"111001000",
63905=>"000000001",
63906=>"110011110",
63907=>"101111110",
63908=>"000000111",
63909=>"110010110",
63910=>"000010111",
63911=>"000110011",
63912=>"010110110",
63913=>"000000000",
63914=>"111000000",
63915=>"000110000",
63916=>"011011111",
63917=>"001000101",
63918=>"100011000",
63919=>"110111101",
63920=>"011111101",
63921=>"101110100",
63922=>"101000101",
63923=>"000000000",
63924=>"111111111",
63925=>"010010101",
63926=>"100000110",
63927=>"000010000",
63928=>"001000100",
63929=>"110111111",
63930=>"110100111",
63931=>"010110001",
63932=>"000010100",
63933=>"000000000",
63934=>"000000001",
63935=>"111000110",
63936=>"010110010",
63937=>"111111010",
63938=>"010000000",
63939=>"111011011",
63940=>"111000000",
63941=>"100100100",
63942=>"010000010",
63943=>"110111111",
63944=>"111001100",
63945=>"111100110",
63946=>"111110000",
63947=>"111111111",
63948=>"010000000",
63949=>"011001110",
63950=>"111000010",
63951=>"111101000",
63952=>"000000000",
63953=>"111011111",
63954=>"111001011",
63955=>"001001000",
63956=>"101111111",
63957=>"110110000",
63958=>"100110010",
63959=>"111000000",
63960=>"110010010",
63961=>"000010111",
63962=>"100000000",
63963=>"000111111",
63964=>"111000100",
63965=>"000001111",
63966=>"000100011",
63967=>"111011010",
63968=>"000101001",
63969=>"111111111",
63970=>"111111101",
63971=>"110111110",
63972=>"100100110",
63973=>"010110001",
63974=>"010000000",
63975=>"111010000",
63976=>"001000000",
63977=>"010000010",
63978=>"010111010",
63979=>"001010000",
63980=>"000000000",
63981=>"001001111",
63982=>"001011000",
63983=>"101011000",
63984=>"000000000",
63985=>"011011001",
63986=>"111000111",
63987=>"010000000",
63988=>"110110000",
63989=>"000111110",
63990=>"000000110",
63991=>"000001001",
63992=>"000000000",
63993=>"110111101",
63994=>"111101111",
63995=>"110111111",
63996=>"000000111",
63997=>"000100000",
63998=>"100100001",
63999=>"110111010",
64000=>"001001111",
64001=>"000111111",
64002=>"110000000",
64003=>"111111111",
64004=>"000010011",
64005=>"000000001",
64006=>"111000000",
64007=>"000011001",
64008=>"000000000",
64009=>"111100001",
64010=>"110000000",
64011=>"111001010",
64012=>"000000101",
64013=>"001101111",
64014=>"010011011",
64015=>"111111111",
64016=>"000000000",
64017=>"001010010",
64018=>"010000000",
64019=>"000010011",
64020=>"101011111",
64021=>"111111011",
64022=>"011111111",
64023=>"111011111",
64024=>"111000000",
64025=>"101111011",
64026=>"000010110",
64027=>"011110111",
64028=>"010000101",
64029=>"110100000",
64030=>"111110111",
64031=>"111111111",
64032=>"100101000",
64033=>"111000011",
64034=>"100111011",
64035=>"111111101",
64036=>"011001011",
64037=>"111110111",
64038=>"100000010",
64039=>"001000000",
64040=>"111000000",
64041=>"111111011",
64042=>"000000000",
64043=>"000101101",
64044=>"001111111",
64045=>"111000000",
64046=>"111111101",
64047=>"111111000",
64048=>"111011000",
64049=>"001001001",
64050=>"100101111",
64051=>"101110000",
64052=>"111011000",
64053=>"110111111",
64054=>"000111111",
64055=>"000110111",
64056=>"111010110",
64057=>"000000111",
64058=>"001100000",
64059=>"101101111",
64060=>"011111011",
64061=>"111010111",
64062=>"000000111",
64063=>"000000000",
64064=>"111101000",
64065=>"111010011",
64066=>"111111101",
64067=>"001010000",
64068=>"111101111",
64069=>"000100000",
64070=>"000000000",
64071=>"111010010",
64072=>"100100111",
64073=>"000000000",
64074=>"000100101",
64075=>"101001111",
64076=>"100000000",
64077=>"000000000",
64078=>"000100110",
64079=>"000011000",
64080=>"000101011",
64081=>"111010000",
64082=>"011000000",
64083=>"111011001",
64084=>"000100111",
64085=>"111111100",
64086=>"011001001",
64087=>"101001000",
64088=>"101110000",
64089=>"001111111",
64090=>"000001001",
64091=>"101111111",
64092=>"110111111",
64093=>"110001001",
64094=>"101000000",
64095=>"000001100",
64096=>"000000111",
64097=>"000000000",
64098=>"100101111",
64099=>"000110110",
64100=>"001111111",
64101=>"100110100",
64102=>"000000000",
64103=>"111111110",
64104=>"000000000",
64105=>"111000000",
64106=>"011000000",
64107=>"111011111",
64108=>"000010000",
64109=>"111100000",
64110=>"011000111",
64111=>"000001000",
64112=>"000001110",
64113=>"111010101",
64114=>"000111011",
64115=>"111011000",
64116=>"111111111",
64117=>"101101101",
64118=>"111111111",
64119=>"101111111",
64120=>"000010000",
64121=>"111111111",
64122=>"000000001",
64123=>"011000000",
64124=>"000111110",
64125=>"111100100",
64126=>"100000000",
64127=>"111101100",
64128=>"111111111",
64129=>"111011000",
64130=>"011011011",
64131=>"010111001",
64132=>"000000000",
64133=>"001111111",
64134=>"111011010",
64135=>"000100111",
64136=>"000111011",
64137=>"000000000",
64138=>"000000000",
64139=>"111100000",
64140=>"000000000",
64141=>"011010010",
64142=>"111011111",
64143=>"000000000",
64144=>"011011111",
64145=>"000010111",
64146=>"101001111",
64147=>"110111000",
64148=>"000100101",
64149=>"111000000",
64150=>"001011011",
64151=>"000111111",
64152=>"001001000",
64153=>"111011000",
64154=>"111010000",
64155=>"000000111",
64156=>"100100100",
64157=>"000011011",
64158=>"111111110",
64159=>"111111111",
64160=>"000000010",
64161=>"101000000",
64162=>"111111111",
64163=>"111010001",
64164=>"111010000",
64165=>"000111111",
64166=>"111111111",
64167=>"000111111",
64168=>"111011000",
64169=>"011010111",
64170=>"000000000",
64171=>"101000000",
64172=>"111011001",
64173=>"110000000",
64174=>"001010110",
64175=>"000111011",
64176=>"000000010",
64177=>"000001111",
64178=>"111101100",
64179=>"000000000",
64180=>"000110110",
64181=>"101111011",
64182=>"000101111",
64183=>"101111000",
64184=>"110111111",
64185=>"000101101",
64186=>"101001010",
64187=>"010010111",
64188=>"001000010",
64189=>"111100000",
64190=>"010000110",
64191=>"101111111",
64192=>"111000100",
64193=>"000111111",
64194=>"011010111",
64195=>"110111111",
64196=>"101001000",
64197=>"001000000",
64198=>"010100000",
64199=>"101001101",
64200=>"010000000",
64201=>"000111111",
64202=>"110001111",
64203=>"000000111",
64204=>"000000000",
64205=>"110111111",
64206=>"000111111",
64207=>"111000100",
64208=>"111000000",
64209=>"000110111",
64210=>"001101001",
64211=>"111000110",
64212=>"111101110",
64213=>"001000110",
64214=>"111000111",
64215=>"101110000",
64216=>"111111111",
64217=>"000000111",
64218=>"100100100",
64219=>"111000000",
64220=>"111110101",
64221=>"111000000",
64222=>"101111111",
64223=>"100000010",
64224=>"101000101",
64225=>"111000100",
64226=>"111000000",
64227=>"000011111",
64228=>"000000010",
64229=>"010111111",
64230=>"000111111",
64231=>"000000000",
64232=>"000000000",
64233=>"000000000",
64234=>"001000000",
64235=>"000011011",
64236=>"000100101",
64237=>"001111101",
64238=>"111000000",
64239=>"111111111",
64240=>"111111101",
64241=>"011000000",
64242=>"111111111",
64243=>"000111111",
64244=>"011110111",
64245=>"000000000",
64246=>"111101011",
64247=>"101000100",
64248=>"101101111",
64249=>"101000000",
64250=>"111111000",
64251=>"000101111",
64252=>"101000101",
64253=>"000000000",
64254=>"101100110",
64255=>"000111011",
64256=>"100100110",
64257=>"010110000",
64258=>"100000001",
64259=>"010010000",
64260=>"011001000",
64261=>"000001110",
64262=>"100000000",
64263=>"111010100",
64264=>"011101001",
64265=>"100000000",
64266=>"111111010",
64267=>"111101001",
64268=>"000010010",
64269=>"011000101",
64270=>"100100100",
64271=>"000000000",
64272=>"100000000",
64273=>"111000001",
64274=>"010111111",
64275=>"100000000",
64276=>"110111111",
64277=>"010111111",
64278=>"001111010",
64279=>"110100000",
64280=>"001000000",
64281=>"111011000",
64282=>"000000110",
64283=>"111000100",
64284=>"100000000",
64285=>"000101101",
64286=>"000001111",
64287=>"100000100",
64288=>"011011000",
64289=>"111111110",
64290=>"100000000",
64291=>"011010000",
64292=>"011001011",
64293=>"000001011",
64294=>"111111111",
64295=>"010000111",
64296=>"010011000",
64297=>"000000000",
64298=>"000100110",
64299=>"000000000",
64300=>"111011011",
64301=>"001010100",
64302=>"000111111",
64303=>"011011011",
64304=>"011111111",
64305=>"111111111",
64306=>"001111010",
64307=>"000010000",
64308=>"000010111",
64309=>"111111111",
64310=>"100101011",
64311=>"100000000",
64312=>"101000111",
64313=>"000000001",
64314=>"010011010",
64315=>"100000000",
64316=>"010111001",
64317=>"111111111",
64318=>"000000000",
64319=>"111001100",
64320=>"000010010",
64321=>"000000110",
64322=>"010011011",
64323=>"110001101",
64324=>"011011011",
64325=>"101111111",
64326=>"100000001",
64327=>"110000111",
64328=>"111111010",
64329=>"111101000",
64330=>"000100110",
64331=>"101001000",
64332=>"101000000",
64333=>"101110110",
64334=>"110011011",
64335=>"011100000",
64336=>"000001000",
64337=>"111000000",
64338=>"100100111",
64339=>"001101011",
64340=>"101111100",
64341=>"001000001",
64342=>"000010000",
64343=>"010000000",
64344=>"111111011",
64345=>"011000100",
64346=>"000110100",
64347=>"011100110",
64348=>"101000000",
64349=>"110110110",
64350=>"010111110",
64351=>"011101101",
64352=>"001001101",
64353=>"000001101",
64354=>"000111111",
64355=>"011011011",
64356=>"011111111",
64357=>"010110111",
64358=>"010000110",
64359=>"111101101",
64360=>"101110000",
64361=>"111101111",
64362=>"000011100",
64363=>"000000011",
64364=>"011000000",
64365=>"011111111",
64366=>"000101101",
64367=>"000010011",
64368=>"110110110",
64369=>"110010001",
64370=>"001101111",
64371=>"000100001",
64372=>"000000000",
64373=>"100111111",
64374=>"000000000",
64375=>"000111111",
64376=>"000010111",
64377=>"111010110",
64378=>"001000101",
64379=>"010100111",
64380=>"011001001",
64381=>"000011111",
64382=>"000101000",
64383=>"111100100",
64384=>"000000010",
64385=>"101100111",
64386=>"111001110",
64387=>"111000000",
64388=>"101000000",
64389=>"111000001",
64390=>"000000100",
64391=>"000010000",
64392=>"111001011",
64393=>"001001111",
64394=>"110000101",
64395=>"000100010",
64396=>"110101000",
64397=>"000100001",
64398=>"110000001",
64399=>"000000000",
64400=>"011111111",
64401=>"001000000",
64402=>"000101100",
64403=>"011111110",
64404=>"100000000",
64405=>"011000000",
64406=>"111111111",
64407=>"011000100",
64408=>"000100001",
64409=>"000010001",
64410=>"111110100",
64411=>"000000000",
64412=>"110100101",
64413=>"011001000",
64414=>"001100111",
64415=>"101001000",
64416=>"111111111",
64417=>"010010100",
64418=>"011011000",
64419=>"101000000",
64420=>"011111011",
64421=>"101100100",
64422=>"110000000",
64423=>"010010010",
64424=>"111111010",
64425=>"000000000",
64426=>"111000000",
64427=>"000110111",
64428=>"010101101",
64429=>"000000101",
64430=>"111011111",
64431=>"011000000",
64432=>"001011001",
64433=>"011110110",
64434=>"010111011",
64435=>"010011001",
64436=>"011000000",
64437=>"001111111",
64438=>"011011010",
64439=>"000000000",
64440=>"011111100",
64441=>"111001001",
64442=>"000000000",
64443=>"100110110",
64444=>"000010100",
64445=>"111111111",
64446=>"010100100",
64447=>"000000000",
64448=>"000010111",
64449=>"101000100",
64450=>"000100100",
64451=>"100110110",
64452=>"010000101",
64453=>"001001000",
64454=>"000000000",
64455=>"000000111",
64456=>"110111111",
64457=>"000000000",
64458=>"100000000",
64459=>"111000111",
64460=>"100100100",
64461=>"110100101",
64462=>"011101100",
64463=>"001111111",
64464=>"111000000",
64465=>"010100110",
64466=>"111111100",
64467=>"010100000",
64468=>"000000001",
64469=>"001011011",
64470=>"011001011",
64471=>"000111111",
64472=>"110100100",
64473=>"101101000",
64474=>"111111011",
64475=>"011111111",
64476=>"110010110",
64477=>"011100000",
64478=>"111000000",
64479=>"000000000",
64480=>"000000000",
64481=>"000010111",
64482=>"110100101",
64483=>"000111011",
64484=>"000000000",
64485=>"000000100",
64486=>"101101000",
64487=>"010110111",
64488=>"000111010",
64489=>"001111000",
64490=>"111010110",
64491=>"000000000",
64492=>"001000000",
64493=>"010000000",
64494=>"101000011",
64495=>"111000100",
64496=>"100111111",
64497=>"001100100",
64498=>"111001110",
64499=>"111011010",
64500=>"001001001",
64501=>"110100000",
64502=>"000000010",
64503=>"111101101",
64504=>"111111110",
64505=>"000100101",
64506=>"100000010",
64507=>"000000100",
64508=>"000010111",
64509=>"111101101",
64510=>"100100010",
64511=>"000001101",
64512=>"101110100",
64513=>"100110000",
64514=>"011001001",
64515=>"100110000",
64516=>"011111000",
64517=>"000100100",
64518=>"001001111",
64519=>"111111011",
64520=>"001011011",
64521=>"011011010",
64522=>"111000001",
64523=>"000000000",
64524=>"000000111",
64525=>"100100000",
64526=>"100001011",
64527=>"011101111",
64528=>"110101000",
64529=>"100000100",
64530=>"111110101",
64531=>"110111001",
64532=>"000100111",
64533=>"000110100",
64534=>"101000101",
64535=>"101000000",
64536=>"100100000",
64537=>"000100100",
64538=>"100110000",
64539=>"111001111",
64540=>"101100110",
64541=>"010011011",
64542=>"000110100",
64543=>"001001011",
64544=>"001011000",
64545=>"100100100",
64546=>"001110110",
64547=>"111011011",
64548=>"001011011",
64549=>"000100000",
64550=>"011001001",
64551=>"110111110",
64552=>"000011000",
64553=>"100100000",
64554=>"000000011",
64555=>"011010000",
64556=>"111111101",
64557=>"110000100",
64558=>"000100110",
64559=>"000100000",
64560=>"000100100",
64561=>"001001001",
64562=>"100110100",
64563=>"100101100",
64564=>"100110011",
64565=>"101000000",
64566=>"001011110",
64567=>"111111011",
64568=>"100100100",
64569=>"100100110",
64570=>"110110100",
64571=>"110110110",
64572=>"000001001",
64573=>"011011011",
64574=>"000100100",
64575=>"011011111",
64576=>"111111111",
64577=>"110100011",
64578=>"101111111",
64579=>"011011110",
64580=>"100110111",
64581=>"100110100",
64582=>"001001110",
64583=>"000011111",
64584=>"100010000",
64585=>"011011000",
64586=>"100100000",
64587=>"101100100",
64588=>"010001001",
64589=>"011000101",
64590=>"000111111",
64591=>"011100000",
64592=>"011011010",
64593=>"011011100",
64594=>"111111110",
64595=>"000100010",
64596=>"011100100",
64597=>"100110001",
64598=>"111111101",
64599=>"111100110",
64600=>"110110110",
64601=>"110110000",
64602=>"001000001",
64603=>"100110110",
64604=>"100100100",
64605=>"000100001",
64606=>"100100100",
64607=>"101011111",
64608=>"011001011",
64609=>"111110000",
64610=>"011001111",
64611=>"110101111",
64612=>"010111111",
64613=>"001011000",
64614=>"111001111",
64615=>"011011011",
64616=>"000110011",
64617=>"110110000",
64618=>"001000110",
64619=>"000110111",
64620=>"100110001",
64621=>"110001010",
64622=>"000001111",
64623=>"000100101",
64624=>"110111001",
64625=>"100110100",
64626=>"011001001",
64627=>"100110011",
64628=>"111110111",
64629=>"100100100",
64630=>"110100000",
64631=>"011001001",
64632=>"001010001",
64633=>"111000000",
64634=>"000100100",
64635=>"100110011",
64636=>"010011001",
64637=>"010110100",
64638=>"011011011",
64639=>"011001011",
64640=>"000101111",
64641=>"010010001",
64642=>"111000110",
64643=>"111110011",
64644=>"010100100",
64645=>"111000111",
64646=>"011110100",
64647=>"111111110",
64648=>"000001011",
64649=>"111011111",
64650=>"111101100",
64651=>"000110111",
64652=>"011001001",
64653=>"101001110",
64654=>"001111001",
64655=>"000100100",
64656=>"000011001",
64657=>"001010011",
64658=>"000011011",
64659=>"011110110",
64660=>"000000010",
64661=>"100100110",
64662=>"101100001",
64663=>"000100100",
64664=>"000001000",
64665=>"001100100",
64666=>"111011000",
64667=>"100001001",
64668=>"100111110",
64669=>"011011011",
64670=>"100100110",
64671=>"000000000",
64672=>"100111011",
64673=>"110100100",
64674=>"011000010",
64675=>"100101001",
64676=>"110000110",
64677=>"001001011",
64678=>"101100100",
64679=>"010001011",
64680=>"100100100",
64681=>"110010000",
64682=>"110111100",
64683=>"110110011",
64684=>"111111011",
64685=>"001000000",
64686=>"011110001",
64687=>"000001011",
64688=>"100000010",
64689=>"001001000",
64690=>"100100110",
64691=>"111110011",
64692=>"011011011",
64693=>"000000011",
64694=>"100110110",
64695=>"000100000",
64696=>"000100110",
64697=>"000000000",
64698=>"001011000",
64699=>"001011111",
64700=>"000100000",
64701=>"011011011",
64702=>"011001001",
64703=>"000000100",
64704=>"001011111",
64705=>"111011011",
64706=>"110111001",
64707=>"001001001",
64708=>"100100000",
64709=>"000100100",
64710=>"000000100",
64711=>"010011000",
64712=>"011001011",
64713=>"010000000",
64714=>"100110001",
64715=>"101011111",
64716=>"001001010",
64717=>"001011011",
64718=>"011011000",
64719=>"001001111",
64720=>"100011111",
64721=>"011101011",
64722=>"001100000",
64723=>"001001110",
64724=>"011011011",
64725=>"111111000",
64726=>"100010000",
64727=>"000110100",
64728=>"001011111",
64729=>"100000000",
64730=>"010100101",
64731=>"100100100",
64732=>"111110100",
64733=>"110110101",
64734=>"110100110",
64735=>"000100100",
64736=>"001000001",
64737=>"000101100",
64738=>"011011111",
64739=>"111011010",
64740=>"101001001",
64741=>"110010100",
64742=>"011011011",
64743=>"011011111",
64744=>"010110100",
64745=>"001000010",
64746=>"000000000",
64747=>"111001000",
64748=>"100000000",
64749=>"111111110",
64750=>"000000000",
64751=>"100000000",
64752=>"001110110",
64753=>"101111100",
64754=>"100100100",
64755=>"111111101",
64756=>"000111110",
64757=>"110111111",
64758=>"100101101",
64759=>"101000000",
64760=>"100100110",
64761=>"110010110",
64762=>"100100100",
64763=>"011111001",
64764=>"111010011",
64765=>"110001101",
64766=>"100010111",
64767=>"111010010",
64768=>"100000000",
64769=>"111110101",
64770=>"110000100",
64771=>"011011011",
64772=>"100000000",
64773=>"111000000",
64774=>"110110110",
64775=>"011110011",
64776=>"000110111",
64777=>"011110100",
64778=>"100100000",
64779=>"100010011",
64780=>"001011111",
64781=>"000011111",
64782=>"000001001",
64783=>"110011011",
64784=>"100100110",
64785=>"000100110",
64786=>"000001011",
64787=>"100110011",
64788=>"100110011",
64789=>"011001000",
64790=>"111010000",
64791=>"100100100",
64792=>"110110110",
64793=>"111111111",
64794=>"000001101",
64795=>"000011001",
64796=>"010011011",
64797=>"000100100",
64798=>"000100110",
64799=>"000000100",
64800=>"111100100",
64801=>"000011001",
64802=>"101100100",
64803=>"110000100",
64804=>"100110000",
64805=>"000111111",
64806=>"100100100",
64807=>"000111000",
64808=>"111010110",
64809=>"000000100",
64810=>"001100100",
64811=>"011000011",
64812=>"001100011",
64813=>"000110111",
64814=>"001000100",
64815=>"011111011",
64816=>"100100011",
64817=>"000001000",
64818=>"000000001",
64819=>"100111111",
64820=>"100000000",
64821=>"100111011",
64822=>"100100110",
64823=>"010111100",
64824=>"011000000",
64825=>"000000100",
64826=>"000000010",
64827=>"100111111",
64828=>"001100110",
64829=>"111111110",
64830=>"000101101",
64831=>"110111110",
64832=>"110110110",
64833=>"100110010",
64834=>"011001000",
64835=>"001001100",
64836=>"110100110",
64837=>"100000100",
64838=>"111110110",
64839=>"011001000",
64840=>"001110110",
64841=>"101011111",
64842=>"100100110",
64843=>"000100101",
64844=>"111110100",
64845=>"000100110",
64846=>"100111110",
64847=>"111100001",
64848=>"000000000",
64849=>"111111001",
64850=>"111110111",
64851=>"000010010",
64852=>"000011011",
64853=>"001000000",
64854=>"001100110",
64855=>"000011011",
64856=>"001011101",
64857=>"010010100",
64858=>"101001100",
64859=>"001001100",
64860=>"010111011",
64861=>"001000101",
64862=>"111111110",
64863=>"110100000",
64864=>"110110110",
64865=>"000000100",
64866=>"110110100",
64867=>"011001011",
64868=>"100000010",
64869=>"000010100",
64870=>"000001011",
64871=>"111001011",
64872=>"101110110",
64873=>"010100100",
64874=>"011011011",
64875=>"111100110",
64876=>"111000111",
64877=>"000000011",
64878=>"011011000",
64879=>"010000111",
64880=>"100110110",
64881=>"001111011",
64882=>"100100100",
64883=>"101000100",
64884=>"011011011",
64885=>"100100100",
64886=>"011011010",
64887=>"000111011",
64888=>"011000011",
64889=>"000100110",
64890=>"100100100",
64891=>"001011111",
64892=>"100110110",
64893=>"100000000",
64894=>"011011100",
64895=>"000011000",
64896=>"110110010",
64897=>"111100000",
64898=>"000111110",
64899=>"000101000",
64900=>"000100011",
64901=>"001101111",
64902=>"110010001",
64903=>"100000001",
64904=>"100100101",
64905=>"100110111",
64906=>"110110100",
64907=>"011111110",
64908=>"101011100",
64909=>"000111111",
64910=>"001111111",
64911=>"100100100",
64912=>"100111110",
64913=>"111111000",
64914=>"000010000",
64915=>"000100110",
64916=>"000000100",
64917=>"000000000",
64918=>"101100111",
64919=>"110000000",
64920=>"111111011",
64921=>"000000011",
64922=>"111000000",
64923=>"001000011",
64924=>"110011001",
64925=>"000100100",
64926=>"000001111",
64927=>"110100111",
64928=>"111110110",
64929=>"100111110",
64930=>"101000000",
64931=>"100110111",
64932=>"000000111",
64933=>"100111110",
64934=>"100100101",
64935=>"111111111",
64936=>"000100000",
64937=>"001011011",
64938=>"111011011",
64939=>"111000000",
64940=>"000011101",
64941=>"000011000",
64942=>"001100111",
64943=>"011001011",
64944=>"111011000",
64945=>"010011010",
64946=>"111101000",
64947=>"001000000",
64948=>"010011011",
64949=>"101101000",
64950=>"000011011",
64951=>"100010111",
64952=>"110000001",
64953=>"000110100",
64954=>"011001000",
64955=>"100000011",
64956=>"111101000",
64957=>"011011011",
64958=>"000001001",
64959=>"111011000",
64960=>"010100100",
64961=>"000001000",
64962=>"001011011",
64963=>"101001000",
64964=>"000000110",
64965=>"100100111",
64966=>"111110000",
64967=>"001000100",
64968=>"000100010",
64969=>"010111111",
64970=>"110010010",
64971=>"100100111",
64972=>"110011000",
64973=>"000000110",
64974=>"110000100",
64975=>"100011011",
64976=>"011011000",
64977=>"000000000",
64978=>"100010011",
64979=>"101111000",
64980=>"111111111",
64981=>"100000101",
64982=>"111100111",
64983=>"111100000",
64984=>"011111111",
64985=>"000000111",
64986=>"101111111",
64987=>"111100111",
64988=>"100110110",
64989=>"000001011",
64990=>"001011111",
64991=>"000000001",
64992=>"010010000",
64993=>"101011011",
64994=>"001011011",
64995=>"100110110",
64996=>"100110000",
64997=>"001000010",
64998=>"011101101",
64999=>"110110001",
65000=>"011011101",
65001=>"100111001",
65002=>"000100110",
65003=>"101000100",
65004=>"011011011",
65005=>"111111110",
65006=>"110000000",
65007=>"000100000",
65008=>"000100100",
65009=>"100000111",
65010=>"011000000",
65011=>"011011010",
65012=>"000110100",
65013=>"111101111",
65014=>"011011111",
65015=>"001001001",
65016=>"100100000",
65017=>"011001001",
65018=>"111100100",
65019=>"000000111",
65020=>"111000000",
65021=>"001011100",
65022=>"100110101",
65023=>"000000111",
65024=>"011001101",
65025=>"110101100",
65026=>"000000110",
65027=>"000000110",
65028=>"001010110",
65029=>"000010010",
65030=>"110110000",
65031=>"011111111",
65032=>"001000111",
65033=>"001000000",
65034=>"000111111",
65035=>"000011110",
65036=>"001001101",
65037=>"000000000",
65038=>"010001011",
65039=>"111100011",
65040=>"111110010",
65041=>"111000000",
65042=>"110101100",
65043=>"011110000",
65044=>"101101101",
65045=>"111111101",
65046=>"110010010",
65047=>"010111000",
65048=>"000111000",
65049=>"111000000",
65050=>"011011000",
65051=>"000010010",
65052=>"101001000",
65053=>"000000000",
65054=>"110111011",
65055=>"000000101",
65056=>"000000111",
65057=>"000000000",
65058=>"000101100",
65059=>"000011010",
65060=>"011000100",
65061=>"110001011",
65062=>"010111111",
65063=>"101001000",
65064=>"111010111",
65065=>"000011000",
65066=>"100111111",
65067=>"111011000",
65068=>"111100001",
65069=>"101101000",
65070=>"111000101",
65071=>"010001000",
65072=>"111000000",
65073=>"001011011",
65074=>"010000000",
65075=>"001000000",
65076=>"110011111",
65077=>"011101101",
65078=>"111110101",
65079=>"111101000",
65080=>"111000000",
65081=>"000000000",
65082=>"000000100",
65083=>"010000001",
65084=>"100000000",
65085=>"010001000",
65086=>"000101100",
65087=>"011111111",
65088=>"110011000",
65089=>"111000101",
65090=>"101000101",
65091=>"001010011",
65092=>"000010000",
65093=>"001101111",
65094=>"001000000",
65095=>"111101000",
65096=>"111001100",
65097=>"000011111",
65098=>"000100101",
65099=>"111111101",
65100=>"111000001",
65101=>"000001011",
65102=>"000000111",
65103=>"111111111",
65104=>"000000000",
65105=>"110000000",
65106=>"111111001",
65107=>"011001110",
65108=>"110111001",
65109=>"111111000",
65110=>"011001001",
65111=>"101010011",
65112=>"000000000",
65113=>"000000101",
65114=>"000111111",
65115=>"110000100",
65116=>"111111000",
65117=>"000001111",
65118=>"011000111",
65119=>"000000110",
65120=>"111111111",
65121=>"000000110",
65122=>"001110111",
65123=>"011000101",
65124=>"000001110",
65125=>"000010001",
65126=>"011111111",
65127=>"001111010",
65128=>"001000110",
65129=>"101000000",
65130=>"101001011",
65131=>"111111000",
65132=>"111000000",
65133=>"000111111",
65134=>"111000000",
65135=>"111011001",
65136=>"101111111",
65137=>"110001100",
65138=>"011111011",
65139=>"101000001",
65140=>"111000001",
65141=>"111000000",
65142=>"000000001",
65143=>"000000101",
65144=>"000111111",
65145=>"111101100",
65146=>"000000000",
65147=>"000000010",
65148=>"000000010",
65149=>"100000110",
65150=>"000010111",
65151=>"000111111",
65152=>"010000000",
65153=>"000000000",
65154=>"111010000",
65155=>"100010010",
65156=>"101101101",
65157=>"110101111",
65158=>"111001101",
65159=>"100000100",
65160=>"000011111",
65161=>"100011111",
65162=>"000111111",
65163=>"100110110",
65164=>"000110111",
65165=>"111111101",
65166=>"010001000",
65167=>"000000001",
65168=>"111001101",
65169=>"000000111",
65170=>"000010000",
65171=>"000000001",
65172=>"010010010",
65173=>"111010010",
65174=>"100011111",
65175=>"000000001",
65176=>"111011000",
65177=>"111110100",
65178=>"000000010",
65179=>"000001111",
65180=>"110001010",
65181=>"000000111",
65182=>"101000000",
65183=>"111000000",
65184=>"000000111",
65185=>"000100000",
65186=>"000111111",
65187=>"100010101",
65188=>"111111000",
65189=>"110000011",
65190=>"011110110",
65191=>"000100111",
65192=>"111010000",
65193=>"000001000",
65194=>"110110111",
65195=>"000000000",
65196=>"111111111",
65197=>"011000010",
65198=>"100101110",
65199=>"001111100",
65200=>"101111110",
65201=>"001001001",
65202=>"000001111",
65203=>"000001100",
65204=>"011111110",
65205=>"000111101",
65206=>"111111100",
65207=>"000011111",
65208=>"001000010",
65209=>"000011010",
65210=>"100010000",
65211=>"101000011",
65212=>"000000101",
65213=>"000001111",
65214=>"000111111",
65215=>"111000000",
65216=>"111101101",
65217=>"110111000",
65218=>"101010000",
65219=>"001001101",
65220=>"111000000",
65221=>"110110100",
65222=>"111111100",
65223=>"000000000",
65224=>"011001111",
65225=>"111010010",
65226=>"111010000",
65227=>"011010010",
65228=>"000110111",
65229=>"000011100",
65230=>"000111100",
65231=>"000110000",
65232=>"000010111",
65233=>"011001110",
65234=>"010000000",
65235=>"001000010",
65236=>"000011001",
65237=>"100101111",
65238=>"100010010",
65239=>"011000000",
65240=>"111100000",
65241=>"011011000",
65242=>"000001111",
65243=>"010000101",
65244=>"111000000",
65245=>"101100111",
65246=>"010110000",
65247=>"000111100",
65248=>"101000010",
65249=>"111000111",
65250=>"000000010",
65251=>"111100110",
65252=>"001100000",
65253=>"010101101",
65254=>"011000111",
65255=>"111101101",
65256=>"100011000",
65257=>"111111101",
65258=>"001010111",
65259=>"111010000",
65260=>"000011111",
65261=>"110000100",
65262=>"000000000",
65263=>"100011100",
65264=>"111111010",
65265=>"111011111",
65266=>"111000010",
65267=>"111111001",
65268=>"110100101",
65269=>"000101111",
65270=>"000001001",
65271=>"110000001",
65272=>"111000000",
65273=>"000111111",
65274=>"111000100",
65275=>"001111101",
65276=>"000111110",
65277=>"111111000",
65278=>"110010111",
65279=>"100100000",
65280=>"000001001",
65281=>"001000111",
65282=>"000000000",
65283=>"000000110",
65284=>"111000101",
65285=>"000000111",
65286=>"000101110",
65287=>"000000010",
65288=>"101000000",
65289=>"000110111",
65290=>"000010110",
65291=>"111000010",
65292=>"000000000",
65293=>"110010001",
65294=>"000000000",
65295=>"110111111",
65296=>"000001001",
65297=>"111111111",
65298=>"010000101",
65299=>"000111110",
65300=>"001100110",
65301=>"001000000",
65302=>"011101100",
65303=>"010010111",
65304=>"000000000",
65305=>"111000111",
65306=>"100100001",
65307=>"000111100",
65308=>"000101110",
65309=>"101100100",
65310=>"101000000",
65311=>"101101101",
65312=>"100001100",
65313=>"110111011",
65314=>"000000010",
65315=>"000111111",
65316=>"000000011",
65317=>"000000111",
65318=>"011001000",
65319=>"000101111",
65320=>"111111010",
65321=>"110100111",
65322=>"000111111",
65323=>"001011110",
65324=>"111011111",
65325=>"000000000",
65326=>"000000000",
65327=>"010101110",
65328=>"001001000",
65329=>"000100000",
65330=>"000000011",
65331=>"000101100",
65332=>"010111111",
65333=>"111111111",
65334=>"110111011",
65335=>"100010011",
65336=>"101000111",
65337=>"000101101",
65338=>"000110000",
65339=>"101000000",
65340=>"100001000",
65341=>"111111000",
65342=>"101010110",
65343=>"010111001",
65344=>"111111111",
65345=>"010101011",
65346=>"011000111",
65347=>"000001111",
65348=>"010111010",
65349=>"001000111",
65350=>"000111111",
65351=>"110001010",
65352=>"000100111",
65353=>"110111111",
65354=>"000001000",
65355=>"000010001",
65356=>"000000010",
65357=>"000011111",
65358=>"111100110",
65359=>"010010111",
65360=>"111111111",
65361=>"111111000",
65362=>"000100110",
65363=>"001100110",
65364=>"110100000",
65365=>"100000110",
65366=>"000101111",
65367=>"000000000",
65368=>"000001101",
65369=>"111001011",
65370=>"000111111",
65371=>"011011110",
65372=>"111111111",
65373=>"000000000",
65374=>"010110101",
65375=>"000010111",
65376=>"110101111",
65377=>"000111110",
65378=>"000101111",
65379=>"010110100",
65380=>"000100100",
65381=>"111111100",
65382=>"010111110",
65383=>"000011111",
65384=>"000101011",
65385=>"000000000",
65386=>"000000110",
65387=>"010001110",
65388=>"010000100",
65389=>"000000010",
65390=>"000001001",
65391=>"111111001",
65392=>"100000010",
65393=>"111110111",
65394=>"011111110",
65395=>"000001011",
65396=>"000000011",
65397=>"000000000",
65398=>"000110011",
65399=>"111111111",
65400=>"011010111",
65401=>"110111101",
65402=>"000001000",
65403=>"111000111",
65404=>"001011010",
65405=>"110000010",
65406=>"111100001",
65407=>"000001000",
65408=>"110110100",
65409=>"111101000",
65410=>"111001000",
65411=>"111111010",
65412=>"001101000",
65413=>"111101100",
65414=>"110100110",
65415=>"001000000",
65416=>"001000100",
65417=>"000001101",
65418=>"010011010",
65419=>"101110111",
65420=>"101101011",
65421=>"111100101",
65422=>"111000000",
65423=>"000000000",
65424=>"001001011",
65425=>"010101111",
65426=>"000000010",
65427=>"000000000",
65428=>"101000100",
65429=>"000000010",
65430=>"100111001",
65431=>"010011011",
65432=>"010000111",
65433=>"001000011",
65434=>"011110111",
65435=>"101000000",
65436=>"000100101",
65437=>"111111010",
65438=>"000000111",
65439=>"100111011",
65440=>"011000000",
65441=>"110000000",
65442=>"111100010",
65443=>"000010000",
65444=>"111001010",
65445=>"110000000",
65446=>"001111000",
65447=>"010110110",
65448=>"000000000",
65449=>"110111000",
65450=>"111010000",
65451=>"000110110",
65452=>"100000101",
65453=>"000101010",
65454=>"000010011",
65455=>"111011110",
65456=>"011000000",
65457=>"000001100",
65458=>"010100000",
65459=>"001000100",
65460=>"111000001",
65461=>"111010100",
65462=>"111111101",
65463=>"001101111",
65464=>"001100000",
65465=>"100000001",
65466=>"001000000",
65467=>"000000010",
65468=>"000010000",
65469=>"000100111",
65470=>"001000000",
65471=>"010010111",
65472=>"000000000",
65473=>"000000000",
65474=>"010000111",
65475=>"000101001",
65476=>"000001000",
65477=>"100000011",
65478=>"000000001",
65479=>"010011000",
65480=>"101000101",
65481=>"110010000",
65482=>"111010010",
65483=>"110000000",
65484=>"000000000",
65485=>"100110110",
65486=>"011010010",
65487=>"111111011",
65488=>"100000010",
65489=>"110100111",
65490=>"111000011",
65491=>"110000010",
65492=>"101101111",
65493=>"000100100",
65494=>"010101111",
65495=>"001111001",
65496=>"000000111",
65497=>"111000000",
65498=>"111110000",
65499=>"000000111",
65500=>"110001001",
65501=>"111110010",
65502=>"111111000",
65503=>"111011001",
65504=>"000111111",
65505=>"001001000",
65506=>"000000110",
65507=>"000000010",
65508=>"010000000",
65509=>"111001000",
65510=>"111000110",
65511=>"111101100",
65512=>"111000111",
65513=>"111111110",
65514=>"000100010",
65515=>"000000111",
65516=>"001001000",
65517=>"111011111",
65518=>"000000000",
65519=>"001111001",
65520=>"111000000",
65521=>"001000010",
65522=>"010000010",
65523=>"111001101",
65524=>"100101111",
65525=>"000001000",
65526=>"000010010",
65527=>"001001101",
65528=>"000000111",
65529=>"000000101",
65530=>"111011110",
65531=>"101001000",
65532=>"000011001",
65533=>"111100110",
65534=>"000111111",
65535=>"000000000",
65536=>"111001011",
65537=>"001101011",
65538=>"000000100",
65539=>"000010111",
65540=>"100000001",
65541=>"111010000",
65542=>"000101011",
65543=>"010000111",
65544=>"000000111",
65545=>"111000000",
65546=>"010000000",
65547=>"000010101",
65548=>"111111111",
65549=>"011000101",
65550=>"100001001",
65551=>"101000000",
65552=>"000000100",
65553=>"111110000",
65554=>"000010000",
65555=>"111000111",
65556=>"111011111",
65557=>"000100010",
65558=>"000010000",
65559=>"011001011",
65560=>"111000000",
65561=>"001101000",
65562=>"000000000",
65563=>"000011000",
65564=>"011000100",
65565=>"100100111",
65566=>"111001100",
65567=>"000101111",
65568=>"000010000",
65569=>"011111111",
65570=>"000010110",
65571=>"010000000",
65572=>"110011111",
65573=>"110110111",
65574=>"000011111",
65575=>"000111111",
65576=>"111111111",
65577=>"111111111",
65578=>"000000000",
65579=>"000110110",
65580=>"011111111",
65581=>"111110011",
65582=>"111101000",
65583=>"000001111",
65584=>"000000000",
65585=>"110000000",
65586=>"000000100",
65587=>"101000000",
65588=>"100000000",
65589=>"111111101",
65590=>"000000000",
65591=>"000000001",
65592=>"111101001",
65593=>"001110110",
65594=>"000010110",
65595=>"111111001",
65596=>"100000111",
65597=>"010111011",
65598=>"000000000",
65599=>"011010110",
65600=>"000000000",
65601=>"111110000",
65602=>"111111111",
65603=>"011001011",
65604=>"100111111",
65605=>"111110010",
65606=>"000000000",
65607=>"010000001",
65608=>"111011110",
65609=>"010000100",
65610=>"010010000",
65611=>"100000000",
65612=>"000000011",
65613=>"110110100",
65614=>"011001100",
65615=>"111111110",
65616=>"000110111",
65617=>"010011000",
65618=>"011101111",
65619=>"011101011",
65620=>"000000010",
65621=>"100110111",
65622=>"001001101",
65623=>"000000000",
65624=>"111111010",
65625=>"111111111",
65626=>"100100111",
65627=>"001100111",
65628=>"000100100",
65629=>"011001001",
65630=>"011111000",
65631=>"100100100",
65632=>"000010111",
65633=>"000010111",
65634=>"111000111",
65635=>"000000010",
65636=>"111111000",
65637=>"000010011",
65638=>"000000111",
65639=>"101100000",
65640=>"011100000",
65641=>"010000110",
65642=>"000000000",
65643=>"111111100",
65644=>"010110101",
65645=>"100011000",
65646=>"000001010",
65647=>"111111001",
65648=>"100100111",
65649=>"000000111",
65650=>"000000000",
65651=>"011111011",
65652=>"111000000",
65653=>"101000000",
65654=>"000010111",
65655=>"011011111",
65656=>"000001111",
65657=>"111100010",
65658=>"001001111",
65659=>"110101100",
65660=>"000000000",
65661=>"110100100",
65662=>"000011110",
65663=>"000000100",
65664=>"111111110",
65665=>"111000100",
65666=>"000010111",
65667=>"101101010",
65668=>"000000010",
65669=>"101101011",
65670=>"011011011",
65671=>"001001100",
65672=>"100001101",
65673=>"001101101",
65674=>"000011000",
65675=>"011011000",
65676=>"000010101",
65677=>"110111100",
65678=>"110011000",
65679=>"000000000",
65680=>"100000100",
65681=>"001000101",
65682=>"101101111",
65683=>"101100000",
65684=>"000001001",
65685=>"000010001",
65686=>"010001000",
65687=>"011011111",
65688=>"010010000",
65689=>"000010011",
65690=>"101000110",
65691=>"000000000",
65692=>"000000000",
65693=>"110110000",
65694=>"001001001",
65695=>"000001000",
65696=>"011000100",
65697=>"101000000",
65698=>"111111111",
65699=>"011001100",
65700=>"010000000",
65701=>"100100110",
65702=>"010110001",
65703=>"010101000",
65704=>"000111000",
65705=>"000000111",
65706=>"010010001",
65707=>"111010000",
65708=>"100110001",
65709=>"111111111",
65710=>"100001000",
65711=>"011111111",
65712=>"011001010",
65713=>"101001011",
65714=>"110010000",
65715=>"010010000",
65716=>"001101110",
65717=>"111110100",
65718=>"000111111",
65719=>"010111000",
65720=>"011100111",
65721=>"100101001",
65722=>"111011000",
65723=>"111000000",
65724=>"111111111",
65725=>"000111011",
65726=>"011011011",
65727=>"000000011",
65728=>"000000000",
65729=>"010111000",
65730=>"000000111",
65731=>"100100111",
65732=>"000011010",
65733=>"011010001",
65734=>"000000100",
65735=>"010111011",
65736=>"000000111",
65737=>"000010010",
65738=>"111111110",
65739=>"001000001",
65740=>"100000101",
65741=>"000000010",
65742=>"001010111",
65743=>"010011000",
65744=>"000011111",
65745=>"110110111",
65746=>"100001010",
65747=>"111101111",
65748=>"000000001",
65749=>"000000100",
65750=>"111111001",
65751=>"000111010",
65752=>"001101111",
65753=>"001000011",
65754=>"111111111",
65755=>"000101010",
65756=>"000000101",
65757=>"010011011",
65758=>"100111111",
65759=>"111101101",
65760=>"100010111",
65761=>"000001001",
65762=>"111111111",
65763=>"100000000",
65764=>"111111111",
65765=>"000000101",
65766=>"010000110",
65767=>"001000000",
65768=>"000010111",
65769=>"100100000",
65770=>"110100000",
65771=>"000000010",
65772=>"011111111",
65773=>"000000110",
65774=>"010000000",
65775=>"000000001",
65776=>"000000111",
65777=>"000001000",
65778=>"111111101",
65779=>"111111111",
65780=>"110100010",
65781=>"000000000",
65782=>"101000000",
65783=>"000000000",
65784=>"000000000",
65785=>"111111010",
65786=>"000000000",
65787=>"000000111",
65788=>"111111100",
65789=>"000000100",
65790=>"000000100",
65791=>"010101000",
65792=>"000000000",
65793=>"110001011",
65794=>"001001001",
65795=>"100111111",
65796=>"101100101",
65797=>"101101111",
65798=>"110010010",
65799=>"100110100",
65800=>"101000111",
65801=>"011011011",
65802=>"111111111",
65803=>"011001011",
65804=>"011011001",
65805=>"000000001",
65806=>"010011100",
65807=>"001000000",
65808=>"001001001",
65809=>"110000111",
65810=>"101100100",
65811=>"000011010",
65812=>"000100100",
65813=>"011011011",
65814=>"011011011",
65815=>"000101101",
65816=>"000000100",
65817=>"100101110",
65818=>"001100000",
65819=>"011011011",
65820=>"010100011",
65821=>"011010000",
65822=>"011011001",
65823=>"001000100",
65824=>"010011000",
65825=>"100100101",
65826=>"010001000",
65827=>"000010011",
65828=>"100100101",
65829=>"100100000",
65830=>"111100100",
65831=>"110100111",
65832=>"100100110",
65833=>"100100110",
65834=>"101001101",
65835=>"011010001",
65836=>"111111100",
65837=>"011001101",
65838=>"010100110",
65839=>"111110110",
65840=>"111001011",
65841=>"101100100",
65842=>"001001011",
65843=>"011101111",
65844=>"111100000",
65845=>"101100101",
65846=>"111010001",
65847=>"000000000",
65848=>"110000100",
65849=>"111000110",
65850=>"000011111",
65851=>"011000111",
65852=>"000010100",
65853=>"100100100",
65854=>"010011011",
65855=>"100101101",
65856=>"111111111",
65857=>"110100100",
65858=>"101100010",
65859=>"011011011",
65860=>"100100000",
65861=>"011000000",
65862=>"001001000",
65863=>"110111110",
65864=>"000011001",
65865=>"101101101",
65866=>"110011000",
65867=>"100100101",
65868=>"111101111",
65869=>"100100100",
65870=>"100100100",
65871=>"101100011",
65872=>"100100100",
65873=>"100000111",
65874=>"100000101",
65875=>"011001000",
65876=>"100110111",
65877=>"111101111",
65878=>"110100101",
65879=>"011011011",
65880=>"100100100",
65881=>"100100000",
65882=>"100100100",
65883=>"000100000",
65884=>"011111111",
65885=>"000000011",
65886=>"011011011",
65887=>"111011000",
65888=>"011011011",
65889=>"101011011",
65890=>"010011111",
65891=>"100110000",
65892=>"000011000",
65893=>"101100001",
65894=>"111111000",
65895=>"000000010",
65896=>"010111111",
65897=>"000001100",
65898=>"110111111",
65899=>"100001011",
65900=>"100101111",
65901=>"000101101",
65902=>"011000001",
65903=>"010100011",
65904=>"111111111",
65905=>"011001010",
65906=>"011101011",
65907=>"110110011",
65908=>"000001111",
65909=>"000000010",
65910=>"111111001",
65911=>"111111010",
65912=>"011010011",
65913=>"100100100",
65914=>"111110110",
65915=>"001011000",
65916=>"100000111",
65917=>"000000110",
65918=>"000011001",
65919=>"111111101",
65920=>"101000000",
65921=>"000000011",
65922=>"011011011",
65923=>"000110110",
65924=>"101111101",
65925=>"111111001",
65926=>"100101110",
65927=>"100100100",
65928=>"100100000",
65929=>"011000100",
65930=>"001011011",
65931=>"011000110",
65932=>"011011001",
65933=>"111111000",
65934=>"111111010",
65935=>"000000111",
65936=>"110110100",
65937=>"101001011",
65938=>"000001111",
65939=>"101111100",
65940=>"100101101",
65941=>"011011011",
65942=>"101100100",
65943=>"001001000",
65944=>"110100110",
65945=>"001111011",
65946=>"001011011",
65947=>"010011010",
65948=>"100010000",
65949=>"010110110",
65950=>"100001100",
65951=>"110110111",
65952=>"000011000",
65953=>"111011011",
65954=>"000000001",
65955=>"000111100",
65956=>"101011110",
65957=>"111110111",
65958=>"100010000",
65959=>"100100000",
65960=>"011000011",
65961=>"011011011",
65962=>"011011011",
65963=>"010000110",
65964=>"000000101",
65965=>"100110110",
65966=>"111101111",
65967=>"000111100",
65968=>"111011001",
65969=>"000110110",
65970=>"101000000",
65971=>"111111111",
65972=>"000000001",
65973=>"001000001",
65974=>"000000000",
65975=>"100100000",
65976=>"011011011",
65977=>"001010111",
65978=>"001001100",
65979=>"101101100",
65980=>"010000000",
65981=>"101100110",
65982=>"001001001",
65983=>"011011011",
65984=>"111111110",
65985=>"110110101",
65986=>"000001111",
65987=>"000100100",
65988=>"011011011",
65989=>"110100000",
65990=>"111101001",
65991=>"000011000",
65992=>"100000101",
65993=>"000111110",
65994=>"101101000",
65995=>"011111100",
65996=>"011010010",
65997=>"111111010",
65998=>"100100100",
65999=>"000011011",
66000=>"100100111",
66001=>"100100100",
66002=>"111001101",
66003=>"100100000",
66004=>"110100100",
66005=>"110101000",
66006=>"101111111",
66007=>"000000111",
66008=>"011011001",
66009=>"100010000",
66010=>"111011101",
66011=>"100100101",
66012=>"101100111",
66013=>"001010010",
66014=>"100000100",
66015=>"011011111",
66016=>"011011001",
66017=>"100100100",
66018=>"011011011",
66019=>"100110101",
66020=>"010011011",
66021=>"011011011",
66022=>"001000101",
66023=>"100110111",
66024=>"000000000",
66025=>"010111001",
66026=>"111101111",
66027=>"001110011",
66028=>"011011011",
66029=>"000101111",
66030=>"000000000",
66031=>"001011011",
66032=>"011001001",
66033=>"000110110",
66034=>"011010010",
66035=>"110111111",
66036=>"101001101",
66037=>"000110101",
66038=>"000010000",
66039=>"000011011",
66040=>"011011011",
66041=>"000000000",
66042=>"110010110",
66043=>"000010100",
66044=>"100100100",
66045=>"001000000",
66046=>"110100100",
66047=>"111111111",
66048=>"011101111",
66049=>"111100100",
66050=>"010010111",
66051=>"101111111",
66052=>"000000111",
66053=>"001111111",
66054=>"101111000",
66055=>"111111000",
66056=>"001000100",
66057=>"000111000",
66058=>"100001001",
66059=>"000011000",
66060=>"000110001",
66061=>"000000000",
66062=>"000110111",
66063=>"000100101",
66064=>"100101100",
66065=>"111111100",
66066=>"110100110",
66067=>"111000000",
66068=>"010000000",
66069=>"101000000",
66070=>"001100000",
66071=>"111010010",
66072=>"101101101",
66073=>"000110101",
66074=>"000000010",
66075=>"010111010",
66076=>"010111000",
66077=>"000000001",
66078=>"000010010",
66079=>"001000000",
66080=>"010111110",
66081=>"101111000",
66082=>"111111110",
66083=>"000000000",
66084=>"000000000",
66085=>"110110100",
66086=>"000000000",
66087=>"000101110",
66088=>"011101111",
66089=>"101000000",
66090=>"000000000",
66091=>"010101111",
66092=>"000011011",
66093=>"000001011",
66094=>"111010111",
66095=>"000000000",
66096=>"000100110",
66097=>"001001000",
66098=>"010000100",
66099=>"101011011",
66100=>"111111110",
66101=>"011110000",
66102=>"011000000",
66103=>"111100100",
66104=>"111111000",
66105=>"111101001",
66106=>"111010000",
66107=>"111111110",
66108=>"100110100",
66109=>"000111111",
66110=>"000010011",
66111=>"110010100",
66112=>"110110000",
66113=>"111010000",
66114=>"000000101",
66115=>"111001001",
66116=>"000000000",
66117=>"101000101",
66118=>"000000110",
66119=>"001100010",
66120=>"001000000",
66121=>"010111010",
66122=>"100000000",
66123=>"111010100",
66124=>"111100000",
66125=>"000000110",
66126=>"010011011",
66127=>"000011010",
66128=>"111000101",
66129=>"111111000",
66130=>"000111011",
66131=>"010111110",
66132=>"010010000",
66133=>"001000000",
66134=>"000110011",
66135=>"010111111",
66136=>"111111111",
66137=>"110111000",
66138=>"111111011",
66139=>"100110000",
66140=>"111111010",
66141=>"010011110",
66142=>"111101111",
66143=>"010100110",
66144=>"101100111",
66145=>"100101101",
66146=>"010111111",
66147=>"111111111",
66148=>"000111011",
66149=>"101111100",
66150=>"110111010",
66151=>"001000101",
66152=>"101111011",
66153=>"111111000",
66154=>"111111101",
66155=>"000010111",
66156=>"000000000",
66157=>"000000000",
66158=>"100111111",
66159=>"111111000",
66160=>"110110100",
66161=>"100111111",
66162=>"011000000",
66163=>"010010110",
66164=>"111111011",
66165=>"001000100",
66166=>"000111111",
66167=>"000100101",
66168=>"111111010",
66169=>"010000000",
66170=>"001000100",
66171=>"010101111",
66172=>"000100110",
66173=>"000010011",
66174=>"000000111",
66175=>"110111110",
66176=>"000111111",
66177=>"010110010",
66178=>"010111111",
66179=>"111111000",
66180=>"000100001",
66181=>"011011000",
66182=>"011011001",
66183=>"000100010",
66184=>"001111111",
66185=>"110000010",
66186=>"010011011",
66187=>"001101010",
66188=>"000000101",
66189=>"110111111",
66190=>"111101111",
66191=>"000000110",
66192=>"010000000",
66193=>"111101000",
66194=>"000101100",
66195=>"111000111",
66196=>"011011111",
66197=>"101111000",
66198=>"110111000",
66199=>"111110100",
66200=>"111111101",
66201=>"111000000",
66202=>"000110000",
66203=>"011111111",
66204=>"001000000",
66205=>"010111101",
66206=>"000101000",
66207=>"000110111",
66208=>"000110011",
66209=>"111111111",
66210=>"010000010",
66211=>"100000000",
66212=>"000000111",
66213=>"110011010",
66214=>"011001010",
66215=>"000110000",
66216=>"001101111",
66217=>"011101101",
66218=>"010000000",
66219=>"000111011",
66220=>"101111111",
66221=>"111111111",
66222=>"010110000",
66223=>"101001101",
66224=>"111011001",
66225=>"001101101",
66226=>"000111000",
66227=>"111111000",
66228=>"000111011",
66229=>"111111010",
66230=>"101111101",
66231=>"011111111",
66232=>"001001001",
66233=>"000100110",
66234=>"111000010",
66235=>"000111111",
66236=>"000010111",
66237=>"010111111",
66238=>"011100101",
66239=>"111100000",
66240=>"111101010",
66241=>"111000000",
66242=>"000100110",
66243=>"000011011",
66244=>"000011000",
66245=>"111011111",
66246=>"001111110",
66247=>"110111000",
66248=>"000101001",
66249=>"110100100",
66250=>"001101110",
66251=>"111100110",
66252=>"000000000",
66253=>"000000011",
66254=>"110010010",
66255=>"110101001",
66256=>"111111010",
66257=>"110011011",
66258=>"111011011",
66259=>"000000010",
66260=>"000011111",
66261=>"110001111",
66262=>"000010010",
66263=>"011001000",
66264=>"111111111",
66265=>"000001011",
66266=>"101011101",
66267=>"110010000",
66268=>"100110111",
66269=>"111101100",
66270=>"111100000",
66271=>"000000000",
66272=>"100111111",
66273=>"000111111",
66274=>"111000000",
66275=>"011111111",
66276=>"010010010",
66277=>"000000111",
66278=>"010111000",
66279=>"110010101",
66280=>"101101111",
66281=>"000100010",
66282=>"001001011",
66283=>"101111111",
66284=>"001001000",
66285=>"101000000",
66286=>"010110010",
66287=>"100011011",
66288=>"111000111",
66289=>"111100111",
66290=>"000111111",
66291=>"010010000",
66292=>"000000111",
66293=>"101000101",
66294=>"000001000",
66295=>"010000000",
66296=>"000000000",
66297=>"101001010",
66298=>"101100111",
66299=>"000111111",
66300=>"111001000",
66301=>"011000101",
66302=>"001110100",
66303=>"000010000",
66304=>"000011111",
66305=>"000000000",
66306=>"000000100",
66307=>"110111010",
66308=>"000000000",
66309=>"000010000",
66310=>"110000001",
66311=>"111110011",
66312=>"000111111",
66313=>"000000000",
66314=>"011001000",
66315=>"000000000",
66316=>"000000000",
66317=>"000111111",
66318=>"000011011",
66319=>"000000000",
66320=>"101111001",
66321=>"110000011",
66322=>"111000000",
66323=>"111111000",
66324=>"101010000",
66325=>"010011010",
66326=>"000000010",
66327=>"111111011",
66328=>"010010000",
66329=>"000110011",
66330=>"000111000",
66331=>"101111111",
66332=>"000001000",
66333=>"111000000",
66334=>"111011111",
66335=>"111000000",
66336=>"000111111",
66337=>"010010000",
66338=>"111001000",
66339=>"000011111",
66340=>"111101110",
66341=>"001110110",
66342=>"000111110",
66343=>"000110110",
66344=>"000010111",
66345=>"000111111",
66346=>"000000000",
66347=>"000010000",
66348=>"011001000",
66349=>"111000111",
66350=>"111111100",
66351=>"000001101",
66352=>"000000111",
66353=>"000011001",
66354=>"000111100",
66355=>"000000001",
66356=>"001000000",
66357=>"010000101",
66358=>"100100001",
66359=>"001101000",
66360=>"001000010",
66361=>"111000001",
66362=>"110101111",
66363=>"111101011",
66364=>"011000001",
66365=>"010111000",
66366=>"001000000",
66367=>"010111111",
66368=>"000110101",
66369=>"101101101",
66370=>"110111111",
66371=>"000110110",
66372=>"110000000",
66373=>"011001000",
66374=>"011100110",
66375=>"111001000",
66376=>"111100100",
66377=>"111111111",
66378=>"010100101",
66379=>"111101100",
66380=>"010000100",
66381=>"001001101",
66382=>"000100100",
66383=>"111101001",
66384=>"101101101",
66385=>"010011000",
66386=>"111111111",
66387=>"111001000",
66388=>"101000101",
66389=>"010100111",
66390=>"111011001",
66391=>"000111111",
66392=>"001111111",
66393=>"011101001",
66394=>"111100100",
66395=>"111111100",
66396=>"101010010",
66397=>"110001001",
66398=>"111000001",
66399=>"000011111",
66400=>"000010110",
66401=>"110000110",
66402=>"000000001",
66403=>"111100110",
66404=>"010111100",
66405=>"110111101",
66406=>"111111110",
66407=>"000001010",
66408=>"101100110",
66409=>"010111111",
66410=>"111111000",
66411=>"111111101",
66412=>"111111111",
66413=>"111100110",
66414=>"001101000",
66415=>"000000000",
66416=>"000110111",
66417=>"010011010",
66418=>"000001100",
66419=>"111000000",
66420=>"111001000",
66421=>"111001111",
66422=>"000001110",
66423=>"000111111",
66424=>"000001010",
66425=>"000111101",
66426=>"101000100",
66427=>"111101001",
66428=>"001010110",
66429=>"111101000",
66430=>"110110000",
66431=>"000000101",
66432=>"101000111",
66433=>"010100100",
66434=>"111111110",
66435=>"111101111",
66436=>"000100110",
66437=>"111111111",
66438=>"100111011",
66439=>"000010011",
66440=>"000001011",
66441=>"101101000",
66442=>"010000010",
66443=>"101101000",
66444=>"000000000",
66445=>"010110110",
66446=>"010000000",
66447=>"001101000",
66448=>"011001011",
66449=>"000100101",
66450=>"001101000",
66451=>"100011101",
66452=>"000110010",
66453=>"000011111",
66454=>"000000101",
66455=>"010110111",
66456=>"000000000",
66457=>"010000111",
66458=>"100000111",
66459=>"111100000",
66460=>"111010010",
66461=>"110011011",
66462=>"100000000",
66463=>"111101101",
66464=>"111000100",
66465=>"010000110",
66466=>"000111111",
66467=>"000011111",
66468=>"111111101",
66469=>"011001111",
66470=>"111001010",
66471=>"000101000",
66472=>"000100000",
66473=>"000111111",
66474=>"101111111",
66475=>"000000000",
66476=>"111101001",
66477=>"000111111",
66478=>"011001000",
66479=>"111111111",
66480=>"100101000",
66481=>"111110001",
66482=>"111000001",
66483=>"010110110",
66484=>"110000100",
66485=>"101000000",
66486=>"000000111",
66487=>"000010111",
66488=>"110000010",
66489=>"000110101",
66490=>"000000010",
66491=>"000010111",
66492=>"110010111",
66493=>"010111111",
66494=>"001011111",
66495=>"000000101",
66496=>"111000111",
66497=>"111011000",
66498=>"000001111",
66499=>"000110111",
66500=>"101000011",
66501=>"011000001",
66502=>"011000011",
66503=>"001000000",
66504=>"111111000",
66505=>"111100000",
66506=>"000001011",
66507=>"110100001",
66508=>"000011111",
66509=>"100010011",
66510=>"101000000",
66511=>"000111000",
66512=>"000010110",
66513=>"001000010",
66514=>"000010000",
66515=>"111000010",
66516=>"000111111",
66517=>"111000011",
66518=>"000000001",
66519=>"000111010",
66520=>"111100000",
66521=>"001000100",
66522=>"110001101",
66523=>"111000010",
66524=>"100001001",
66525=>"000000111",
66526=>"110100111",
66527=>"011111000",
66528=>"111000100",
66529=>"000000001",
66530=>"000111111",
66531=>"110111111",
66532=>"000010111",
66533=>"000000111",
66534=>"001111111",
66535=>"111111101",
66536=>"010111110",
66537=>"010111111",
66538=>"110100000",
66539=>"101000000",
66540=>"000000111",
66541=>"000110111",
66542=>"000010000",
66543=>"101000010",
66544=>"111000000",
66545=>"100000100",
66546=>"101111110",
66547=>"010001000",
66548=>"000100111",
66549=>"111000000",
66550=>"000000110",
66551=>"111100001",
66552=>"101000000",
66553=>"111000010",
66554=>"111111111",
66555=>"000000000",
66556=>"001000000",
66557=>"111011011",
66558=>"110101111",
66559=>"111110000",
66560=>"010001000",
66561=>"000111111",
66562=>"000000000",
66563=>"000000111",
66564=>"110110110",
66565=>"110111110",
66566=>"101111100",
66567=>"000001111",
66568=>"000000000",
66569=>"101101011",
66570=>"010011100",
66571=>"101000101",
66572=>"111111100",
66573=>"100000011",
66574=>"011100011",
66575=>"110000000",
66576=>"000000111",
66577=>"110010000",
66578=>"111000101",
66579=>"111101000",
66580=>"000000011",
66581=>"111111100",
66582=>"011110100",
66583=>"000001010",
66584=>"111000000",
66585=>"111111111",
66586=>"000001000",
66587=>"000000001",
66588=>"000000110",
66589=>"001101010",
66590=>"111100000",
66591=>"100111001",
66592=>"110111111",
66593=>"111111011",
66594=>"000010001",
66595=>"010010000",
66596=>"000001100",
66597=>"111111111",
66598=>"111100000",
66599=>"000110000",
66600=>"100011111",
66601=>"101101010",
66602=>"000000011",
66603=>"010101111",
66604=>"001001011",
66605=>"111110110",
66606=>"101111111",
66607=>"000000111",
66608=>"110001101",
66609=>"110110110",
66610=>"000010001",
66611=>"010010000",
66612=>"000001100",
66613=>"010000000",
66614=>"110110100",
66615=>"000000110",
66616=>"010101001",
66617=>"000000000",
66618=>"011100000",
66619=>"011010011",
66620=>"011011110",
66621=>"111111010",
66622=>"000000000",
66623=>"110110110",
66624=>"010101111",
66625=>"101111100",
66626=>"110111010",
66627=>"011001111",
66628=>"000110110",
66629=>"000110110",
66630=>"010000000",
66631=>"011000000",
66632=>"001000110",
66633=>"111010111",
66634=>"101100111",
66635=>"111000000",
66636=>"000011001",
66637=>"110110010",
66638=>"111111111",
66639=>"100110110",
66640=>"110010000",
66641=>"111000010",
66642=>"111000010",
66643=>"000000000",
66644=>"101001111",
66645=>"011010110",
66646=>"010011001",
66647=>"111001111",
66648=>"000000100",
66649=>"100100001",
66650=>"001101101",
66651=>"100000000",
66652=>"111100100",
66653=>"000001000",
66654=>"001100011",
66655=>"100101001",
66656=>"101010000",
66657=>"000001111",
66658=>"100010010",
66659=>"000000100",
66660=>"001001000",
66661=>"110000000",
66662=>"111011111",
66663=>"010001000",
66664=>"111010111",
66665=>"000000000",
66666=>"000010101",
66667=>"001011111",
66668=>"100001101",
66669=>"010111111",
66670=>"110010000",
66671=>"000000110",
66672=>"001000000",
66673=>"000111111",
66674=>"111011100",
66675=>"111110011",
66676=>"101110111",
66677=>"000000000",
66678=>"000111101",
66679=>"000000000",
66680=>"101101100",
66681=>"000010000",
66682=>"000110111",
66683=>"111000001",
66684=>"011100111",
66685=>"100000000",
66686=>"101001111",
66687=>"001000101",
66688=>"001001110",
66689=>"010000111",
66690=>"100000010",
66691=>"010101111",
66692=>"101101110",
66693=>"000000000",
66694=>"100011111",
66695=>"110100111",
66696=>"000101001",
66697=>"100000010",
66698=>"001101101",
66699=>"111100101",
66700=>"001001001",
66701=>"111111001",
66702=>"000000000",
66703=>"001000000",
66704=>"011001100",
66705=>"100101001",
66706=>"010001001",
66707=>"101001100",
66708=>"100010011",
66709=>"000110100",
66710=>"111010010",
66711=>"000001111",
66712=>"110110000",
66713=>"101100101",
66714=>"101101111",
66715=>"000000000",
66716=>"101000100",
66717=>"111010111",
66718=>"010000000",
66719=>"111011111",
66720=>"000111110",
66721=>"000000110",
66722=>"000011001",
66723=>"101000111",
66724=>"001000000",
66725=>"001011010",
66726=>"110110000",
66727=>"000000000",
66728=>"110011000",
66729=>"000000000",
66730=>"101101010",
66731=>"110010000",
66732=>"011111101",
66733=>"110110000",
66734=>"100001010",
66735=>"110010000",
66736=>"101000111",
66737=>"010001000",
66738=>"000001101",
66739=>"001100000",
66740=>"101101100",
66741=>"001100111",
66742=>"111111111",
66743=>"010111111",
66744=>"100011011",
66745=>"110010110",
66746=>"111000000",
66747=>"001000111",
66748=>"111110010",
66749=>"100010111",
66750=>"011000011",
66751=>"110100000",
66752=>"111001111",
66753=>"101111111",
66754=>"000111110",
66755=>"001100110",
66756=>"000010000",
66757=>"100100011",
66758=>"110100110",
66759=>"111111111",
66760=>"001110111",
66761=>"000101000",
66762=>"000111111",
66763=>"010111111",
66764=>"111101101",
66765=>"110011011",
66766=>"000010111",
66767=>"111111111",
66768=>"000001001",
66769=>"000000110",
66770=>"111001111",
66771=>"000111111",
66772=>"111011101",
66773=>"000000011",
66774=>"001000000",
66775=>"100000001",
66776=>"111101110",
66777=>"001000100",
66778=>"100000001",
66779=>"000000000",
66780=>"010011001",
66781=>"000101101",
66782=>"111111000",
66783=>"110010001",
66784=>"111110000",
66785=>"000010000",
66786=>"001000001",
66787=>"111111000",
66788=>"101000100",
66789=>"111111001",
66790=>"011001101",
66791=>"001011010",
66792=>"000110111",
66793=>"110110100",
66794=>"000000011",
66795=>"001111110",
66796=>"000000111",
66797=>"111101100",
66798=>"000000000",
66799=>"110110000",
66800=>"010100000",
66801=>"011011010",
66802=>"001000000",
66803=>"001001001",
66804=>"011010000",
66805=>"000000101",
66806=>"010010010",
66807=>"000000001",
66808=>"000000111",
66809=>"101001000",
66810=>"001101111",
66811=>"001001000",
66812=>"110110000",
66813=>"011011101",
66814=>"011010000",
66815=>"000000000",
66816=>"100100100",
66817=>"101000110",
66818=>"000000101",
66819=>"101000000",
66820=>"111101011",
66821=>"101101000",
66822=>"000000010",
66823=>"110111111",
66824=>"010000000",
66825=>"000000000",
66826=>"001110000",
66827=>"000101100",
66828=>"011000100",
66829=>"111111000",
66830=>"011000000",
66831=>"111100100",
66832=>"111000001",
66833=>"100000000",
66834=>"100101110",
66835=>"110111011",
66836=>"000101101",
66837=>"000111111",
66838=>"111011111",
66839=>"000110111",
66840=>"000000101",
66841=>"010111101",
66842=>"000000000",
66843=>"000000000",
66844=>"100000011",
66845=>"100010000",
66846=>"000001000",
66847=>"001111010",
66848=>"101000101",
66849=>"111111111",
66850=>"111101111",
66851=>"111110111",
66852=>"111000000",
66853=>"000011100",
66854=>"000010000",
66855=>"111111000",
66856=>"010111111",
66857=>"000001000",
66858=>"101101000",
66859=>"011111010",
66860=>"000100111",
66861=>"111010100",
66862=>"101110000",
66863=>"101111110",
66864=>"101011101",
66865=>"111000000",
66866=>"000111111",
66867=>"000100000",
66868=>"000010011",
66869=>"111111111",
66870=>"001011110",
66871=>"111010000",
66872=>"111100111",
66873=>"000101000",
66874=>"000100010",
66875=>"011000111",
66876=>"001011111",
66877=>"010111010",
66878=>"000000000",
66879=>"001100000",
66880=>"100000111",
66881=>"000100000",
66882=>"111110010",
66883=>"110100000",
66884=>"000000000",
66885=>"000101001",
66886=>"100101100",
66887=>"101100010",
66888=>"111111110",
66889=>"101101111",
66890=>"001010010",
66891=>"000000000",
66892=>"010000100",
66893=>"100100100",
66894=>"011000000",
66895=>"001000001",
66896=>"010010000",
66897=>"111010111",
66898=>"001000101",
66899=>"000000000",
66900=>"000000111",
66901=>"011010110",
66902=>"011000000",
66903=>"101100000",
66904=>"000000010",
66905=>"110000000",
66906=>"000011011",
66907=>"100000010",
66908=>"011000001",
66909=>"001001111",
66910=>"100101101",
66911=>"011001001",
66912=>"111000000",
66913=>"111110010",
66914=>"000000000",
66915=>"000110110",
66916=>"110000001",
66917=>"100000000",
66918=>"111100101",
66919=>"100000100",
66920=>"101111010",
66921=>"111111111",
66922=>"101101111",
66923=>"111000000",
66924=>"100010100",
66925=>"100011000",
66926=>"010000000",
66927=>"000101111",
66928=>"111000000",
66929=>"100101101",
66930=>"000111111",
66931=>"111000000",
66932=>"101001000",
66933=>"000000000",
66934=>"001001000",
66935=>"010000000",
66936=>"001000000",
66937=>"000100000",
66938=>"101100001",
66939=>"000000001",
66940=>"101100111",
66941=>"001001001",
66942=>"011111111",
66943=>"000001010",
66944=>"110101101",
66945=>"000111011",
66946=>"000000111",
66947=>"101001100",
66948=>"000000101",
66949=>"101111010",
66950=>"000110000",
66951=>"011001000",
66952=>"111000100",
66953=>"000110010",
66954=>"000000000",
66955=>"010000000",
66956=>"101000100",
66957=>"101101000",
66958=>"111010100",
66959=>"010000000",
66960=>"110101001",
66961=>"000001000",
66962=>"000000000",
66963=>"000100111",
66964=>"101100000",
66965=>"101000101",
66966=>"111111011",
66967=>"000101100",
66968=>"100000000",
66969=>"000110010",
66970=>"000011111",
66971=>"111000001",
66972=>"011000000",
66973=>"101111111",
66974=>"101111111",
66975=>"010101101",
66976=>"111111111",
66977=>"000010011",
66978=>"011111011",
66979=>"111111011",
66980=>"001101000",
66981=>"011000000",
66982=>"111101000",
66983=>"111111111",
66984=>"110110000",
66985=>"010011000",
66986=>"110111111",
66987=>"101100010",
66988=>"011000000",
66989=>"110100100",
66990=>"001111110",
66991=>"011101101",
66992=>"100000101",
66993=>"111011011",
66994=>"001111111",
66995=>"100100111",
66996=>"101001011",
66997=>"100100111",
66998=>"001001111",
66999=>"111001000",
67000=>"010111110",
67001=>"111010000",
67002=>"010111111",
67003=>"011010000",
67004=>"101011011",
67005=>"111111111",
67006=>"000100100",
67007=>"011011000",
67008=>"000000101",
67009=>"101100001",
67010=>"111111000",
67011=>"110000001",
67012=>"000000000",
67013=>"001101000",
67014=>"110100000",
67015=>"101010010",
67016=>"111010111",
67017=>"111001000",
67018=>"111010011",
67019=>"101101000",
67020=>"111100000",
67021=>"011011110",
67022=>"000000000",
67023=>"001000000",
67024=>"000001001",
67025=>"111011000",
67026=>"011001010",
67027=>"111101000",
67028=>"111101111",
67029=>"110111111",
67030=>"010011000",
67031=>"001001000",
67032=>"000000000",
67033=>"101111111",
67034=>"011001100",
67035=>"001101001",
67036=>"110101110",
67037=>"111111000",
67038=>"001000110",
67039=>"000000000",
67040=>"111000000",
67041=>"000001010",
67042=>"000101111",
67043=>"010001000",
67044=>"000000001",
67045=>"001101101",
67046=>"000000000",
67047=>"000101011",
67048=>"111000111",
67049=>"101111111",
67050=>"000010000",
67051=>"001000000",
67052=>"111111001",
67053=>"111111010",
67054=>"010000010",
67055=>"001101100",
67056=>"100000000",
67057=>"100100000",
67058=>"101101100",
67059=>"011100110",
67060=>"001001001",
67061=>"001111010",
67062=>"010010000",
67063=>"111101011",
67064=>"000000111",
67065=>"000111111",
67066=>"100101011",
67067=>"101010000",
67068=>"111111111",
67069=>"011111101",
67070=>"000001111",
67071=>"100000000",
67072=>"001000001",
67073=>"100000100",
67074=>"101101111",
67075=>"110010110",
67076=>"110100100",
67077=>"100001000",
67078=>"111011010",
67079=>"111111010",
67080=>"000000000",
67081=>"010010000",
67082=>"001001011",
67083=>"101101101",
67084=>"110000001",
67085=>"110011000",
67086=>"100100010",
67087=>"010110011",
67088=>"011000000",
67089=>"010010000",
67090=>"010100101",
67091=>"111011000",
67092=>"010111001",
67093=>"100100101",
67094=>"101101101",
67095=>"101101110",
67096=>"010010010",
67097=>"110100001",
67098=>"110110111",
67099=>"101100000",
67100=>"011011000",
67101=>"001001001",
67102=>"110010000",
67103=>"111011010",
67104=>"001101111",
67105=>"010000111",
67106=>"110111111",
67107=>"000000000",
67108=>"011011111",
67109=>"100100000",
67110=>"000000000",
67111=>"111111111",
67112=>"010111011",
67113=>"100111110",
67114=>"100000000",
67115=>"111111111",
67116=>"100010010",
67117=>"100101001",
67118=>"000000011",
67119=>"100000010",
67120=>"000010010",
67121=>"101101101",
67122=>"111000000",
67123=>"111100100",
67124=>"000000100",
67125=>"111101000",
67126=>"000100100",
67127=>"111011110",
67128=>"101101101",
67129=>"111100110",
67130=>"000000101",
67131=>"111111010",
67132=>"110110100",
67133=>"111111111",
67134=>"000100101",
67135=>"101101100",
67136=>"000010010",
67137=>"010100010",
67138=>"101111111",
67139=>"111001001",
67140=>"010010000",
67141=>"010000000",
67142=>"100000000",
67143=>"011110110",
67144=>"001100110",
67145=>"111010010",
67146=>"000001001",
67147=>"111000000",
67148=>"110000000",
67149=>"011110110",
67150=>"111111000",
67151=>"101111011",
67152=>"100100000",
67153=>"111111111",
67154=>"011001100",
67155=>"000001111",
67156=>"110100110",
67157=>"111101111",
67158=>"000100100",
67159=>"100100101",
67160=>"101000000",
67161=>"011100001",
67162=>"010000010",
67163=>"000000101",
67164=>"010111010",
67165=>"010001101",
67166=>"100000000",
67167=>"100000100",
67168=>"000110000",
67169=>"001001000",
67170=>"111101101",
67171=>"000110110",
67172=>"001000100",
67173=>"000000000",
67174=>"111101111",
67175=>"110101111",
67176=>"111110110",
67177=>"000010110",
67178=>"000000000",
67179=>"111001001",
67180=>"000000011",
67181=>"111111110",
67182=>"000000111",
67183=>"000000001",
67184=>"001100000",
67185=>"100101101",
67186=>"000001001",
67187=>"101011001",
67188=>"010011010",
67189=>"000000000",
67190=>"000010000",
67191=>"101011000",
67192=>"000000101",
67193=>"111111000",
67194=>"100101111",
67195=>"000001111",
67196=>"100000111",
67197=>"001010100",
67198=>"101100110",
67199=>"001101001",
67200=>"101000010",
67201=>"111011010",
67202=>"010111000",
67203=>"001111011",
67204=>"001000110",
67205=>"110100000",
67206=>"001001001",
67207=>"100101011",
67208=>"100110100",
67209=>"000000000",
67210=>"000110000",
67211=>"000000001",
67212=>"110110101",
67213=>"111111000",
67214=>"111111111",
67215=>"001000000",
67216=>"000100111",
67217=>"111100100",
67218=>"010000011",
67219=>"110010110",
67220=>"001011010",
67221=>"101100111",
67222=>"000010000",
67223=>"110000111",
67224=>"010010110",
67225=>"110111111",
67226=>"000000000",
67227=>"011111111",
67228=>"000000010",
67229=>"111001111",
67230=>"010011000",
67231=>"000000000",
67232=>"000000011",
67233=>"010100011",
67234=>"000101011",
67235=>"010110010",
67236=>"001111011",
67237=>"000000100",
67238=>"010110001",
67239=>"100000000",
67240=>"110010000",
67241=>"110111100",
67242=>"000000000",
67243=>"000011010",
67244=>"111101101",
67245=>"000101111",
67246=>"111110110",
67247=>"000110000",
67248=>"101000101",
67249=>"001000110",
67250=>"111101111",
67251=>"000001000",
67252=>"011111110",
67253=>"000010011",
67254=>"010011010",
67255=>"101100001",
67256=>"111001001",
67257=>"000000110",
67258=>"000010010",
67259=>"000010110",
67260=>"101001011",
67261=>"111111111",
67262=>"000000000",
67263=>"001000100",
67264=>"101000100",
67265=>"000000010",
67266=>"000000000",
67267=>"101100000",
67268=>"100010011",
67269=>"100100011",
67270=>"000000011",
67271=>"000000000",
67272=>"100111100",
67273=>"001000000",
67274=>"000100010",
67275=>"000000000",
67276=>"010100000",
67277=>"111010110",
67278=>"000100110",
67279=>"110110100",
67280=>"111001010",
67281=>"101000011",
67282=>"111100000",
67283=>"000011111",
67284=>"111000001",
67285=>"101101111",
67286=>"101111111",
67287=>"010000010",
67288=>"101000101",
67289=>"000001100",
67290=>"000111110",
67291=>"111100000",
67292=>"111111101",
67293=>"000111111",
67294=>"111000111",
67295=>"000000000",
67296=>"111101101",
67297=>"101000000",
67298=>"111011000",
67299=>"011011111",
67300=>"000000000",
67301=>"111100000",
67302=>"000000000",
67303=>"010010110",
67304=>"001111010",
67305=>"000010000",
67306=>"111100111",
67307=>"000000111",
67308=>"000000000",
67309=>"111111110",
67310=>"111111000",
67311=>"000010010",
67312=>"111101100",
67313=>"011101111",
67314=>"000000101",
67315=>"111110000",
67316=>"000001100",
67317=>"101100111",
67318=>"000000000",
67319=>"101111001",
67320=>"000000000",
67321=>"001010111",
67322=>"011001011",
67323=>"011111111",
67324=>"000000101",
67325=>"101111101",
67326=>"001011001",
67327=>"011111111",
67328=>"001001011",
67329=>"000000000",
67330=>"101100000",
67331=>"110111111",
67332=>"101100101",
67333=>"111101000",
67334=>"000111010",
67335=>"110111010",
67336=>"000000101",
67337=>"111101000",
67338=>"111100000",
67339=>"000000111",
67340=>"111100101",
67341=>"000000111",
67342=>"000100110",
67343=>"010010010",
67344=>"111101001",
67345=>"010010000",
67346=>"101111010",
67347=>"000001010",
67348=>"100000000",
67349=>"001000000",
67350=>"111110000",
67351=>"001111111",
67352=>"101101101",
67353=>"000000000",
67354=>"000011111",
67355=>"000000111",
67356=>"000011001",
67357=>"110111011",
67358=>"111100101",
67359=>"000010010",
67360=>"011010101",
67361=>"000111101",
67362=>"110111010",
67363=>"001010111",
67364=>"100101011",
67365=>"000000000",
67366=>"010111000",
67367=>"000000000",
67368=>"001111111",
67369=>"010111111",
67370=>"000000100",
67371=>"110110010",
67372=>"000110000",
67373=>"111110000",
67374=>"010011001",
67375=>"000000001",
67376=>"000101101",
67377=>"100001011",
67378=>"111111111",
67379=>"000111111",
67380=>"101011111",
67381=>"111010100",
67382=>"010000000",
67383=>"100100011",
67384=>"010011101",
67385=>"101000000",
67386=>"000010111",
67387=>"010010011",
67388=>"001000010",
67389=>"101111111",
67390=>"101101000",
67391=>"001000001",
67392=>"111101010",
67393=>"010000101",
67394=>"111111110",
67395=>"011001100",
67396=>"111000010",
67397=>"000000101",
67398=>"110111110",
67399=>"111110111",
67400=>"111111100",
67401=>"000010101",
67402=>"111001001",
67403=>"000110111",
67404=>"011111000",
67405=>"000000110",
67406=>"001000111",
67407=>"000010111",
67408=>"000111111",
67409=>"010111010",
67410=>"000011111",
67411=>"001001001",
67412=>"000000111",
67413=>"011011000",
67414=>"001111111",
67415=>"111101101",
67416=>"100010110",
67417=>"000010010",
67418=>"000011011",
67419=>"000000011",
67420=>"000010000",
67421=>"100111111",
67422=>"111111001",
67423=>"100100110",
67424=>"101001000",
67425=>"110110010",
67426=>"111101100",
67427=>"000110110",
67428=>"000001111",
67429=>"000011011",
67430=>"000000111",
67431=>"111000000",
67432=>"000010010",
67433=>"111101101",
67434=>"000101100",
67435=>"011111010",
67436=>"000010010",
67437=>"000101000",
67438=>"101111101",
67439=>"000111111",
67440=>"000000110",
67441=>"000100101",
67442=>"000001001",
67443=>"111001000",
67444=>"111011000",
67445=>"000001111",
67446=>"000000000",
67447=>"111101101",
67448=>"010010000",
67449=>"000010010",
67450=>"101111111",
67451=>"000000000",
67452=>"000010010",
67453=>"000100110",
67454=>"000011010",
67455=>"101001010",
67456=>"000001001",
67457=>"110111100",
67458=>"011000111",
67459=>"000001000",
67460=>"100101111",
67461=>"111111100",
67462=>"100000100",
67463=>"100001111",
67464=>"001101110",
67465=>"111000110",
67466=>"111111000",
67467=>"111000000",
67468=>"111101111",
67469=>"111000000",
67470=>"000010011",
67471=>"100000000",
67472=>"000111111",
67473=>"101000010",
67474=>"001000000",
67475=>"101111111",
67476=>"000001011",
67477=>"111101101",
67478=>"111110000",
67479=>"000100111",
67480=>"010011010",
67481=>"101001000",
67482=>"001101111",
67483=>"010111101",
67484=>"000111111",
67485=>"000000101",
67486=>"111011111",
67487=>"101101000",
67488=>"101011001",
67489=>"010111111",
67490=>"000110010",
67491=>"000000010",
67492=>"001011100",
67493=>"000100100",
67494=>"000001000",
67495=>"000000111",
67496=>"000000101",
67497=>"010000010",
67498=>"010111111",
67499=>"000111110",
67500=>"010110111",
67501=>"111101100",
67502=>"100111110",
67503=>"000011111",
67504=>"000110111",
67505=>"000111011",
67506=>"010000110",
67507=>"001101001",
67508=>"000000000",
67509=>"000001011",
67510=>"011100001",
67511=>"000110111",
67512=>"000000000",
67513=>"001001011",
67514=>"010111000",
67515=>"000010000",
67516=>"010010011",
67517=>"111001111",
67518=>"110101101",
67519=>"011111111",
67520=>"111111100",
67521=>"110110011",
67522=>"111111101",
67523=>"101001111",
67524=>"100000010",
67525=>"111111101",
67526=>"001111011",
67527=>"111101000",
67528=>"111001111",
67529=>"111011111",
67530=>"101000110",
67531=>"101000010",
67532=>"000000111",
67533=>"100010010",
67534=>"100111111",
67535=>"000000100",
67536=>"111101000",
67537=>"000101110",
67538=>"100000111",
67539=>"010010000",
67540=>"101101111",
67541=>"001111010",
67542=>"000010001",
67543=>"010110111",
67544=>"000010011",
67545=>"000000010",
67546=>"011111110",
67547=>"111101101",
67548=>"111011010",
67549=>"101101111",
67550=>"010000010",
67551=>"110110111",
67552=>"101000001",
67553=>"111111101",
67554=>"111111100",
67555=>"110011011",
67556=>"100000100",
67557=>"010010000",
67558=>"000000110",
67559=>"000110110",
67560=>"010111111",
67561=>"000011000",
67562=>"011101001",
67563=>"000101110",
67564=>"111101001",
67565=>"111111011",
67566=>"110111000",
67567=>"000000100",
67568=>"001000011",
67569=>"100010001",
67570=>"001111111",
67571=>"000110000",
67572=>"000010110",
67573=>"101100111",
67574=>"111000100",
67575=>"000100100",
67576=>"000101111",
67577=>"100111111",
67578=>"100111100",
67579=>"101111001",
67580=>"100010111",
67581=>"000010000",
67582=>"110000111",
67583=>"000011011",
67584=>"000100001",
67585=>"111111000",
67586=>"000000100",
67587=>"000000000",
67588=>"011111111",
67589=>"101000101",
67590=>"110101101",
67591=>"000111010",
67592=>"000000010",
67593=>"101101101",
67594=>"100000001",
67595=>"000010110",
67596=>"100000000",
67597=>"000101000",
67598=>"001011001",
67599=>"000010001",
67600=>"000010111",
67601=>"111101111",
67602=>"000100000",
67603=>"011100000",
67604=>"111111111",
67605=>"110100000",
67606=>"111011011",
67607=>"111000111",
67608=>"010101000",
67609=>"101110010",
67610=>"011001000",
67611=>"000000000",
67612=>"111111110",
67613=>"100100001",
67614=>"111000100",
67615=>"000100000",
67616=>"000101100",
67617=>"111100000",
67618=>"000100010",
67619=>"000010010",
67620=>"111001011",
67621=>"111011000",
67622=>"000000000",
67623=>"001000110",
67624=>"010111011",
67625=>"100110010",
67626=>"000000000",
67627=>"100011010",
67628=>"010101110",
67629=>"111101000",
67630=>"101101101",
67631=>"111101010",
67632=>"111000100",
67633=>"111111111",
67634=>"101111010",
67635=>"100000111",
67636=>"110100001",
67637=>"010111010",
67638=>"110000001",
67639=>"000001111",
67640=>"010010011",
67641=>"010000101",
67642=>"101101000",
67643=>"000000100",
67644=>"110010100",
67645=>"110101000",
67646=>"101100000",
67647=>"011001000",
67648=>"000011011",
67649=>"111010100",
67650=>"111111000",
67651=>"110000001",
67652=>"010000111",
67653=>"001011011",
67654=>"101001101",
67655=>"111001001",
67656=>"111001100",
67657=>"100000101",
67658=>"010000000",
67659=>"101000001",
67660=>"111101100",
67661=>"111110110",
67662=>"110111111",
67663=>"010010010",
67664=>"000000000",
67665=>"111000000",
67666=>"001101111",
67667=>"011000111",
67668=>"100111101",
67669=>"110100000",
67670=>"000000110",
67671=>"111000000",
67672=>"101101001",
67673=>"111000100",
67674=>"100110000",
67675=>"010011100",
67676=>"111010110",
67677=>"001001000",
67678=>"100111010",
67679=>"000001100",
67680=>"011111111",
67681=>"111000000",
67682=>"111000000",
67683=>"000111010",
67684=>"000110000",
67685=>"100011011",
67686=>"111111101",
67687=>"000111001",
67688=>"000000111",
67689=>"101100101",
67690=>"100000111",
67691=>"000000000",
67692=>"010110011",
67693=>"000010000",
67694=>"111100101",
67695=>"011001100",
67696=>"110110011",
67697=>"000000101",
67698=>"001000100",
67699=>"000001000",
67700=>"100000000",
67701=>"101101101",
67702=>"101101100",
67703=>"111110100",
67704=>"101001000",
67705=>"010000100",
67706=>"001111111",
67707=>"101101111",
67708=>"000111010",
67709=>"110100100",
67710=>"011000000",
67711=>"010000100",
67712=>"010010000",
67713=>"101000000",
67714=>"111111110",
67715=>"000000100",
67716=>"000011101",
67717=>"101111001",
67718=>"111010000",
67719=>"000001001",
67720=>"110001010",
67721=>"000000001",
67722=>"000101000",
67723=>"000111000",
67724=>"000010110",
67725=>"100000111",
67726=>"110000011",
67727=>"100000001",
67728=>"001011111",
67729=>"110100010",
67730=>"001000000",
67731=>"000011011",
67732=>"000000010",
67733=>"101000000",
67734=>"111101111",
67735=>"000011011",
67736=>"111110111",
67737=>"101001000",
67738=>"111000111",
67739=>"101100101",
67740=>"111000100",
67741=>"111100000",
67742=>"111000011",
67743=>"111101000",
67744=>"011011001",
67745=>"011000010",
67746=>"010001001",
67747=>"000101100",
67748=>"010000110",
67749=>"000110100",
67750=>"100110000",
67751=>"010001000",
67752=>"111111101",
67753=>"000000111",
67754=>"011100000",
67755=>"011000000",
67756=>"000101101",
67757=>"111000000",
67758=>"110001001",
67759=>"111111111",
67760=>"101111010",
67761=>"000001100",
67762=>"110001010",
67763=>"001100100",
67764=>"000001001",
67765=>"000100000",
67766=>"000011111",
67767=>"010011010",
67768=>"011011000",
67769=>"000000000",
67770=>"100100000",
67771=>"111101101",
67772=>"000101101",
67773=>"111111111",
67774=>"111100010",
67775=>"000010001",
67776=>"111100101",
67777=>"111101101",
67778=>"101000000",
67779=>"101110111",
67780=>"000000000",
67781=>"110110001",
67782=>"000000110",
67783=>"000000111",
67784=>"000000101",
67785=>"000111010",
67786=>"000111111",
67787=>"000011001",
67788=>"000000010",
67789=>"000111111",
67790=>"000111000",
67791=>"000111110",
67792=>"100100000",
67793=>"000110111",
67794=>"000010000",
67795=>"000000101",
67796=>"111000010",
67797=>"000001000",
67798=>"111000100",
67799=>"000000111",
67800=>"000000010",
67801=>"000011011",
67802=>"110110110",
67803=>"001000000",
67804=>"111110010",
67805=>"100111000",
67806=>"100011111",
67807=>"001000101",
67808=>"000000000",
67809=>"111100100",
67810=>"000010110",
67811=>"100000011",
67812=>"101000101",
67813=>"111101111",
67814=>"111101111",
67815=>"011111110",
67816=>"111111111",
67817=>"100111001",
67818=>"011100100",
67819=>"000000110",
67820=>"010111000",
67821=>"010010101",
67822=>"000000000",
67823=>"011110110",
67824=>"000001111",
67825=>"011011100",
67826=>"000010001",
67827=>"110101101",
67828=>"110001110",
67829=>"001101000",
67830=>"000000101",
67831=>"101100101",
67832=>"000000010",
67833=>"001101011",
67834=>"111001101",
67835=>"000000001",
67836=>"110001111",
67837=>"001000000",
67838=>"110011111",
67839=>"111101101",
67840=>"000110111",
67841=>"000000000",
67842=>"101111111",
67843=>"000111000",
67844=>"000100001",
67845=>"000111110",
67846=>"000000010",
67847=>"111000100",
67848=>"110111001",
67849=>"010111011",
67850=>"111111011",
67851=>"111011000",
67852=>"111111111",
67853=>"000110110",
67854=>"111111111",
67855=>"001111111",
67856=>"111111001",
67857=>"111100000",
67858=>"111111110",
67859=>"000000001",
67860=>"000000111",
67861=>"000000000",
67862=>"000000000",
67863=>"110111011",
67864=>"111111011",
67865=>"101001001",
67866=>"000000000",
67867=>"101111111",
67868=>"111111111",
67869=>"111111101",
67870=>"111111111",
67871=>"111000011",
67872=>"111110111",
67873=>"000010000",
67874=>"111111111",
67875=>"110111010",
67876=>"000000000",
67877=>"001011011",
67878=>"110111111",
67879=>"000111111",
67880=>"000000101",
67881=>"000000111",
67882=>"101111000",
67883=>"100000101",
67884=>"100000100",
67885=>"001101001",
67886=>"000111001",
67887=>"111000000",
67888=>"011111000",
67889=>"001000110",
67890=>"001000011",
67891=>"000000101",
67892=>"100110111",
67893=>"001000111",
67894=>"111110000",
67895=>"000000000",
67896=>"111000101",
67897=>"111111111",
67898=>"000000111",
67899=>"110101011",
67900=>"010110111",
67901=>"011010010",
67902=>"000000000",
67903=>"111011011",
67904=>"001101001",
67905=>"110111111",
67906=>"000000001",
67907=>"100111011",
67908=>"000000001",
67909=>"111101101",
67910=>"000001111",
67911=>"101001000",
67912=>"011011111",
67913=>"111111111",
67914=>"111001111",
67915=>"111111010",
67916=>"110000000",
67917=>"001000011",
67918=>"000000000",
67919=>"001000101",
67920=>"011111001",
67921=>"111010000",
67922=>"000101100",
67923=>"110100010",
67924=>"111000010",
67925=>"010011011",
67926=>"000001001",
67927=>"111111111",
67928=>"000000100",
67929=>"000000000",
67930=>"000000000",
67931=>"111010000",
67932=>"111111000",
67933=>"010110010",
67934=>"100111111",
67935=>"011111110",
67936=>"000000000",
67937=>"111110010",
67938=>"000010000",
67939=>"100000000",
67940=>"111000011",
67941=>"100100010",
67942=>"111111111",
67943=>"111111111",
67944=>"001000000",
67945=>"100111111",
67946=>"001101000",
67947=>"111111101",
67948=>"000001001",
67949=>"010010010",
67950=>"001111000",
67951=>"000000111",
67952=>"011000011",
67953=>"000000000",
67954=>"110111001",
67955=>"111110111",
67956=>"000000110",
67957=>"101000000",
67958=>"000000001",
67959=>"000000001",
67960=>"000101000",
67961=>"000111111",
67962=>"101101001",
67963=>"000010010",
67964=>"001001011",
67965=>"011011010",
67966=>"001111001",
67967=>"111111111",
67968=>"000101101",
67969=>"011011111",
67970=>"111111000",
67971=>"110010000",
67972=>"000000000",
67973=>"111111111",
67974=>"110010111",
67975=>"001000111",
67976=>"111001110",
67977=>"000000000",
67978=>"010111111",
67979=>"000101010",
67980=>"000111111",
67981=>"000001000",
67982=>"111111111",
67983=>"100000000",
67984=>"010000001",
67985=>"101101111",
67986=>"110100000",
67987=>"000000000",
67988=>"001011111",
67989=>"111111101",
67990=>"000111111",
67991=>"110010000",
67992=>"000000000",
67993=>"000100000",
67994=>"111111000",
67995=>"010111000",
67996=>"101011010",
67997=>"000000000",
67998=>"100000010",
67999=>"110110010",
68000=>"000100111",
68001=>"111101000",
68002=>"000000111",
68003=>"111111010",
68004=>"101001100",
68005=>"000000000",
68006=>"101111111",
68007=>"110111111",
68008=>"001101000",
68009=>"000000001",
68010=>"001000000",
68011=>"110111000",
68012=>"000000000",
68013=>"100000000",
68014=>"010011001",
68015=>"001000000",
68016=>"111101111",
68017=>"110000111",
68018=>"100111111",
68019=>"100100000",
68020=>"111111111",
68021=>"011011011",
68022=>"000100000",
68023=>"101101111",
68024=>"100011111",
68025=>"100001101",
68026=>"111111100",
68027=>"111111010",
68028=>"000000110",
68029=>"000111111",
68030=>"011100100",
68031=>"001000000",
68032=>"010111111",
68033=>"111011000",
68034=>"101111101",
68035=>"101000010",
68036=>"001001010",
68037=>"001001011",
68038=>"111101000",
68039=>"111111111",
68040=>"110001111",
68041=>"111010110",
68042=>"010111000",
68043=>"101101111",
68044=>"111111010",
68045=>"101100100",
68046=>"000000000",
68047=>"000010000",
68048=>"110110010",
68049=>"010010011",
68050=>"100101001",
68051=>"000101111",
68052=>"111111000",
68053=>"101011100",
68054=>"010111111",
68055=>"110000000",
68056=>"001000111",
68057=>"000100001",
68058=>"011001000",
68059=>"000111111",
68060=>"001000001",
68061=>"111110101",
68062=>"000000000",
68063=>"001101000",
68064=>"000000000",
68065=>"111010101",
68066=>"001000101",
68067=>"100000000",
68068=>"000110010",
68069=>"001001111",
68070=>"110110010",
68071=>"000010100",
68072=>"000111000",
68073=>"100000000",
68074=>"111111110",
68075=>"111111111",
68076=>"101101111",
68077=>"001000101",
68078=>"110111111",
68079=>"010111110",
68080=>"111110110",
68081=>"100100101",
68082=>"101111111",
68083=>"010010001",
68084=>"110101110",
68085=>"100100101",
68086=>"110000000",
68087=>"111001111",
68088=>"111001011",
68089=>"101000010",
68090=>"110111111",
68091=>"010111111",
68092=>"011011000",
68093=>"000110111",
68094=>"000000000",
68095=>"111000000",
68096=>"011011000",
68097=>"001000000",
68098=>"000000001",
68099=>"101110110",
68100=>"100111011",
68101=>"110100000",
68102=>"111010011",
68103=>"000010010",
68104=>"001111100",
68105=>"001000110",
68106=>"101000000",
68107=>"111000000",
68108=>"010111000",
68109=>"000001000",
68110=>"100011011",
68111=>"110100111",
68112=>"111110111",
68113=>"000000000",
68114=>"000000000",
68115=>"000000010",
68116=>"111001001",
68117=>"000101101",
68118=>"000101101",
68119=>"000000110",
68120=>"100111110",
68121=>"000110111",
68122=>"000101000",
68123=>"111101000",
68124=>"000000000",
68125=>"001000111",
68126=>"110000110",
68127=>"000001000",
68128=>"100000011",
68129=>"010111010",
68130=>"101000001",
68131=>"000010000",
68132=>"110111001",
68133=>"111111101",
68134=>"111000111",
68135=>"011110000",
68136=>"111111111",
68137=>"111010010",
68138=>"000010010",
68139=>"111011111",
68140=>"011001011",
68141=>"000101010",
68142=>"011000101",
68143=>"000000110",
68144=>"000001010",
68145=>"101011011",
68146=>"000000000",
68147=>"101000111",
68148=>"111000001",
68149=>"111111000",
68150=>"100100001",
68151=>"000000001",
68152=>"100000100",
68153=>"111001000",
68154=>"011100010",
68155=>"011001000",
68156=>"110110000",
68157=>"001101000",
68158=>"000000000",
68159=>"011010000",
68160=>"111111000",
68161=>"111101101",
68162=>"110111010",
68163=>"001100000",
68164=>"000000110",
68165=>"111000101",
68166=>"011001001",
68167=>"011111111",
68168=>"000000000",
68169=>"110010010",
68170=>"111000101",
68171=>"000110000",
68172=>"010000000",
68173=>"000100100",
68174=>"001101100",
68175=>"111111111",
68176=>"000001000",
68177=>"111111001",
68178=>"000001000",
68179=>"001000000",
68180=>"110000101",
68181=>"000000001",
68182=>"000101100",
68183=>"000000000",
68184=>"110100001",
68185=>"111111011",
68186=>"010100000",
68187=>"110111000",
68188=>"111011000",
68189=>"001001011",
68190=>"111111111",
68191=>"001101001",
68192=>"101000000",
68193=>"111111010",
68194=>"101000111",
68195=>"000011000",
68196=>"000111000",
68197=>"111100100",
68198=>"111111000",
68199=>"111111101",
68200=>"000000000",
68201=>"111111000",
68202=>"111110110",
68203=>"111111111",
68204=>"000000111",
68205=>"000001010",
68206=>"111110100",
68207=>"000001001",
68208=>"111001000",
68209=>"010110111",
68210=>"001000100",
68211=>"101010111",
68212=>"001011000",
68213=>"100100000",
68214=>"000110110",
68215=>"111010001",
68216=>"101111101",
68217=>"110101000",
68218=>"000000000",
68219=>"001101111",
68220=>"000110110",
68221=>"100100001",
68222=>"101111110",
68223=>"000000000",
68224=>"111111000",
68225=>"111000001",
68226=>"010000000",
68227=>"111111111",
68228=>"000101000",
68229=>"001000000",
68230=>"011101010",
68231=>"011011000",
68232=>"000101000",
68233=>"001110001",
68234=>"111111011",
68235=>"010010111",
68236=>"001000101",
68237=>"001001111",
68238=>"001000000",
68239=>"011000001",
68240=>"011001101",
68241=>"111000000",
68242=>"000000101",
68243=>"001000100",
68244=>"000110111",
68245=>"000000111",
68246=>"010111101",
68247=>"110000001",
68248=>"111111000",
68249=>"111001110",
68250=>"000000000",
68251=>"101000000",
68252=>"000000010",
68253=>"000000001",
68254=>"110001000",
68255=>"001000011",
68256=>"000000001",
68257=>"111111011",
68258=>"001010010",
68259=>"111111000",
68260=>"000000001",
68261=>"110110000",
68262=>"001001101",
68263=>"111110111",
68264=>"000000011",
68265=>"111010111",
68266=>"111111111",
68267=>"000000000",
68268=>"011000100",
68269=>"111111000",
68270=>"100000001",
68271=>"000101011",
68272=>"010000010",
68273=>"000000000",
68274=>"010001111",
68275=>"001100100",
68276=>"100101010",
68277=>"000000011",
68278=>"010110011",
68279=>"111110111",
68280=>"011011100",
68281=>"000111110",
68282=>"111101010",
68283=>"001001111",
68284=>"110110000",
68285=>"001001001",
68286=>"101110000",
68287=>"001001101",
68288=>"110101000",
68289=>"010010000",
68290=>"111000000",
68291=>"101011000",
68292=>"011010010",
68293=>"001001111",
68294=>"000100111",
68295=>"110110000",
68296=>"111110010",
68297=>"001001001",
68298=>"110111100",
68299=>"110110111",
68300=>"110010000",
68301=>"000011011",
68302=>"010000000",
68303=>"111111101",
68304=>"000000010",
68305=>"011100010",
68306=>"111111010",
68307=>"110110010",
68308=>"000000001",
68309=>"101000000",
68310=>"111111000",
68311=>"001101010",
68312=>"000001001",
68313=>"011000000",
68314=>"110100001",
68315=>"000000111",
68316=>"001100011",
68317=>"011011111",
68318=>"010100101",
68319=>"000010111",
68320=>"110111001",
68321=>"000010001",
68322=>"000001000",
68323=>"011111011",
68324=>"001001001",
68325=>"000010011",
68326=>"110110100",
68327=>"011000100",
68328=>"111101000",
68329=>"000000000",
68330=>"001100000",
68331=>"001111111",
68332=>"000110110",
68333=>"101001001",
68334=>"000000000",
68335=>"000001011",
68336=>"101001111",
68337=>"100100111",
68338=>"000000010",
68339=>"001110110",
68340=>"110101001",
68341=>"000000000",
68342=>"000010000",
68343=>"110000110",
68344=>"000000101",
68345=>"010011110",
68346=>"111111101",
68347=>"110111111",
68348=>"111100001",
68349=>"001000010",
68350=>"111111000",
68351=>"111110010",
68352=>"011011011",
68353=>"000001000",
68354=>"101000000",
68355=>"001001101",
68356=>"111100100",
68357=>"111000000",
68358=>"000111100",
68359=>"001000011",
68360=>"000111011",
68361=>"001001111",
68362=>"000000001",
68363=>"000110000",
68364=>"000010010",
68365=>"010011100",
68366=>"000100111",
68367=>"000010110",
68368=>"000000000",
68369=>"101000111",
68370=>"111010000",
68371=>"111000000",
68372=>"101101111",
68373=>"111101000",
68374=>"100100000",
68375=>"000101111",
68376=>"000000000",
68377=>"001111110",
68378=>"000001000",
68379=>"111001111",
68380=>"001001111",
68381=>"100001000",
68382=>"110100000",
68383=>"100000110",
68384=>"011001000",
68385=>"001101111",
68386=>"000111000",
68387=>"000000000",
68388=>"100110110",
68389=>"110000110",
68390=>"101000000",
68391=>"000110000",
68392=>"000010010",
68393=>"001001001",
68394=>"000000000",
68395=>"111101111",
68396=>"011111111",
68397=>"000111111",
68398=>"111111100",
68399=>"001101000",
68400=>"110101000",
68401=>"001001010",
68402=>"111111000",
68403=>"101000000",
68404=>"001000000",
68405=>"111110111",
68406=>"110000001",
68407=>"101011110",
68408=>"111101111",
68409=>"101001101",
68410=>"111111000",
68411=>"000001011",
68412=>"100000101",
68413=>"010111010",
68414=>"001000000",
68415=>"000000010",
68416=>"001010110",
68417=>"110000011",
68418=>"000000111",
68419=>"001001001",
68420=>"110010110",
68421=>"001001000",
68422=>"001000000",
68423=>"010010010",
68424=>"010111111",
68425=>"111001000",
68426=>"101000101",
68427=>"111000101",
68428=>"000010010",
68429=>"011111110",
68430=>"000110110",
68431=>"100111110",
68432=>"100000011",
68433=>"010111000",
68434=>"010111000",
68435=>"011011001",
68436=>"000000001",
68437=>"000100100",
68438=>"010011011",
68439=>"101000001",
68440=>"110111110",
68441=>"001001000",
68442=>"100101011",
68443=>"000011010",
68444=>"001000010",
68445=>"100001001",
68446=>"111111011",
68447=>"000000010",
68448=>"010000000",
68449=>"110101101",
68450=>"110000101",
68451=>"001001000",
68452=>"001100111",
68453=>"111000101",
68454=>"011001101",
68455=>"111011000",
68456=>"100110000",
68457=>"000100000",
68458=>"110001101",
68459=>"101111000",
68460=>"111001001",
68461=>"101011001",
68462=>"000000110",
68463=>"001101101",
68464=>"111111111",
68465=>"001000000",
68466=>"001000100",
68467=>"000010000",
68468=>"000100010",
68469=>"101001000",
68470=>"001000110",
68471=>"110110100",
68472=>"110001101",
68473=>"011011111",
68474=>"001111110",
68475=>"000111111",
68476=>"001001000",
68477=>"010100101",
68478=>"011000100",
68479=>"101000001",
68480=>"000110111",
68481=>"111000000",
68482=>"111001001",
68483=>"000110110",
68484=>"100011000",
68485=>"111111111",
68486=>"011100110",
68487=>"000100001",
68488=>"101111110",
68489=>"100000000",
68490=>"101100100",
68491=>"110010000",
68492=>"001001111",
68493=>"000110010",
68494=>"011001000",
68495=>"001000110",
68496=>"100100110",
68497=>"101110110",
68498=>"101000011",
68499=>"111101000",
68500=>"001110000",
68501=>"111000001",
68502=>"101111111",
68503=>"000010000",
68504=>"001000100",
68505=>"101110100",
68506=>"000010000",
68507=>"000000101",
68508=>"101001001",
68509=>"111111011",
68510=>"011001111",
68511=>"010000010",
68512=>"000011111",
68513=>"001000100",
68514=>"111001001",
68515=>"010101001",
68516=>"010111000",
68517=>"000110110",
68518=>"000110000",
68519=>"000000000",
68520=>"110010011",
68521=>"110111101",
68522=>"110111000",
68523=>"101000111",
68524=>"000010010",
68525=>"111001001",
68526=>"011001110",
68527=>"000110010",
68528=>"100000000",
68529=>"100011010",
68530=>"010001110",
68531=>"001000000",
68532=>"100011010",
68533=>"000000101",
68534=>"000011011",
68535=>"011110100",
68536=>"011000001",
68537=>"000111110",
68538=>"111000111",
68539=>"010000001",
68540=>"100110001",
68541=>"000110110",
68542=>"011011011",
68543=>"111110010",
68544=>"101000000",
68545=>"001000000",
68546=>"001101111",
68547=>"000100110",
68548=>"111000000",
68549=>"000011011",
68550=>"000100100",
68551=>"000101111",
68552=>"111101000",
68553=>"000010100",
68554=>"111001000",
68555=>"111010010",
68556=>"111000100",
68557=>"000000000",
68558=>"101000100",
68559=>"010111000",
68560=>"010110000",
68561=>"011011110",
68562=>"101010010",
68563=>"000010111",
68564=>"000011111",
68565=>"001100110",
68566=>"001001101",
68567=>"000001111",
68568=>"110010000",
68569=>"000000000",
68570=>"001111110",
68571=>"101001001",
68572=>"000001001",
68573=>"110110101",
68574=>"111110110",
68575=>"001110100",
68576=>"110000110",
68577=>"101001000",
68578=>"010011110",
68579=>"011101111",
68580=>"111000000",
68581=>"010001011",
68582=>"010111111",
68583=>"111001111",
68584=>"111000000",
68585=>"111110001",
68586=>"101000000",
68587=>"000000000",
68588=>"000001010",
68589=>"010110010",
68590=>"100000000",
68591=>"000111001",
68592=>"010010010",
68593=>"000001110",
68594=>"110111101",
68595=>"000110010",
68596=>"100111110",
68597=>"111000000",
68598=>"000000000",
68599=>"001000000",
68600=>"001000111",
68601=>"100010101",
68602=>"000101110",
68603=>"000111111",
68604=>"110000011",
68605=>"111101000",
68606=>"100110001",
68607=>"111010001",
68608=>"011011010",
68609=>"110110110",
68610=>"110110010",
68611=>"110010010",
68612=>"110111010",
68613=>"100111110",
68614=>"000000111",
68615=>"010110010",
68616=>"100000000",
68617=>"100100110",
68618=>"110011010",
68619=>"111100100",
68620=>"110010010",
68621=>"101000000",
68622=>"000100110",
68623=>"000010110",
68624=>"110110000",
68625=>"111101101",
68626=>"001011001",
68627=>"100100110",
68628=>"101000000",
68629=>"000010100",
68630=>"110100110",
68631=>"001011011",
68632=>"000101111",
68633=>"000110000",
68634=>"111101001",
68635=>"110110110",
68636=>"101111111",
68637=>"100010110",
68638=>"100011110",
68639=>"010000010",
68640=>"111011010",
68641=>"010011011",
68642=>"011101001",
68643=>"000111010",
68644=>"110100110",
68645=>"011001011",
68646=>"110110110",
68647=>"000000100",
68648=>"001111111",
68649=>"001000101",
68650=>"110110110",
68651=>"110010010",
68652=>"011111111",
68653=>"000110110",
68654=>"000000010",
68655=>"111111110",
68656=>"110000000",
68657=>"000000010",
68658=>"001011011",
68659=>"110110110",
68660=>"011011000",
68661=>"110000000",
68662=>"110110011",
68663=>"110110100",
68664=>"010010100",
68665=>"111001011",
68666=>"001101001",
68667=>"110110010",
68668=>"110010100",
68669=>"011011011",
68670=>"100000100",
68671=>"100000000",
68672=>"110110110",
68673=>"111111111",
68674=>"111000000",
68675=>"110110110",
68676=>"111011000",
68677=>"011001000",
68678=>"100000110",
68679=>"001000111",
68680=>"110010100",
68681=>"011101111",
68682=>"100110110",
68683=>"110100010",
68684=>"001001001",
68685=>"001000101",
68686=>"000111111",
68687=>"011010011",
68688=>"110111111",
68689=>"000000000",
68690=>"110010111",
68691=>"110110100",
68692=>"100110010",
68693=>"000100100",
68694=>"100100100",
68695=>"000111111",
68696=>"101101000",
68697=>"001111111",
68698=>"110110011",
68699=>"110110000",
68700=>"110100100",
68701=>"100100100",
68702=>"110110110",
68703=>"100011110",
68704=>"110110110",
68705=>"110110000",
68706=>"110110110",
68707=>"011100110",
68708=>"110110111",
68709=>"001111110",
68710=>"000001000",
68711=>"100000100",
68712=>"000010010",
68713=>"000000100",
68714=>"000111000",
68715=>"100010101",
68716=>"111011010",
68717=>"001001001",
68718=>"111000110",
68719=>"110111110",
68720=>"110100000",
68721=>"110010000",
68722=>"110110110",
68723=>"000000110",
68724=>"011010100",
68725=>"100100100",
68726=>"111110011",
68727=>"110110000",
68728=>"100100000",
68729=>"111001000",
68730=>"000001010",
68731=>"011101111",
68732=>"100110000",
68733=>"001001000",
68734=>"101101001",
68735=>"100100111",
68736=>"110110000",
68737=>"000100110",
68738=>"110110000",
68739=>"110011111",
68740=>"000000010",
68741=>"111010111",
68742=>"000010100",
68743=>"110100100",
68744=>"111111111",
68745=>"110000010",
68746=>"100100110",
68747=>"000001001",
68748=>"001000011",
68749=>"011110011",
68750=>"111100111",
68751=>"100100110",
68752=>"110000000",
68753=>"011111110",
68754=>"000000111",
68755=>"110000000",
68756=>"100110110",
68757=>"010110110",
68758=>"010011010",
68759=>"101000100",
68760=>"010110110",
68761=>"111000001",
68762=>"000010000",
68763=>"100110010",
68764=>"110000000",
68765=>"100111000",
68766=>"001010101",
68767=>"001011111",
68768=>"110110100",
68769=>"110110001",
68770=>"000000000",
68771=>"111111110",
68772=>"100011111",
68773=>"110110010",
68774=>"011001001",
68775=>"000001001",
68776=>"110110110",
68777=>"110100000",
68778=>"011010011",
68779=>"111000110",
68780=>"101001001",
68781=>"000000100",
68782=>"110011010",
68783=>"000000000",
68784=>"000011111",
68785=>"100100010",
68786=>"000001001",
68787=>"110010000",
68788=>"001001111",
68789=>"111110111",
68790=>"000010101",
68791=>"000011111",
68792=>"110110100",
68793=>"011011011",
68794=>"010010000",
68795=>"100110000",
68796=>"101000100",
68797=>"011011011",
68798=>"000000000",
68799=>"100000110",
68800=>"100010000",
68801=>"110110010",
68802=>"000011011",
68803=>"001011111",
68804=>"111101101",
68805=>"100110100",
68806=>"110010110",
68807=>"011011011",
68808=>"000101101",
68809=>"111110010",
68810=>"110010100",
68811=>"100100110",
68812=>"100100100",
68813=>"110000111",
68814=>"100111111",
68815=>"011011011",
68816=>"011111011",
68817=>"100000000",
68818=>"110000100",
68819=>"010010010",
68820=>"000011011",
68821=>"111111000",
68822=>"110010110",
68823=>"011110111",
68824=>"110110100",
68825=>"100100110",
68826=>"011100101",
68827=>"001101101",
68828=>"110110000",
68829=>"001000001",
68830=>"000100100",
68831=>"110110110",
68832=>"000000000",
68833=>"000000010",
68834=>"000011111",
68835=>"110110000",
68836=>"110110110",
68837=>"111111010",
68838=>"110010110",
68839=>"000010111",
68840=>"001000000",
68841=>"111011000",
68842=>"011011011",
68843=>"111111111",
68844=>"100110110",
68845=>"110010010",
68846=>"011011011",
68847=>"000100111",
68848=>"111000100",
68849=>"011001111",
68850=>"100100110",
68851=>"100100100",
68852=>"111101111",
68853=>"110000000",
68854=>"000000110",
68855=>"100100101",
68856=>"100110110",
68857=>"011000000",
68858=>"000000001",
68859=>"000111111",
68860=>"000111111",
68861=>"010011110",
68862=>"000010111",
68863=>"111110111",
68864=>"001000111",
68865=>"110010100",
68866=>"100000111",
68867=>"010110100",
68868=>"000100110",
68869=>"110101011",
68870=>"111111011",
68871=>"111111111",
68872=>"101000010",
68873=>"101000010",
68874=>"010011000",
68875=>"000101101",
68876=>"001101000",
68877=>"101101111",
68878=>"100100110",
68879=>"111100000",
68880=>"111101000",
68881=>"101000000",
68882=>"100000000",
68883=>"100010000",
68884=>"110110001",
68885=>"101000111",
68886=>"111011000",
68887=>"011000000",
68888=>"000100100",
68889=>"101001011",
68890=>"101101111",
68891=>"101101101",
68892=>"101101101",
68893=>"111010111",
68894=>"000111111",
68895=>"101000111",
68896=>"000000000",
68897=>"000000000",
68898=>"011010011",
68899=>"000011000",
68900=>"101001001",
68901=>"001001011",
68902=>"000110111",
68903=>"011011000",
68904=>"011010010",
68905=>"010100111",
68906=>"110000110",
68907=>"010010000",
68908=>"010000010",
68909=>"000111111",
68910=>"000100110",
68911=>"100000001",
68912=>"000000000",
68913=>"001111101",
68914=>"000000000",
68915=>"101101101",
68916=>"010010001",
68917=>"111000101",
68918=>"111110100",
68919=>"100000010",
68920=>"000000001",
68921=>"000000111",
68922=>"101111110",
68923=>"111000000",
68924=>"100001001",
68925=>"111111000",
68926=>"000000000",
68927=>"100110100",
68928=>"000000000",
68929=>"000101100",
68930=>"001000000",
68931=>"011011001",
68932=>"001101010",
68933=>"111000000",
68934=>"000010110",
68935=>"111000011",
68936=>"111001101",
68937=>"111111011",
68938=>"000001011",
68939=>"000101111",
68940=>"000100111",
68941=>"100100000",
68942=>"000001011",
68943=>"110000111",
68944=>"000000010",
68945=>"000100000",
68946=>"111111111",
68947=>"111001000",
68948=>"000000111",
68949=>"110011001",
68950=>"000100101",
68951=>"000000000",
68952=>"001110111",
68953=>"001011110",
68954=>"000000111",
68955=>"001001111",
68956=>"000000110",
68957=>"001111111",
68958=>"101111001",
68959=>"110110110",
68960=>"100101101",
68961=>"010110010",
68962=>"000000111",
68963=>"011011000",
68964=>"000111110",
68965=>"111100011",
68966=>"111111100",
68967=>"101000010",
68968=>"000100111",
68969=>"011101100",
68970=>"101010111",
68971=>"011101111",
68972=>"000110101",
68973=>"000000010",
68974=>"101000011",
68975=>"100010011",
68976=>"000100100",
68977=>"000000000",
68978=>"110111001",
68979=>"000101111",
68980=>"000000000",
68981=>"001001101",
68982=>"101000000",
68983=>"110010100",
68984=>"011000101",
68985=>"111110101",
68986=>"000110001",
68987=>"111000101",
68988=>"010111001",
68989=>"100000000",
68990=>"111111000",
68991=>"010010011",
68992=>"101000000",
68993=>"100100010",
68994=>"001011111",
68995=>"111010010",
68996=>"000111111",
68997=>"011010001",
68998=>"100110100",
68999=>"000000010",
69000=>"001011000",
69001=>"000010010",
69002=>"101111110",
69003=>"010000000",
69004=>"110000000",
69005=>"110000100",
69006=>"101001000",
69007=>"100000000",
69008=>"100000111",
69009=>"111000000",
69010=>"111000000",
69011=>"000111011",
69012=>"111010010",
69013=>"100000000",
69014=>"101110111",
69015=>"101110111",
69016=>"111111000",
69017=>"010000111",
69018=>"101100111",
69019=>"110000000",
69020=>"000000011",
69021=>"101101110",
69022=>"010101101",
69023=>"000011000",
69024=>"011110110",
69025=>"111110000",
69026=>"011010010",
69027=>"101111000",
69028=>"000010110",
69029=>"000100111",
69030=>"110101101",
69031=>"000000111",
69032=>"000100110",
69033=>"000101101",
69034=>"100000001",
69035=>"000000000",
69036=>"000111111",
69037=>"001111010",
69038=>"010011010",
69039=>"111111010",
69040=>"001110000",
69041=>"001001011",
69042=>"100110001",
69043=>"111011011",
69044=>"111100000",
69045=>"111001100",
69046=>"111000110",
69047=>"000100101",
69048=>"101100110",
69049=>"000000100",
69050=>"101110111",
69051=>"101111001",
69052=>"010111111",
69053=>"111000000",
69054=>"001001101",
69055=>"010000000",
69056=>"101101101",
69057=>"101000000",
69058=>"111101100",
69059=>"000000100",
69060=>"000000000",
69061=>"111111011",
69062=>"000111011",
69063=>"000000001",
69064=>"010000110",
69065=>"000100000",
69066=>"111011011",
69067=>"010000101",
69068=>"100100011",
69069=>"000110100",
69070=>"110101000",
69071=>"000000100",
69072=>"000110111",
69073=>"001001011",
69074=>"100111111",
69075=>"011111111",
69076=>"001001010",
69077=>"101101000",
69078=>"000101111",
69079=>"000000000",
69080=>"011111000",
69081=>"101111110",
69082=>"110101111",
69083=>"000000100",
69084=>"111111000",
69085=>"000010111",
69086=>"000001100",
69087=>"001000111",
69088=>"001000000",
69089=>"000100100",
69090=>"111111111",
69091=>"000110110",
69092=>"001000000",
69093=>"111111001",
69094=>"000010110",
69095=>"111110110",
69096=>"100111000",
69097=>"000001100",
69098=>"010110001",
69099=>"101101111",
69100=>"110010000",
69101=>"001110111",
69102=>"000010010",
69103=>"101110111",
69104=>"000100000",
69105=>"011100100",
69106=>"000110010",
69107=>"110110010",
69108=>"100101011",
69109=>"000000111",
69110=>"001000110",
69111=>"010010010",
69112=>"000000000",
69113=>"100100000",
69114=>"111111010",
69115=>"010101000",
69116=>"101100111",
69117=>"011011101",
69118=>"000111110",
69119=>"000000111",
69120=>"110101011",
69121=>"111110000",
69122=>"000000000",
69123=>"111000110",
69124=>"111000000",
69125=>"111100000",
69126=>"111000101",
69127=>"000111111",
69128=>"000101010",
69129=>"010010001",
69130=>"100100000",
69131=>"011000000",
69132=>"000011111",
69133=>"110100010",
69134=>"111111111",
69135=>"111000011",
69136=>"101101101",
69137=>"100000100",
69138=>"000000100",
69139=>"111000000",
69140=>"101000111",
69141=>"000001000",
69142=>"101001001",
69143=>"001110010",
69144=>"000101011",
69145=>"100010010",
69146=>"111111100",
69147=>"111101101",
69148=>"101100010",
69149=>"001000111",
69150=>"011010000",
69151=>"111101000",
69152=>"000111011",
69153=>"000000001",
69154=>"000111111",
69155=>"000010010",
69156=>"000010110",
69157=>"010110000",
69158=>"101111011",
69159=>"001110111",
69160=>"000000111",
69161=>"111101101",
69162=>"111000000",
69163=>"010001010",
69164=>"111011111",
69165=>"111001111",
69166=>"011000000",
69167=>"000011000",
69168=>"000010001",
69169=>"011100110",
69170=>"000111000",
69171=>"010001111",
69172=>"000000001",
69173=>"010000100",
69174=>"010000000",
69175=>"000111000",
69176=>"100010000",
69177=>"100000000",
69178=>"000100000",
69179=>"000000010",
69180=>"000000000",
69181=>"001111010",
69182=>"000000000",
69183=>"111011000",
69184=>"111111111",
69185=>"111110000",
69186=>"010010000",
69187=>"101110100",
69188=>"110000010",
69189=>"101010000",
69190=>"010110100",
69191=>"111110111",
69192=>"011101011",
69193=>"000111011",
69194=>"111101101",
69195=>"111010100",
69196=>"111011010",
69197=>"110110110",
69198=>"011001001",
69199=>"111100111",
69200=>"101000000",
69201=>"111111111",
69202=>"001101111",
69203=>"010001001",
69204=>"010000100",
69205=>"111100100",
69206=>"000111011",
69207=>"111010111",
69208=>"011111001",
69209=>"011010000",
69210=>"101111101",
69211=>"001011011",
69212=>"110010010",
69213=>"110001000",
69214=>"111101101",
69215=>"000101000",
69216=>"111011001",
69217=>"101000000",
69218=>"000000001",
69219=>"100011011",
69220=>"110110010",
69221=>"110111101",
69222=>"010111110",
69223=>"010111010",
69224=>"000010111",
69225=>"001000000",
69226=>"000010101",
69227=>"111111111",
69228=>"001111110",
69229=>"111101101",
69230=>"000011011",
69231=>"111111101",
69232=>"111101001",
69233=>"010000000",
69234=>"111000000",
69235=>"000111110",
69236=>"000000000",
69237=>"101000000",
69238=>"011111111",
69239=>"010000000",
69240=>"101001001",
69241=>"010110111",
69242=>"101000000",
69243=>"000000101",
69244=>"100100100",
69245=>"000100100",
69246=>"011001001",
69247=>"101100111",
69248=>"000010010",
69249=>"011111001",
69250=>"000000010",
69251=>"010000000",
69252=>"110101101",
69253=>"111110000",
69254=>"110011100",
69255=>"000000010",
69256=>"110000110",
69257=>"001000000",
69258=>"111101111",
69259=>"000010111",
69260=>"111101101",
69261=>"000101111",
69262=>"110111111",
69263=>"100000000",
69264=>"100101101",
69265=>"101111110",
69266=>"111111001",
69267=>"110011111",
69268=>"000100011",
69269=>"111100000",
69270=>"011111111",
69271=>"111101100",
69272=>"011111010",
69273=>"011000000",
69274=>"000010010",
69275=>"111000000",
69276=>"000110111",
69277=>"000101101",
69278=>"010010100",
69279=>"000010010",
69280=>"000110001",
69281=>"100000010",
69282=>"010110010",
69283=>"000111111",
69284=>"111100100",
69285=>"000110110",
69286=>"000110110",
69287=>"010010000",
69288=>"101000000",
69289=>"100111000",
69290=>"010100000",
69291=>"101100000",
69292=>"000011010",
69293=>"111000001",
69294=>"110010001",
69295=>"100100000",
69296=>"011000000",
69297=>"001001001",
69298=>"111000011",
69299=>"010100101",
69300=>"010001001",
69301=>"011011010",
69302=>"000011001",
69303=>"010011110",
69304=>"001001000",
69305=>"001101110",
69306=>"111010010",
69307=>"111010011",
69308=>"010111111",
69309=>"111111010",
69310=>"111111110",
69311=>"000000000",
69312=>"101000001",
69313=>"000000111",
69314=>"001010011",
69315=>"011011011",
69316=>"000000011",
69317=>"011100101",
69318=>"111111110",
69319=>"000010010",
69320=>"011001000",
69321=>"111010111",
69322=>"000111111",
69323=>"010000000",
69324=>"111000100",
69325=>"000111100",
69326=>"010010000",
69327=>"111101101",
69328=>"000111111",
69329=>"110011010",
69330=>"001000000",
69331=>"111101111",
69332=>"000010010",
69333=>"110100110",
69334=>"000100000",
69335=>"111101000",
69336=>"010110100",
69337=>"100101000",
69338=>"110001000",
69339=>"011000101",
69340=>"111111001",
69341=>"010101101",
69342=>"000010010",
69343=>"101101000",
69344=>"101000110",
69345=>"010100101",
69346=>"110111111",
69347=>"010000010",
69348=>"110000101",
69349=>"111111100",
69350=>"011100000",
69351=>"111110100",
69352=>"111100111",
69353=>"001000100",
69354=>"101000000",
69355=>"000111110",
69356=>"111101001",
69357=>"010000000",
69358=>"000000001",
69359=>"000000111",
69360=>"011100000",
69361=>"111001110",
69362=>"010110100",
69363=>"110100000",
69364=>"010011011",
69365=>"101101101",
69366=>"001000000",
69367=>"000000100",
69368=>"111111010",
69369=>"101111010",
69370=>"010000000",
69371=>"001101111",
69372=>"100000011",
69373=>"011000000",
69374=>"000001011",
69375=>"000010110",
69376=>"101100010",
69377=>"011111011",
69378=>"100110010",
69379=>"111111000",
69380=>"000000110",
69381=>"111001111",
69382=>"111100111",
69383=>"000111101",
69384=>"000010110",
69385=>"000000111",
69386=>"111001100",
69387=>"000101110",
69388=>"000000000",
69389=>"000010111",
69390=>"000000000",
69391=>"111111010",
69392=>"110000011",
69393=>"111000000",
69394=>"100010111",
69395=>"000111100",
69396=>"111100100",
69397=>"000001111",
69398=>"011110010",
69399=>"011111000",
69400=>"100100101",
69401=>"000011110",
69402=>"010011011",
69403=>"000010011",
69404=>"011100010",
69405=>"000000011",
69406=>"000001000",
69407=>"010110110",
69408=>"111111000",
69409=>"011111000",
69410=>"111110101",
69411=>"111111101",
69412=>"110100110",
69413=>"011011000",
69414=>"000100010",
69415=>"000111010",
69416=>"000100010",
69417=>"011101111",
69418=>"000000101",
69419=>"000010111",
69420=>"000000000",
69421=>"000110111",
69422=>"111111110",
69423=>"111000101",
69424=>"000000010",
69425=>"101111110",
69426=>"111111011",
69427=>"111101100",
69428=>"111101111",
69429=>"111000000",
69430=>"000000011",
69431=>"000100100",
69432=>"000000010",
69433=>"000000100",
69434=>"110000100",
69435=>"011011101",
69436=>"111000000",
69437=>"001111111",
69438=>"110000000",
69439=>"000011011",
69440=>"111111000",
69441=>"101111001",
69442=>"111111011",
69443=>"001100000",
69444=>"011111011",
69445=>"101111100",
69446=>"000111110",
69447=>"111111111",
69448=>"100010000",
69449=>"100101000",
69450=>"010010010",
69451=>"111000000",
69452=>"111111000",
69453=>"011111111",
69454=>"000011001",
69455=>"000000000",
69456=>"000000000",
69457=>"011111110",
69458=>"111101100",
69459=>"110110100",
69460=>"000010111",
69461=>"000000100",
69462=>"000100111",
69463=>"101000001",
69464=>"110111110",
69465=>"111111000",
69466=>"010010001",
69467=>"111111010",
69468=>"000010010",
69469=>"111110010",
69470=>"000000001",
69471=>"100000001",
69472=>"110100000",
69473=>"111011000",
69474=>"000100111",
69475=>"001001000",
69476=>"010011011",
69477=>"011111011",
69478=>"000000000",
69479=>"111011010",
69480=>"111111111",
69481=>"000000111",
69482=>"000000111",
69483=>"001010000",
69484=>"000000000",
69485=>"010111000",
69486=>"000000100",
69487=>"111000000",
69488=>"100111110",
69489=>"110001001",
69490=>"101000110",
69491=>"111011111",
69492=>"100111111",
69493=>"011011001",
69494=>"000001000",
69495=>"000000100",
69496=>"111110111",
69497=>"011011000",
69498=>"111101111",
69499=>"110110100",
69500=>"000001100",
69501=>"010011011",
69502=>"101111111",
69503=>"000010011",
69504=>"101000101",
69505=>"111010001",
69506=>"000111011",
69507=>"111111100",
69508=>"011100000",
69509=>"000000000",
69510=>"110110000",
69511=>"100100000",
69512=>"001111011",
69513=>"110100100",
69514=>"100000000",
69515=>"000111111",
69516=>"000000111",
69517=>"111100000",
69518=>"000000000",
69519=>"011000000",
69520=>"111100111",
69521=>"101000100",
69522=>"000000111",
69523=>"000010000",
69524=>"010101000",
69525=>"111000000",
69526=>"111001000",
69527=>"000000000",
69528=>"000000000",
69529=>"011000011",
69530=>"011111111",
69531=>"111000100",
69532=>"111101111",
69533=>"011111111",
69534=>"000111111",
69535=>"100000000",
69536=>"111111000",
69537=>"111011000",
69538=>"000001111",
69539=>"011111000",
69540=>"100000110",
69541=>"111011011",
69542=>"011010010",
69543=>"000100000",
69544=>"011011101",
69545=>"000111101",
69546=>"011000101",
69547=>"111000100",
69548=>"101101111",
69549=>"111111101",
69550=>"111001000",
69551=>"000000000",
69552=>"101001111",
69553=>"000110000",
69554=>"011011010",
69555=>"111011001",
69556=>"111111110",
69557=>"111000010",
69558=>"100111011",
69559=>"000100111",
69560=>"011000010",
69561=>"001001100",
69562=>"000000001",
69563=>"001111111",
69564=>"110000001",
69565=>"010111111",
69566=>"000111100",
69567=>"000000111",
69568=>"111111000",
69569=>"000000101",
69570=>"010001000",
69571=>"111111011",
69572=>"000000001",
69573=>"011111011",
69574=>"111111100",
69575=>"111000101",
69576=>"111111101",
69577=>"000111111",
69578=>"101111111",
69579=>"000000011",
69580=>"100100110",
69581=>"110110000",
69582=>"111111111",
69583=>"111010100",
69584=>"000111111",
69585=>"100000000",
69586=>"101101101",
69587=>"100101100",
69588=>"001100101",
69589=>"010011011",
69590=>"111100000",
69591=>"110100100",
69592=>"100000111",
69593=>"000111100",
69594=>"111111000",
69595=>"111011000",
69596=>"000000011",
69597=>"100011000",
69598=>"010000000",
69599=>"100111111",
69600=>"000111110",
69601=>"001000000",
69602=>"111000001",
69603=>"000001000",
69604=>"101000000",
69605=>"010000000",
69606=>"111111111",
69607=>"110110000",
69608=>"100111110",
69609=>"000010111",
69610=>"100000001",
69611=>"001000000",
69612=>"111001001",
69613=>"000001111",
69614=>"010000110",
69615=>"011000100",
69616=>"111000101",
69617=>"111110111",
69618=>"000100011",
69619=>"111111011",
69620=>"001011001",
69621=>"000000111",
69622=>"001001000",
69623=>"011000000",
69624=>"110111111",
69625=>"111111111",
69626=>"001000000",
69627=>"111101101",
69628=>"111011000",
69629=>"000000111",
69630=>"000110011",
69631=>"011111010",
69632=>"001001010",
69633=>"111110010",
69634=>"010000011",
69635=>"001110110",
69636=>"100011001",
69637=>"000011111",
69638=>"011110101",
69639=>"010000000",
69640=>"111110000",
69641=>"111111000",
69642=>"100100100",
69643=>"000000111",
69644=>"010000000",
69645=>"000000011",
69646=>"011001010",
69647=>"001000000",
69648=>"111111111",
69649=>"010111001",
69650=>"000000000",
69651=>"111000011",
69652=>"110110100",
69653=>"011000000",
69654=>"011000001",
69655=>"001000011",
69656=>"010010110",
69657=>"111111111",
69658=>"100111111",
69659=>"111111011",
69660=>"111111100",
69661=>"010100000",
69662=>"000111011",
69663=>"101101111",
69664=>"111100001",
69665=>"010110111",
69666=>"111001011",
69667=>"010111010",
69668=>"001001000",
69669=>"100100000",
69670=>"000011110",
69671=>"101111000",
69672=>"110100000",
69673=>"000110100",
69674=>"111001001",
69675=>"100000000",
69676=>"101001111",
69677=>"110111010",
69678=>"001110111",
69679=>"101000000",
69680=>"111111000",
69681=>"101101001",
69682=>"010001000",
69683=>"111011101",
69684=>"101000000",
69685=>"101111011",
69686=>"100100001",
69687=>"000111000",
69688=>"001000101",
69689=>"000100111",
69690=>"100100111",
69691=>"100001001",
69692=>"011101000",
69693=>"101101011",
69694=>"010000000",
69695=>"100000000",
69696=>"011110010",
69697=>"100101010",
69698=>"010111100",
69699=>"000100100",
69700=>"000000111",
69701=>"001000000",
69702=>"110111101",
69703=>"010000111",
69704=>"001000000",
69705=>"111110100",
69706=>"010010010",
69707=>"000000000",
69708=>"000111101",
69709=>"101101111",
69710=>"001101100",
69711=>"111010111",
69712=>"101111111",
69713=>"000000111",
69714=>"001111010",
69715=>"111000000",
69716=>"101111111",
69717=>"000100100",
69718=>"111101100",
69719=>"110011000",
69720=>"111001101",
69721=>"100101001",
69722=>"100111001",
69723=>"100100000",
69724=>"010111101",
69725=>"001100001",
69726=>"010111111",
69727=>"001001001",
69728=>"100010011",
69729=>"010010110",
69730=>"110111001",
69731=>"111111110",
69732=>"100000100",
69733=>"001001101",
69734=>"111111111",
69735=>"111111000",
69736=>"010101001",
69737=>"000111111",
69738=>"111101000",
69739=>"101100101",
69740=>"000101111",
69741=>"011110010",
69742=>"111111011",
69743=>"111101101",
69744=>"100000100",
69745=>"000111111",
69746=>"000001001",
69747=>"000000010",
69748=>"111001100",
69749=>"000000010",
69750=>"000010110",
69751=>"111111000",
69752=>"010101010",
69753=>"110110111",
69754=>"011000000",
69755=>"001000101",
69756=>"000000001",
69757=>"100000000",
69758=>"111000000",
69759=>"000010111",
69760=>"111010000",
69761=>"000111000",
69762=>"111100000",
69763=>"111000101",
69764=>"110111000",
69765=>"101110110",
69766=>"001001000",
69767=>"010000001",
69768=>"001000000",
69769=>"010000110",
69770=>"000011111",
69771=>"000010101",
69772=>"111100010",
69773=>"011001001",
69774=>"111111101",
69775=>"001010000",
69776=>"101100011",
69777=>"010000010",
69778=>"101000000",
69779=>"011010011",
69780=>"011011111",
69781=>"111110111",
69782=>"101101101",
69783=>"000000000",
69784=>"111011101",
69785=>"100111110",
69786=>"011011000",
69787=>"010011110",
69788=>"000011100",
69789=>"110111111",
69790=>"101100110",
69791=>"111000111",
69792=>"100000100",
69793=>"010000000",
69794=>"101001000",
69795=>"111111111",
69796=>"110110111",
69797=>"000000000",
69798=>"000010000",
69799=>"000000010",
69800=>"111111111",
69801=>"010010111",
69802=>"101000000",
69803=>"000010111",
69804=>"000000111",
69805=>"000111101",
69806=>"100100100",
69807=>"110111111",
69808=>"010100001",
69809=>"000011000",
69810=>"000001111",
69811=>"000100100",
69812=>"101100101",
69813=>"011100001",
69814=>"010100000",
69815=>"010011111",
69816=>"100001000",
69817=>"110100100",
69818=>"110011001",
69819=>"111101111",
69820=>"111000010",
69821=>"011111001",
69822=>"001001100",
69823=>"010101000",
69824=>"001101101",
69825=>"000000100",
69826=>"000001110",
69827=>"101000001",
69828=>"111000101",
69829=>"100010001",
69830=>"101001101",
69831=>"010011000",
69832=>"001001111",
69833=>"110111010",
69834=>"000000010",
69835=>"000001101",
69836=>"111101000",
69837=>"100000000",
69838=>"000001000",
69839=>"000101110",
69840=>"110101100",
69841=>"001000000",
69842=>"010111101",
69843=>"100100110",
69844=>"011111101",
69845=>"000111000",
69846=>"000001101",
69847=>"100101111",
69848=>"101000000",
69849=>"010010000",
69850=>"100000000",
69851=>"010000110",
69852=>"001001011",
69853=>"111010000",
69854=>"001111000",
69855=>"100101111",
69856=>"110111100",
69857=>"011011011",
69858=>"010100101",
69859=>"110110111",
69860=>"111001110",
69861=>"111101101",
69862=>"000001011",
69863=>"001011001",
69864=>"010111111",
69865=>"111111010",
69866=>"001001001",
69867=>"111111111",
69868=>"010110011",
69869=>"100110110",
69870=>"000000001",
69871=>"111001001",
69872=>"001000010",
69873=>"110101000",
69874=>"010010111",
69875=>"000001100",
69876=>"100100001",
69877=>"011111111",
69878=>"001111000",
69879=>"001111101",
69880=>"000000000",
69881=>"100111111",
69882=>"111111011",
69883=>"101000111",
69884=>"101101101",
69885=>"010000101",
69886=>"001000000",
69887=>"000010101",
69888=>"011001010",
69889=>"000000000",
69890=>"001000101",
69891=>"110000000",
69892=>"111111111",
69893=>"101101111",
69894=>"110010010",
69895=>"000110000",
69896=>"111110000",
69897=>"101001101",
69898=>"100101100",
69899=>"011011010",
69900=>"000000111",
69901=>"010111010",
69902=>"111011001",
69903=>"000111111",
69904=>"111111011",
69905=>"111001000",
69906=>"000000111",
69907=>"100000000",
69908=>"101101111",
69909=>"001111001",
69910=>"001101101",
69911=>"000111111",
69912=>"101100110",
69913=>"110000000",
69914=>"111110001",
69915=>"000000000",
69916=>"000000110",
69917=>"110110111",
69918=>"111101000",
69919=>"000000000",
69920=>"111100000",
69921=>"001111111",
69922=>"110001000",
69923=>"111000001",
69924=>"011011000",
69925=>"110100000",
69926=>"101101111",
69927=>"110000111",
69928=>"000101000",
69929=>"100110000",
69930=>"000100111",
69931=>"000001111",
69932=>"111111111",
69933=>"111100111",
69934=>"111010000",
69935=>"100100010",
69936=>"101001100",
69937=>"001111010",
69938=>"001111110",
69939=>"101001000",
69940=>"010000111",
69941=>"000001100",
69942=>"000111111",
69943=>"010110110",
69944=>"000101000",
69945=>"000000011",
69946=>"110100000",
69947=>"001000000",
69948=>"100111100",
69949=>"111000010",
69950=>"110000000",
69951=>"001000000",
69952=>"101000110",
69953=>"111001000",
69954=>"111011000",
69955=>"100100000",
69956=>"000000011",
69957=>"010000000",
69958=>"111111001",
69959=>"101011000",
69960=>"011111111",
69961=>"000000000",
69962=>"000000010",
69963=>"010111000",
69964=>"111000000",
69965=>"011011010",
69966=>"100100100",
69967=>"101101111",
69968=>"111000000",
69969=>"000010010",
69970=>"111101000",
69971=>"101001001",
69972=>"000000111",
69973=>"000011111",
69974=>"110110100",
69975=>"001000000",
69976=>"000110100",
69977=>"001000011",
69978=>"100000111",
69979=>"111111111",
69980=>"111001101",
69981=>"011011000",
69982=>"010110111",
69983=>"011001000",
69984=>"111111000",
69985=>"000000000",
69986=>"101000000",
69987=>"100110110",
69988=>"101000000",
69989=>"010111111",
69990=>"000010000",
69991=>"111000110",
69992=>"000111111",
69993=>"101111110",
69994=>"010000111",
69995=>"111000100",
69996=>"000110110",
69997=>"000000100",
69998=>"000010111",
69999=>"100111111",
70000=>"100101000",
70001=>"011111110",
70002=>"011100111",
70003=>"111111000",
70004=>"111111111",
70005=>"001000000",
70006=>"010000101",
70007=>"110000101",
70008=>"100000110",
70009=>"110000000",
70010=>"001001111",
70011=>"000000101",
70012=>"100011001",
70013=>"100100000",
70014=>"000111111",
70015=>"000000001",
70016=>"101000001",
70017=>"101010110",
70018=>"000000111",
70019=>"010000111",
70020=>"111000000",
70021=>"010100101",
70022=>"001100110",
70023=>"110000100",
70024=>"001000000",
70025=>"000001000",
70026=>"101100101",
70027=>"010000000",
70028=>"000110100",
70029=>"111111000",
70030=>"001000101",
70031=>"110000001",
70032=>"110110000",
70033=>"111111111",
70034=>"000110000",
70035=>"101101000",
70036=>"110100000",
70037=>"101001101",
70038=>"111010000",
70039=>"011011011",
70040=>"001101000",
70041=>"000011010",
70042=>"000111010",
70043=>"101100000",
70044=>"101010010",
70045=>"000000000",
70046=>"111110111",
70047=>"101100101",
70048=>"000110111",
70049=>"101001010",
70050=>"000101110",
70051=>"111000011",
70052=>"001011111",
70053=>"110001000",
70054=>"111110110",
70055=>"110110000",
70056=>"110101111",
70057=>"111110000",
70058=>"001000000",
70059=>"111000000",
70060=>"111000000",
70061=>"000000001",
70062=>"100110100",
70063=>"011000000",
70064=>"000110110",
70065=>"001011011",
70066=>"000000000",
70067=>"000000100",
70068=>"110110000",
70069=>"111111101",
70070=>"010000000",
70071=>"011011101",
70072=>"011011000",
70073=>"011001000",
70074=>"111100010",
70075=>"111111100",
70076=>"000010010",
70077=>"111111011",
70078=>"110110000",
70079=>"011111000",
70080=>"100001111",
70081=>"000101111",
70082=>"101111110",
70083=>"001011000",
70084=>"000000111",
70085=>"011000100",
70086=>"010000000",
70087=>"101001000",
70088=>"111000000",
70089=>"000000001",
70090=>"011001101",
70091=>"101001110",
70092=>"100000000",
70093=>"011110100",
70094=>"000011111",
70095=>"001000111",
70096=>"000000111",
70097=>"110110000",
70098=>"111000000",
70099=>"110010111",
70100=>"010000000",
70101=>"100110100",
70102=>"111110100",
70103=>"110000111",
70104=>"000111111",
70105=>"110000010",
70106=>"100000101",
70107=>"000000111",
70108=>"101101111",
70109=>"000110110",
70110=>"111101110",
70111=>"000110111",
70112=>"000000001",
70113=>"101000000",
70114=>"000000111",
70115=>"111111000",
70116=>"100011011",
70117=>"010110000",
70118=>"010110110",
70119=>"011111000",
70120=>"000000111",
70121=>"010011001",
70122=>"001101001",
70123=>"000010001",
70124=>"110110011",
70125=>"110000000",
70126=>"000000000",
70127=>"010100001",
70128=>"000000000",
70129=>"101001111",
70130=>"010011000",
70131=>"110100111",
70132=>"110001010",
70133=>"001000101",
70134=>"010000000",
70135=>"010001110",
70136=>"000110111",
70137=>"111111111",
70138=>"001000111",
70139=>"110011001",
70140=>"111111001",
70141=>"000000111",
70142=>"100100000",
70143=>"111000110",
70144=>"000000000",
70145=>"111111111",
70146=>"010111101",
70147=>"111111111",
70148=>"000100111",
70149=>"110000000",
70150=>"101111110",
70151=>"011111111",
70152=>"011111010",
70153=>"000001000",
70154=>"110000000",
70155=>"000000001",
70156=>"011011000",
70157=>"101101000",
70158=>"000000000",
70159=>"000000100",
70160=>"111111111",
70161=>"000001101",
70162=>"000000110",
70163=>"000000010",
70164=>"000000000",
70165=>"011110100",
70166=>"111111111",
70167=>"111111111",
70168=>"000000111",
70169=>"110101001",
70170=>"000000000",
70171=>"000111111",
70172=>"000110010",
70173=>"111111001",
70174=>"110010011",
70175=>"111111111",
70176=>"000000000",
70177=>"111011101",
70178=>"000001000",
70179=>"001010110",
70180=>"000000111",
70181=>"100101010",
70182=>"011001001",
70183=>"001100010",
70184=>"010000101",
70185=>"000000000",
70186=>"101000100",
70187=>"111111111",
70188=>"110010011",
70189=>"001000110",
70190=>"001011111",
70191=>"110111011",
70192=>"000000000",
70193=>"001011001",
70194=>"000000000",
70195=>"111100000",
70196=>"000000000",
70197=>"010111101",
70198=>"111110100",
70199=>"000000010",
70200=>"000000000",
70201=>"000000000",
70202=>"010000000",
70203=>"100111110",
70204=>"000000001",
70205=>"111111111",
70206=>"010000000",
70207=>"000000010",
70208=>"000000100",
70209=>"000111101",
70210=>"110010000",
70211=>"111111101",
70212=>"000000000",
70213=>"000000000",
70214=>"101000100",
70215=>"101001111",
70216=>"000000000",
70217=>"000001001",
70218=>"000110000",
70219=>"000100111",
70220=>"000000100",
70221=>"000000001",
70222=>"110110010",
70223=>"111111111",
70224=>"010111111",
70225=>"111111111",
70226=>"000000111",
70227=>"001001001",
70228=>"111110000",
70229=>"011000001",
70230=>"100010110",
70231=>"000000000",
70232=>"111001101",
70233=>"001100111",
70234=>"011110010",
70235=>"001011100",
70236=>"000000000",
70237=>"001000100",
70238=>"001111111",
70239=>"111110000",
70240=>"000001011",
70241=>"110000000",
70242=>"000111000",
70243=>"111111111",
70244=>"000010010",
70245=>"000000011",
70246=>"100010000",
70247=>"000000000",
70248=>"010000000",
70249=>"000000000",
70250=>"000011011",
70251=>"000000000",
70252=>"000001000",
70253=>"000000000",
70254=>"110000000",
70255=>"000110101",
70256=>"000110011",
70257=>"000010010",
70258=>"111011011",
70259=>"001000001",
70260=>"000000000",
70261=>"000000000",
70262=>"101000000",
70263=>"000000000",
70264=>"111111111",
70265=>"000100111",
70266=>"000000000",
70267=>"000001010",
70268=>"010000011",
70269=>"100100000",
70270=>"111111110",
70271=>"000000000",
70272=>"101010110",
70273=>"111011011",
70274=>"000110010",
70275=>"111110111",
70276=>"001010111",
70277=>"111111111",
70278=>"000110100",
70279=>"000000000",
70280=>"001000000",
70281=>"000111111",
70282=>"000000000",
70283=>"000000011",
70284=>"111111111",
70285=>"110111101",
70286=>"000000110",
70287=>"000000000",
70288=>"110110110",
70289=>"111001111",
70290=>"000000110",
70291=>"111111001",
70292=>"000000000",
70293=>"001000000",
70294=>"101001001",
70295=>"110000000",
70296=>"010111011",
70297=>"000010101",
70298=>"010111010",
70299=>"011111011",
70300=>"000000000",
70301=>"010010110",
70302=>"000010000",
70303=>"101111011",
70304=>"111000001",
70305=>"111110111",
70306=>"111111000",
70307=>"100111111",
70308=>"010001101",
70309=>"100010010",
70310=>"111010011",
70311=>"110101010",
70312=>"111111111",
70313=>"010001001",
70314=>"111111111",
70315=>"000000100",
70316=>"111101111",
70317=>"000000000",
70318=>"110110100",
70319=>"010001111",
70320=>"111111101",
70321=>"111001001",
70322=>"000100010",
70323=>"000000011",
70324=>"011111000",
70325=>"000010111",
70326=>"001011111",
70327=>"100101111",
70328=>"000000110",
70329=>"011000001",
70330=>"000000010",
70331=>"010000111",
70332=>"100100000",
70333=>"101101111",
70334=>"000011000",
70335=>"111101011",
70336=>"110111110",
70337=>"000000011",
70338=>"000000000",
70339=>"001011001",
70340=>"000000000",
70341=>"001001000",
70342=>"000000100",
70343=>"000000011",
70344=>"111000000",
70345=>"001001110",
70346=>"000000000",
70347=>"010110001",
70348=>"110101011",
70349=>"110110110",
70350=>"111011111",
70351=>"001101111",
70352=>"100111100",
70353=>"111011100",
70354=>"000000000",
70355=>"000000001",
70356=>"111111111",
70357=>"110110111",
70358=>"000010100",
70359=>"000011000",
70360=>"111111110",
70361=>"000001011",
70362=>"011001111",
70363=>"011001001",
70364=>"110110111",
70365=>"111001001",
70366=>"010000001",
70367=>"000000000",
70368=>"010101000",
70369=>"101000011",
70370=>"111110111",
70371=>"000110111",
70372=>"000101000",
70373=>"110000111",
70374=>"001000000",
70375=>"110110111",
70376=>"000000011",
70377=>"001001000",
70378=>"001001001",
70379=>"001000001",
70380=>"000000000",
70381=>"111111111",
70382=>"101110000",
70383=>"010111010",
70384=>"111101100",
70385=>"000000000",
70386=>"101000011",
70387=>"100111010",
70388=>"000001010",
70389=>"111111111",
70390=>"000000000",
70391=>"111111111",
70392=>"010110000",
70393=>"100111111",
70394=>"011111111",
70395=>"010010000",
70396=>"000000000",
70397=>"010110000",
70398=>"000010110",
70399=>"000110111",
70400=>"111001111",
70401=>"000000011",
70402=>"000101111",
70403=>"001010000",
70404=>"111111111",
70405=>"000000101",
70406=>"000100000",
70407=>"011000100",
70408=>"000110111",
70409=>"001111111",
70410=>"111101101",
70411=>"110001000",
70412=>"000000111",
70413=>"000100000",
70414=>"111001011",
70415=>"111000111",
70416=>"011000100",
70417=>"100101101",
70418=>"000000000",
70419=>"000001000",
70420=>"011010001",
70421=>"000000110",
70422=>"001001011",
70423=>"111111000",
70424=>"101000000",
70425=>"111001010",
70426=>"011011011",
70427=>"000111111",
70428=>"000101000",
70429=>"111000001",
70430=>"000000001",
70431=>"111000000",
70432=>"111111010",
70433=>"111011000",
70434=>"011011000",
70435=>"000010110",
70436=>"100000001",
70437=>"110100000",
70438=>"111100000",
70439=>"010111010",
70440=>"111000000",
70441=>"010000110",
70442=>"111101000",
70443=>"000100001",
70444=>"001001001",
70445=>"101000000",
70446=>"110000000",
70447=>"001111011",
70448=>"000000110",
70449=>"011100100",
70450=>"000000111",
70451=>"111100000",
70452=>"111111110",
70453=>"111011111",
70454=>"100111111",
70455=>"101111111",
70456=>"100001101",
70457=>"000101111",
70458=>"000111000",
70459=>"111010010",
70460=>"000000000",
70461=>"111011000",
70462=>"000000000",
70463=>"110011000",
70464=>"000100010",
70465=>"010000101",
70466=>"110000100",
70467=>"000100111",
70468=>"000000000",
70469=>"111000001",
70470=>"000110000",
70471=>"101100111",
70472=>"110100001",
70473=>"000000000",
70474=>"000111111",
70475=>"111000000",
70476=>"000000000",
70477=>"100110110",
70478=>"111111001",
70479=>"111010000",
70480=>"101101111",
70481=>"000011011",
70482=>"001001111",
70483=>"011010000",
70484=>"000000000",
70485=>"010110111",
70486=>"111001000",
70487=>"000000001",
70488=>"000100000",
70489=>"011010000",
70490=>"110100100",
70491=>"111010000",
70492=>"000000000",
70493=>"001000000",
70494=>"100110111",
70495=>"110001111",
70496=>"000111111",
70497=>"000000011",
70498=>"100111111",
70499=>"101001001",
70500=>"010100100",
70501=>"111100001",
70502=>"101000000",
70503=>"111010001",
70504=>"111111000",
70505=>"111010000",
70506=>"010110111",
70507=>"010000111",
70508=>"111110010",
70509=>"111011001",
70510=>"001010000",
70511=>"011000000",
70512=>"100100101",
70513=>"111000000",
70514=>"001110011",
70515=>"101000011",
70516=>"010000000",
70517=>"000000000",
70518=>"000000000",
70519=>"111011111",
70520=>"000111000",
70521=>"111111111",
70522=>"101111111",
70523=>"101111111",
70524=>"110010010",
70525=>"010001000",
70526=>"010010000",
70527=>"100100111",
70528=>"011000000",
70529=>"111000111",
70530=>"000000000",
70531=>"111111111",
70532=>"010101100",
70533=>"011001101",
70534=>"001001100",
70535=>"011010100",
70536=>"001001111",
70537=>"001001101",
70538=>"111110001",
70539=>"010011111",
70540=>"000000000",
70541=>"111111011",
70542=>"000111111",
70543=>"110111111",
70544=>"111100001",
70545=>"101000000",
70546=>"010000000",
70547=>"010101111",
70548=>"011010010",
70549=>"010010101",
70550=>"101101111",
70551=>"011001011",
70552=>"011011000",
70553=>"011010101",
70554=>"000000111",
70555=>"111111000",
70556=>"000000000",
70557=>"000000110",
70558=>"000000101",
70559=>"000001111",
70560=>"001101001",
70561=>"000000000",
70562=>"000000101",
70563=>"100111110",
70564=>"110101011",
70565=>"110001000",
70566=>"111000000",
70567=>"011111000",
70568=>"000011111",
70569=>"010110010",
70570=>"100001101",
70571=>"000100011",
70572=>"111111111",
70573=>"000111010",
70574=>"000000001",
70575=>"011000111",
70576=>"111011111",
70577=>"000001001",
70578=>"111111000",
70579=>"010000001",
70580=>"011000100",
70581=>"000011100",
70582=>"010001010",
70583=>"111000000",
70584=>"000000001",
70585=>"110110000",
70586=>"011000000",
70587=>"000111111",
70588=>"011000000",
70589=>"000000111",
70590=>"001011011",
70591=>"000000000",
70592=>"011000000",
70593=>"111000000",
70594=>"000100100",
70595=>"111110110",
70596=>"000011000",
70597=>"011001011",
70598=>"011011000",
70599=>"101111111",
70600=>"010000000",
70601=>"000001111",
70602=>"000111110",
70603=>"111111111",
70604=>"010000000",
70605=>"011110010",
70606=>"110101001",
70607=>"011000000",
70608=>"011000000",
70609=>"011101111",
70610=>"111010000",
70611=>"011111000",
70612=>"010000000",
70613=>"100100110",
70614=>"001001111",
70615=>"011010000",
70616=>"111000000",
70617=>"111101100",
70618=>"110110100",
70619=>"000111111",
70620=>"000000110",
70621=>"001000111",
70622=>"111100000",
70623=>"111011010",
70624=>"111011000",
70625=>"000100111",
70626=>"111010001",
70627=>"110101111",
70628=>"010000000",
70629=>"001000111",
70630=>"000101111",
70631=>"000011011",
70632=>"000100111",
70633=>"100111111",
70634=>"101001001",
70635=>"000000011",
70636=>"000111111",
70637=>"000000111",
70638=>"000000000",
70639=>"000000000",
70640=>"000000000",
70641=>"111000101",
70642=>"011111111",
70643=>"110100000",
70644=>"000000100",
70645=>"000001001",
70646=>"100001010",
70647=>"111010000",
70648=>"111111001",
70649=>"111001000",
70650=>"001001111",
70651=>"111010001",
70652=>"011111010",
70653=>"111111100",
70654=>"000101111",
70655=>"100000001",
70656=>"000000000",
70657=>"001100000",
70658=>"111011000",
70659=>"011100110",
70660=>"001011011",
70661=>"000000011",
70662=>"111111000",
70663=>"011111111",
70664=>"101101111",
70665=>"000101100",
70666=>"001001111",
70667=>"111000010",
70668=>"111010000",
70669=>"010000001",
70670=>"001011001",
70671=>"001111111",
70672=>"111111111",
70673=>"010000001",
70674=>"000000001",
70675=>"101110000",
70676=>"000111011",
70677=>"000100110",
70678=>"010001000",
70679=>"000001000",
70680=>"111100000",
70681=>"000000000",
70682=>"101111000",
70683=>"111000000",
70684=>"000000100",
70685=>"101111111",
70686=>"001000000",
70687=>"111111010",
70688=>"000100111",
70689=>"111100111",
70690=>"100111111",
70691=>"000111010",
70692=>"001101000",
70693=>"000000001",
70694=>"110000111",
70695=>"110000000",
70696=>"010111101",
70697=>"001111110",
70698=>"100000000",
70699=>"101000001",
70700=>"011001000",
70701=>"111101011",
70702=>"000000001",
70703=>"000000111",
70704=>"000000010",
70705=>"011101111",
70706=>"000011111",
70707=>"000000000",
70708=>"010010000",
70709=>"000010010",
70710=>"110110100",
70711=>"000111111",
70712=>"000000000",
70713=>"000000000",
70714=>"010110111",
70715=>"001101100",
70716=>"110001101",
70717=>"111111111",
70718=>"111000000",
70719=>"100111110",
70720=>"111101000",
70721=>"111011011",
70722=>"100111011",
70723=>"000100110",
70724=>"111100100",
70725=>"010011010",
70726=>"101111110",
70727=>"011000011",
70728=>"111111111",
70729=>"111110000",
70730=>"111011111",
70731=>"101100010",
70732=>"000001001",
70733=>"011001001",
70734=>"100110110",
70735=>"111111011",
70736=>"111000000",
70737=>"000100111",
70738=>"000000000",
70739=>"101100000",
70740=>"011000000",
70741=>"011001111",
70742=>"011101100",
70743=>"011010000",
70744=>"010000000",
70745=>"001000010",
70746=>"110110000",
70747=>"100100100",
70748=>"001000000",
70749=>"001001011",
70750=>"000011000",
70751=>"011001011",
70752=>"000111000",
70753=>"111110000",
70754=>"111010000",
70755=>"011011111",
70756=>"100100000",
70757=>"000001111",
70758=>"110111111",
70759=>"000111111",
70760=>"000000000",
70761=>"010000101",
70762=>"110111111",
70763=>"000101111",
70764=>"101100100",
70765=>"000010111",
70766=>"100111000",
70767=>"000000111",
70768=>"100111011",
70769=>"000000110",
70770=>"001010001",
70771=>"000010000",
70772=>"000101111",
70773=>"000000000",
70774=>"110000000",
70775=>"111111111",
70776=>"011011111",
70777=>"101100000",
70778=>"101000000",
70779=>"000001001",
70780=>"110100001",
70781=>"100001000",
70782=>"000111010",
70783=>"111010000",
70784=>"000000000",
70785=>"000000010",
70786=>"111111111",
70787=>"111101111",
70788=>"101101001",
70789=>"000000000",
70790=>"001001011",
70791=>"111011000",
70792=>"001001110",
70793=>"000100100",
70794=>"000110011",
70795=>"010000000",
70796=>"000000000",
70797=>"000000000",
70798=>"101100100",
70799=>"000010000",
70800=>"100110101",
70801=>"010000000",
70802=>"010111010",
70803=>"011000100",
70804=>"100001000",
70805=>"000001111",
70806=>"110101111",
70807=>"000001011",
70808=>"110000111",
70809=>"010000111",
70810=>"010111111",
70811=>"000001111",
70812=>"000001010",
70813=>"000000111",
70814=>"000100111",
70815=>"111000000",
70816=>"110111101",
70817=>"000000111",
70818=>"111000000",
70819=>"111111111",
70820=>"000000111",
70821=>"011011000",
70822=>"100110110",
70823=>"100101111",
70824=>"001000000",
70825=>"001101111",
70826=>"110110111",
70827=>"111110001",
70828=>"000000000",
70829=>"111111000",
70830=>"000001001",
70831=>"111111001",
70832=>"000000000",
70833=>"001000001",
70834=>"000000111",
70835=>"110110100",
70836=>"110100001",
70837=>"000000000",
70838=>"010010000",
70839=>"000000000",
70840=>"001000101",
70841=>"011001000",
70842=>"011010111",
70843=>"000111111",
70844=>"000010110",
70845=>"000000111",
70846=>"001011011",
70847=>"000010111",
70848=>"101000000",
70849=>"101101001",
70850=>"000111011",
70851=>"101100000",
70852=>"000000101",
70853=>"000001001",
70854=>"001111111",
70855=>"010001111",
70856=>"101111010",
70857=>"111111000",
70858=>"000000000",
70859=>"101111010",
70860=>"000000011",
70861=>"001100100",
70862=>"000000000",
70863=>"001111100",
70864=>"111111010",
70865=>"101100110",
70866=>"111111000",
70867=>"000001000",
70868=>"111011000",
70869=>"000000101",
70870=>"011010111",
70871=>"000111111",
70872=>"000000000",
70873=>"100111111",
70874=>"001101101",
70875=>"011000000",
70876=>"110100001",
70877=>"110111111",
70878=>"010010000",
70879=>"000000001",
70880=>"111111010",
70881=>"000000101",
70882=>"111011000",
70883=>"100100100",
70884=>"100000111",
70885=>"111010110",
70886=>"111111001",
70887=>"101001111",
70888=>"111000111",
70889=>"010001000",
70890=>"100100111",
70891=>"011111111",
70892=>"101110000",
70893=>"000010000",
70894=>"110000000",
70895=>"010000011",
70896=>"010000010",
70897=>"001101100",
70898=>"101100011",
70899=>"100001001",
70900=>"111101000",
70901=>"100000000",
70902=>"010010111",
70903=>"000000101",
70904=>"111010111",
70905=>"000111111",
70906=>"101111111",
70907=>"111100000",
70908=>"000101011",
70909=>"111010000",
70910=>"110100101",
70911=>"000110011",
70912=>"110000000",
70913=>"000000000",
70914=>"111001111",
70915=>"001000011",
70916=>"101111011",
70917=>"110110000",
70918=>"000111111",
70919=>"000010111",
70920=>"101001000",
70921=>"000000111",
70922=>"001100110",
70923=>"110110100",
70924=>"111010000",
70925=>"110110000",
70926=>"110000011",
70927=>"000001101",
70928=>"101111111",
70929=>"000000111",
70930=>"111010010",
70931=>"000000111",
70932=>"001111111",
70933=>"110000111",
70934=>"000110000",
70935=>"000000010",
70936=>"111001001",
70937=>"000101111",
70938=>"000011010",
70939=>"111000110",
70940=>"000000100",
70941=>"001111001",
70942=>"000011111",
70943=>"101001001",
70944=>"111000010",
70945=>"111110000",
70946=>"110110011",
70947=>"110000000",
70948=>"110111001",
70949=>"000000000",
70950=>"101000000",
70951=>"110000001",
70952=>"111001000",
70953=>"110110101",
70954=>"000101101",
70955=>"011111000",
70956=>"000111111",
70957=>"001111010",
70958=>"000110111",
70959=>"000111000",
70960=>"000111111",
70961=>"111011000",
70962=>"111110100",
70963=>"000111111",
70964=>"000101111",
70965=>"100000111",
70966=>"000001011",
70967=>"000000000",
70968=>"000111000",
70969=>"000001111",
70970=>"000000001",
70971=>"000000000",
70972=>"011001000",
70973=>"001000101",
70974=>"100000001",
70975=>"011011001",
70976=>"101110111",
70977=>"110011010",
70978=>"000000000",
70979=>"011100110",
70980=>"110110000",
70981=>"000000001",
70982=>"000001110",
70983=>"101001101",
70984=>"011000010",
70985=>"000111111",
70986=>"000111111",
70987=>"000101001",
70988=>"011000000",
70989=>"110110000",
70990=>"110110100",
70991=>"100110111",
70992=>"101001000",
70993=>"111111010",
70994=>"000111111",
70995=>"101101100",
70996=>"000101111",
70997=>"000110100",
70998=>"011011001",
70999=>"000101111",
71000=>"010101001",
71001=>"011001000",
71002=>"000100000",
71003=>"011100100",
71004=>"000001011",
71005=>"010001001",
71006=>"101111010",
71007=>"100011010",
71008=>"111100000",
71009=>"011110111",
71010=>"111001000",
71011=>"000001011",
71012=>"100100000",
71013=>"000000011",
71014=>"000000111",
71015=>"001111110",
71016=>"110000001",
71017=>"000000111",
71018=>"111110000",
71019=>"000001111",
71020=>"100111100",
71021=>"000001111",
71022=>"000000001",
71023=>"000000000",
71024=>"110110000",
71025=>"010110100",
71026=>"000100110",
71027=>"000010111",
71028=>"111111111",
71029=>"000000101",
71030=>"100000000",
71031=>"110110011",
71032=>"001000111",
71033=>"000000110",
71034=>"111010001",
71035=>"111111000",
71036=>"111110110",
71037=>"000011000",
71038=>"001000000",
71039=>"010000000",
71040=>"100100110",
71041=>"101000000",
71042=>"000010010",
71043=>"101111111",
71044=>"001111111",
71045=>"001000000",
71046=>"000000101",
71047=>"101100011",
71048=>"011000000",
71049=>"010110111",
71050=>"000110111",
71051=>"001001111",
71052=>"110000000",
71053=>"100000001",
71054=>"000110111",
71055=>"000001111",
71056=>"000100001",
71057=>"100101100",
71058=>"010000000",
71059=>"001001111",
71060=>"100111111",
71061=>"001111000",
71062=>"101000101",
71063=>"111111100",
71064=>"101101111",
71065=>"001001100",
71066=>"011000000",
71067=>"001001010",
71068=>"000111110",
71069=>"111100000",
71070=>"000111111",
71071=>"000111100",
71072=>"011011000",
71073=>"000111111",
71074=>"111010000",
71075=>"001111111",
71076=>"000000010",
71077=>"110111111",
71078=>"000001111",
71079=>"101111111",
71080=>"000111111",
71081=>"110110100",
71082=>"111010000",
71083=>"111111000",
71084=>"111011000",
71085=>"110000000",
71086=>"011001001",
71087=>"010001111",
71088=>"111111001",
71089=>"111110110",
71090=>"001111000",
71091=>"111010000",
71092=>"001001101",
71093=>"001111111",
71094=>"111111010",
71095=>"000010100",
71096=>"100000000",
71097=>"101111111",
71098=>"000110111",
71099=>"000111111",
71100=>"000001110",
71101=>"111111101",
71102=>"111100000",
71103=>"000011111",
71104=>"001001111",
71105=>"111101111",
71106=>"011000111",
71107=>"000001000",
71108=>"110000000",
71109=>"111110111",
71110=>"000101011",
71111=>"111000000",
71112=>"110101110",
71113=>"111110000",
71114=>"111110000",
71115=>"110100011",
71116=>"000101101",
71117=>"111100001",
71118=>"100111101",
71119=>"111111011",
71120=>"000011101",
71121=>"110111001",
71122=>"000000100",
71123=>"110000101",
71124=>"111001111",
71125=>"000010000",
71126=>"111111000",
71127=>"001111111",
71128=>"000001111",
71129=>"000000000",
71130=>"110100001",
71131=>"000000111",
71132=>"001111101",
71133=>"001111000",
71134=>"000101101",
71135=>"010100111",
71136=>"000000110",
71137=>"110111111",
71138=>"000000001",
71139=>"111010000",
71140=>"000000010",
71141=>"001111110",
71142=>"111111000",
71143=>"000000001",
71144=>"111000000",
71145=>"000000001",
71146=>"000001011",
71147=>"100000001",
71148=>"110110000",
71149=>"111111100",
71150=>"110000000",
71151=>"110110000",
71152=>"010000001",
71153=>"100111011",
71154=>"000010001",
71155=>"110011011",
71156=>"011000000",
71157=>"000011111",
71158=>"000000111",
71159=>"111111000",
71160=>"111111000",
71161=>"111111000",
71162=>"000110110",
71163=>"000011111",
71164=>"000101111",
71165=>"000110000",
71166=>"011100100",
71167=>"000101111",
71168=>"101000000",
71169=>"010010011",
71170=>"100001000",
71171=>"110111111",
71172=>"000000000",
71173=>"100100101",
71174=>"011011011",
71175=>"001001001",
71176=>"001100110",
71177=>"000100000",
71178=>"001100000",
71179=>"001000001",
71180=>"100110110",
71181=>"110100100",
71182=>"100100000",
71183=>"000111101",
71184=>"111001100",
71185=>"011011001",
71186=>"100011001",
71187=>"011011011",
71188=>"100100000",
71189=>"001001011",
71190=>"011101001",
71191=>"000110111",
71192=>"001100000",
71193=>"111011110",
71194=>"011011011",
71195=>"001000000",
71196=>"011110110",
71197=>"100100110",
71198=>"011010000",
71199=>"110010010",
71200=>"100101100",
71201=>"000011111",
71202=>"100000011",
71203=>"100100011",
71204=>"111111111",
71205=>"011101101",
71206=>"011011011",
71207=>"100111111",
71208=>"010000110",
71209=>"110111101",
71210=>"011111001",
71211=>"111001011",
71212=>"000001100",
71213=>"111101011",
71214=>"001100000",
71215=>"000100010",
71216=>"100001110",
71217=>"000000000",
71218=>"100001101",
71219=>"100000001",
71220=>"000000000",
71221=>"011001001",
71222=>"011011001",
71223=>"001001001",
71224=>"001001111",
71225=>"010100101",
71226=>"100100100",
71227=>"000100010",
71228=>"010100100",
71229=>"100110110",
71230=>"010000100",
71231=>"000111001",
71232=>"001001111",
71233=>"011110100",
71234=>"101111001",
71235=>"010001000",
71236=>"010110110",
71237=>"000000000",
71238=>"001011001",
71239=>"111101010",
71240=>"100101110",
71241=>"010010110",
71242=>"000000000",
71243=>"001000000",
71244=>"011011001",
71245=>"000000000",
71246=>"111111111",
71247=>"100100011",
71248=>"011011010",
71249=>"011100110",
71250=>"000000000",
71251=>"000000010",
71252=>"001000010",
71253=>"111101110",
71254=>"111110110",
71255=>"101001100",
71256=>"111110110",
71257=>"001001000",
71258=>"101001101",
71259=>"100001011",
71260=>"100100100",
71261=>"000000000",
71262=>"111011101",
71263=>"001011011",
71264=>"000011000",
71265=>"010110010",
71266=>"100001100",
71267=>"001111111",
71268=>"110110110",
71269=>"101111111",
71270=>"100000010",
71271=>"100000100",
71272=>"100111011",
71273=>"111100100",
71274=>"011001001",
71275=>"000011111",
71276=>"110100110",
71277=>"100100100",
71278=>"001100111",
71279=>"001100100",
71280=>"000000000",
71281=>"000000101",
71282=>"011001010",
71283=>"111011001",
71284=>"011000011",
71285=>"001000000",
71286=>"001011011",
71287=>"011011001",
71288=>"100011001",
71289=>"110110110",
71290=>"001011001",
71291=>"100100110",
71292=>"111000100",
71293=>"111100100",
71294=>"110001100",
71295=>"000000110",
71296=>"100000100",
71297=>"100110000",
71298=>"001000000",
71299=>"100100100",
71300=>"010000000",
71301=>"000001110",
71302=>"001000000",
71303=>"001001000",
71304=>"111111111",
71305=>"011010110",
71306=>"111110110",
71307=>"001001100",
71308=>"000001100",
71309=>"001001101",
71310=>"010000001",
71311=>"101000100",
71312=>"111110011",
71313=>"010000011",
71314=>"000000000",
71315=>"011010011",
71316=>"011011000",
71317=>"000001000",
71318=>"111111111",
71319=>"001000011",
71320=>"001000000",
71321=>"000010010",
71322=>"011100110",
71323=>"100100010",
71324=>"000001010",
71325=>"011101100",
71326=>"001111011",
71327=>"001001001",
71328=>"100000100",
71329=>"110100111",
71330=>"100011111",
71331=>"111100100",
71332=>"011111100",
71333=>"000000100",
71334=>"000011011",
71335=>"000100010",
71336=>"001001001",
71337=>"010010011",
71338=>"110100100",
71339=>"011010001",
71340=>"000101010",
71341=>"011011000",
71342=>"110100101",
71343=>"000001001",
71344=>"110101110",
71345=>"101100100",
71346=>"100100110",
71347=>"100000100",
71348=>"111100111",
71349=>"000000001",
71350=>"111110100",
71351=>"000011101",
71352=>"100011011",
71353=>"000000000",
71354=>"011000001",
71355=>"101000001",
71356=>"100011100",
71357=>"111011111",
71358=>"000001000",
71359=>"100011011",
71360=>"001000001",
71361=>"011011001",
71362=>"001001011",
71363=>"000111101",
71364=>"000100100",
71365=>"111100111",
71366=>"000110110",
71367=>"111101100",
71368=>"101100100",
71369=>"011011010",
71370=>"100110110",
71371=>"001001001",
71372=>"011001010",
71373=>"011010011",
71374=>"001000100",
71375=>"001110000",
71376=>"011011011",
71377=>"111101111",
71378=>"011011010",
71379=>"001011011",
71380=>"011011011",
71381=>"000100100",
71382=>"000000000",
71383=>"100000000",
71384=>"110111011",
71385=>"110011011",
71386=>"101101111",
71387=>"101100100",
71388=>"111100110",
71389=>"100110010",
71390=>"011000010",
71391=>"111001000",
71392=>"001000010",
71393=>"100001101",
71394=>"001011001",
71395=>"100110111",
71396=>"100000010",
71397=>"000100110",
71398=>"001011011",
71399=>"100000100",
71400=>"000011001",
71401=>"100001011",
71402=>"111000000",
71403=>"100110100",
71404=>"001011010",
71405=>"000001111",
71406=>"000100000",
71407=>"000100110",
71408=>"010110110",
71409=>"000100101",
71410=>"011111000",
71411=>"100110100",
71412=>"111111101",
71413=>"101000001",
71414=>"000001011",
71415=>"011011011",
71416=>"000000111",
71417=>"000111011",
71418=>"110100100",
71419=>"101000010",
71420=>"001001000",
71421=>"110100110",
71422=>"111111101",
71423=>"011111001",
71424=>"111011001",
71425=>"011100000",
71426=>"001110100",
71427=>"010101000",
71428=>"111111110",
71429=>"111111110",
71430=>"000111000",
71431=>"011101000",
71432=>"110000000",
71433=>"000000011",
71434=>"001010011",
71435=>"101111011",
71436=>"100100000",
71437=>"101110011",
71438=>"011001011",
71439=>"111100010",
71440=>"000011101",
71441=>"000000110",
71442=>"111000000",
71443=>"000000011",
71444=>"001100000",
71445=>"011100100",
71446=>"111001100",
71447=>"000100101",
71448=>"001110000",
71449=>"010000111",
71450=>"110010001",
71451=>"011011000",
71452=>"111111111",
71453=>"100000000",
71454=>"001000101",
71455=>"101101011",
71456=>"111000000",
71457=>"000001101",
71458=>"000111000",
71459=>"111101000",
71460=>"100100100",
71461=>"110111111",
71462=>"000000000",
71463=>"000100010",
71464=>"010111111",
71465=>"110111111",
71466=>"000000010",
71467=>"111010010",
71468=>"111101011",
71469=>"000000101",
71470=>"001101011",
71471=>"001001000",
71472=>"000011101",
71473=>"111101111",
71474=>"000000000",
71475=>"000010100",
71476=>"101111010",
71477=>"011000000",
71478=>"110100100",
71479=>"111100000",
71480=>"010111000",
71481=>"010110010",
71482=>"111100000",
71483=>"010110100",
71484=>"100000010",
71485=>"011101101",
71486=>"000000000",
71487=>"111111110",
71488=>"000000000",
71489=>"111111111",
71490=>"100100110",
71491=>"110110001",
71492=>"111111100",
71493=>"111001110",
71494=>"100000000",
71495=>"110100001",
71496=>"000111001",
71497=>"010011000",
71498=>"010000000",
71499=>"001111101",
71500=>"000111111",
71501=>"100111011",
71502=>"110110110",
71503=>"111111001",
71504=>"001001010",
71505=>"001010111",
71506=>"111110010",
71507=>"001001001",
71508=>"111000000",
71509=>"000000010",
71510=>"000101011",
71511=>"011001111",
71512=>"100000001",
71513=>"111101111",
71514=>"111110111",
71515=>"000011111",
71516=>"100010010",
71517=>"001001001",
71518=>"010010111",
71519=>"001011000",
71520=>"110000000",
71521=>"000000000",
71522=>"111111111",
71523=>"100101001",
71524=>"100111111",
71525=>"001011001",
71526=>"110010010",
71527=>"000000000",
71528=>"110000000",
71529=>"010010010",
71530=>"000110011",
71531=>"111111000",
71532=>"000111111",
71533=>"000011100",
71534=>"100001000",
71535=>"111111010",
71536=>"111101001",
71537=>"111111000",
71538=>"001000100",
71539=>"000101111",
71540=>"000101111",
71541=>"101000000",
71542=>"000000000",
71543=>"111110110",
71544=>"011000000",
71545=>"011010111",
71546=>"101000000",
71547=>"010000000",
71548=>"110000000",
71549=>"100100100",
71550=>"010010111",
71551=>"000110000",
71552=>"011111100",
71553=>"010001111",
71554=>"001111111",
71555=>"010111010",
71556=>"000000110",
71557=>"110110000",
71558=>"011111111",
71559=>"000001010",
71560=>"100100100",
71561=>"010110010",
71562=>"010011101",
71563=>"111000100",
71564=>"000000010",
71565=>"001111010",
71566=>"000101101",
71567=>"000001000",
71568=>"100101100",
71569=>"111111111",
71570=>"010011001",
71571=>"111000000",
71572=>"000000000",
71573=>"000000000",
71574=>"111111100",
71575=>"001011010",
71576=>"101111011",
71577=>"000101111",
71578=>"111101101",
71579=>"000100100",
71580=>"110111101",
71581=>"111101101",
71582=>"010011001",
71583=>"111001101",
71584=>"111010101",
71585=>"000100000",
71586=>"010000000",
71587=>"011101000",
71588=>"111110100",
71589=>"000000010",
71590=>"100100001",
71591=>"111111010",
71592=>"000000111",
71593=>"000000000",
71594=>"000100100",
71595=>"111010111",
71596=>"000110011",
71597=>"100000100",
71598=>"110010001",
71599=>"111000011",
71600=>"111111111",
71601=>"001001001",
71602=>"000111111",
71603=>"100100110",
71604=>"000100100",
71605=>"111111010",
71606=>"000000011",
71607=>"111010110",
71608=>"001000000",
71609=>"000000000",
71610=>"111001010",
71611=>"111101111",
71612=>"110101011",
71613=>"111111110",
71614=>"001000000",
71615=>"000110010",
71616=>"001101000",
71617=>"000010111",
71618=>"000000111",
71619=>"011111001",
71620=>"000010000",
71621=>"000001000",
71622=>"010000010",
71623=>"010110000",
71624=>"000101111",
71625=>"001000111",
71626=>"011111011",
71627=>"111001101",
71628=>"000000001",
71629=>"011000000",
71630=>"000000000",
71631=>"101100000",
71632=>"000010010",
71633=>"100111101",
71634=>"100000000",
71635=>"111111110",
71636=>"110101000",
71637=>"100100000",
71638=>"111000000",
71639=>"110110010",
71640=>"101100000",
71641=>"100000000",
71642=>"010110101",
71643=>"000000010",
71644=>"001000000",
71645=>"111101000",
71646=>"000101100",
71647=>"000001000",
71648=>"000000011",
71649=>"000000000",
71650=>"000000000",
71651=>"011101010",
71652=>"010000111",
71653=>"111111101",
71654=>"010011101",
71655=>"110011000",
71656=>"000010110",
71657=>"000000000",
71658=>"110110111",
71659=>"111111110",
71660=>"000000000",
71661=>"111110010",
71662=>"001000100",
71663=>"010010111",
71664=>"100110001",
71665=>"000000000",
71666=>"111110010",
71667=>"000001011",
71668=>"110110110",
71669=>"000111111",
71670=>"000000010",
71671=>"101000111",
71672=>"000000000",
71673=>"000001000",
71674=>"001001111",
71675=>"000000000",
71676=>"110101011",
71677=>"111111101",
71678=>"011111000",
71679=>"000100100",
71680=>"101110111",
71681=>"110011110",
71682=>"100100100",
71683=>"000001111",
71684=>"001111011",
71685=>"100100101",
71686=>"011001000",
71687=>"101011001",
71688=>"000100100",
71689=>"100100100",
71690=>"011011110",
71691=>"000011011",
71692=>"000011011",
71693=>"000011111",
71694=>"101110110",
71695=>"111000011",
71696=>"110000000",
71697=>"101000100",
71698=>"101101011",
71699=>"111111000",
71700=>"111101110",
71701=>"111100010",
71702=>"100101110",
71703=>"111111100",
71704=>"000100100",
71705=>"101111111",
71706=>"010100110",
71707=>"000000100",
71708=>"101100111",
71709=>"000001011",
71710=>"000100101",
71711=>"000000001",
71712=>"111100000",
71713=>"111111010",
71714=>"001101111",
71715=>"000000000",
71716=>"111110101",
71717=>"000011011",
71718=>"001011000",
71719=>"100000000",
71720=>"111110110",
71721=>"010111101",
71722=>"110111111",
71723=>"001000000",
71724=>"111111011",
71725=>"011011111",
71726=>"111011000",
71727=>"000000011",
71728=>"011100100",
71729=>"111001001",
71730=>"101101000",
71731=>"000000000",
71732=>"001111111",
71733=>"111011011",
71734=>"010000000",
71735=>"010111001",
71736=>"111000000",
71737=>"110000100",
71738=>"011101011",
71739=>"100100100",
71740=>"001001000",
71741=>"110010010",
71742=>"100100100",
71743=>"000010000",
71744=>"111000001",
71745=>"000100010",
71746=>"100110111",
71747=>"111100011",
71748=>"100100000",
71749=>"010000000",
71750=>"001011111",
71751=>"111100111",
71752=>"101011001",
71753=>"011100101",
71754=>"111000110",
71755=>"111000000",
71756=>"101100100",
71757=>"101011001",
71758=>"110110111",
71759=>"110011111",
71760=>"000000100",
71761=>"111111111",
71762=>"110010111",
71763=>"000000001",
71764=>"000011001",
71765=>"011000010",
71766=>"100110001",
71767=>"100100000",
71768=>"110010111",
71769=>"000000001",
71770=>"000100001",
71771=>"100000100",
71772=>"111100111",
71773=>"001000001",
71774=>"011011011",
71775=>"110110000",
71776=>"010000001",
71777=>"000001001",
71778=>"100100100",
71779=>"100110111",
71780=>"111000001",
71781=>"000001000",
71782=>"011011011",
71783=>"000001001",
71784=>"000000000",
71785=>"100101011",
71786=>"000111011",
71787=>"110111111",
71788=>"000100000",
71789=>"101011001",
71790=>"111100100",
71791=>"100100000",
71792=>"100000000",
71793=>"100000010",
71794=>"001000100",
71795=>"000011110",
71796=>"000000001",
71797=>"100100101",
71798=>"010010011",
71799=>"000000100",
71800=>"000100110",
71801=>"010100000",
71802=>"100100000",
71803=>"101111001",
71804=>"011101000",
71805=>"000001000",
71806=>"000000000",
71807=>"000000100",
71808=>"011100001",
71809=>"111110110",
71810=>"000000101",
71811=>"100111111",
71812=>"011001000",
71813=>"111100111",
71814=>"110110100",
71815=>"111000000",
71816=>"111111111",
71817=>"111010100",
71818=>"000001000",
71819=>"000100000",
71820=>"011000001",
71821=>"111101111",
71822=>"000100011",
71823=>"111100000",
71824=>"100110101",
71825=>"000101111",
71826=>"011000000",
71827=>"010111000",
71828=>"110101000",
71829=>"100100100",
71830=>"000010111",
71831=>"001101110",
71832=>"100100100",
71833=>"100011000",
71834=>"000000110",
71835=>"100100000",
71836=>"111010011",
71837=>"100100000",
71838=>"000000011",
71839=>"000100111",
71840=>"100011001",
71841=>"000000100",
71842=>"000011000",
71843=>"100101111",
71844=>"000100111",
71845=>"011100111",
71846=>"000001100",
71847=>"001100000",
71848=>"111111110",
71849=>"011010011",
71850=>"000100111",
71851=>"111000100",
71852=>"101111111",
71853=>"100100100",
71854=>"000000110",
71855=>"011011000",
71856=>"000110100",
71857=>"111110000",
71858=>"000100111",
71859=>"100000000",
71860=>"010001101",
71861=>"110111111",
71862=>"000100100",
71863=>"000000000",
71864=>"110100000",
71865=>"001001100",
71866=>"010000000",
71867=>"111111111",
71868=>"110001001",
71869=>"111110100",
71870=>"000100100",
71871=>"000000011",
71872=>"110000000",
71873=>"010100100",
71874=>"010011011",
71875=>"000000001",
71876=>"001000001",
71877=>"001101111",
71878=>"001110111",
71879=>"011100100",
71880=>"111111010",
71881=>"010000000",
71882=>"010011110",
71883=>"110111111",
71884=>"000100000",
71885=>"011010000",
71886=>"100100101",
71887=>"111000011",
71888=>"100111111",
71889=>"000011011",
71890=>"110100000",
71891=>"100110001",
71892=>"100100100",
71893=>"100000000",
71894=>"000000000",
71895=>"000111010",
71896=>"010011011",
71897=>"000001011",
71898=>"111001111",
71899=>"101100100",
71900=>"111111010",
71901=>"100000011",
71902=>"000000011",
71903=>"101101100",
71904=>"000000100",
71905=>"001100100",
71906=>"000011011",
71907=>"011001000",
71908=>"010000000",
71909=>"000010010",
71910=>"111100000",
71911=>"110110111",
71912=>"111100100",
71913=>"111011000",
71914=>"100001000",
71915=>"100100100",
71916=>"000010000",
71917=>"011010001",
71918=>"010000000",
71919=>"000100111",
71920=>"000000000",
71921=>"110110111",
71922=>"100000100",
71923=>"100100011",
71924=>"011000100",
71925=>"100101100",
71926=>"000000101",
71927=>"111000000",
71928=>"000000000",
71929=>"111011011",
71930=>"111110111",
71931=>"101111111",
71932=>"111111111",
71933=>"000111111",
71934=>"111111111",
71935=>"011000000",
71936=>"000000001",
71937=>"000000111",
71938=>"111000000",
71939=>"010001111",
71940=>"110000111",
71941=>"000000000",
71942=>"000010110",
71943=>"001001111",
71944=>"111100101",
71945=>"000010000",
71946=>"001011011",
71947=>"000000000",
71948=>"101000001",
71949=>"000000101",
71950=>"100000110",
71951=>"110100100",
71952=>"101111001",
71953=>"000010000",
71954=>"000100000",
71955=>"000000111",
71956=>"111111100",
71957=>"111000000",
71958=>"010111101",
71959=>"111000111",
71960=>"000000000",
71961=>"001111001",
71962=>"000000100",
71963=>"111111000",
71964=>"000000110",
71965=>"010000111",
71966=>"111111100",
71967=>"101000000",
71968=>"000000111",
71969=>"000101111",
71970=>"101111101",
71971=>"100100111",
71972=>"000000011",
71973=>"011011000",
71974=>"000000000",
71975=>"000101101",
71976=>"100011101",
71977=>"100010001",
71978=>"000010000",
71979=>"010001000",
71980=>"000111111",
71981=>"111111111",
71982=>"000011010",
71983=>"111111010",
71984=>"000000111",
71985=>"111001000",
71986=>"111111000",
71987=>"111111111",
71988=>"001010000",
71989=>"110010111",
71990=>"000111110",
71991=>"101001001",
71992=>"110111110",
71993=>"111001011",
71994=>"011111110",
71995=>"110001100",
71996=>"001001011",
71997=>"111110111",
71998=>"000000000",
71999=>"011100101",
72000=>"111001000",
72001=>"101111000",
72002=>"111111111",
72003=>"011110010",
72004=>"000000000",
72005=>"111110000",
72006=>"110000111",
72007=>"111111000",
72008=>"010110111",
72009=>"110111010",
72010=>"000101101",
72011=>"111100000",
72012=>"101110000",
72013=>"111000100",
72014=>"110000000",
72015=>"111001111",
72016=>"000000000",
72017=>"111110111",
72018=>"000000110",
72019=>"001100110",
72020=>"000000110",
72021=>"001001100",
72022=>"110011100",
72023=>"000000001",
72024=>"001111000",
72025=>"111110011",
72026=>"011000000",
72027=>"000100100",
72028=>"000000000",
72029=>"110000001",
72030=>"111111111",
72031=>"101111110",
72032=>"001101111",
72033=>"111001000",
72034=>"000010011",
72035=>"110000000",
72036=>"111001000",
72037=>"111111001",
72038=>"000111100",
72039=>"111000000",
72040=>"001000110",
72041=>"111111000",
72042=>"101111000",
72043=>"110000111",
72044=>"010010111",
72045=>"001010111",
72046=>"111000000",
72047=>"001111110",
72048=>"111011111",
72049=>"000010000",
72050=>"000111011",
72051=>"000000000",
72052=>"101110010",
72053=>"110000000",
72054=>"101110111",
72055=>"001100001",
72056=>"101111011",
72057=>"101111000",
72058=>"100000011",
72059=>"111100000",
72060=>"001101010",
72061=>"000100000",
72062=>"000000010",
72063=>"110000000",
72064=>"000101111",
72065=>"010011011",
72066=>"000000101",
72067=>"010001101",
72068=>"000000111",
72069=>"111111010",
72070=>"000110010",
72071=>"000100000",
72072=>"010000000",
72073=>"111000000",
72074=>"111000100",
72075=>"101100000",
72076=>"000000000",
72077=>"101000101",
72078=>"010000000",
72079=>"011000000",
72080=>"111111111",
72081=>"111101000",
72082=>"010000000",
72083=>"101100000",
72084=>"000001111",
72085=>"000111101",
72086=>"111010000",
72087=>"000000011",
72088=>"000110111",
72089=>"001000111",
72090=>"111000000",
72091=>"111000010",
72092=>"111100100",
72093=>"111000011",
72094=>"101111111",
72095=>"111000000",
72096=>"001100011",
72097=>"111111000",
72098=>"000101101",
72099=>"001000101",
72100=>"001011000",
72101=>"010111111",
72102=>"000111110",
72103=>"000111111",
72104=>"000000110",
72105=>"000111111",
72106=>"110000000",
72107=>"011010000",
72108=>"111001100",
72109=>"001001000",
72110=>"111000000",
72111=>"001000111",
72112=>"111111001",
72113=>"000000000",
72114=>"000000011",
72115=>"000001100",
72116=>"111100111",
72117=>"111110000",
72118=>"011000101",
72119=>"011101101",
72120=>"000000101",
72121=>"000000111",
72122=>"000000000",
72123=>"000101001",
72124=>"000000000",
72125=>"110111111",
72126=>"110001000",
72127=>"011110000",
72128=>"111000000",
72129=>"111000000",
72130=>"111111111",
72131=>"111101110",
72132=>"111111000",
72133=>"111100000",
72134=>"010110111",
72135=>"111010001",
72136=>"011100001",
72137=>"101000111",
72138=>"000000000",
72139=>"100000001",
72140=>"111100000",
72141=>"000101010",
72142=>"111111101",
72143=>"000111111",
72144=>"100000000",
72145=>"110000001",
72146=>"100100100",
72147=>"110111111",
72148=>"101000001",
72149=>"011100000",
72150=>"001111111",
72151=>"111001111",
72152=>"001101110",
72153=>"000011011",
72154=>"011001110",
72155=>"000000000",
72156=>"010111101",
72157=>"000001100",
72158=>"000000000",
72159=>"001111110",
72160=>"111111001",
72161=>"111000000",
72162=>"111000000",
72163=>"111000010",
72164=>"000001000",
72165=>"000010111",
72166=>"000000111",
72167=>"111000000",
72168=>"111101010",
72169=>"000000110",
72170=>"100110010",
72171=>"010000101",
72172=>"011100101",
72173=>"101100000",
72174=>"010000000",
72175=>"111000000",
72176=>"000000000",
72177=>"111001010",
72178=>"000111110",
72179=>"110111110",
72180=>"001000000",
72181=>"010000000",
72182=>"111000000",
72183=>"111101001",
72184=>"000111101",
72185=>"100000110",
72186=>"111000111",
72187=>"110001101",
72188=>"111010111",
72189=>"000010000",
72190=>"110001001",
72191=>"100100000",
72192=>"010110000",
72193=>"100000011",
72194=>"101000000",
72195=>"000111111",
72196=>"100111111",
72197=>"000000000",
72198=>"100000000",
72199=>"000001111",
72200=>"101000000",
72201=>"000010000",
72202=>"011110110",
72203=>"111111111",
72204=>"100000000",
72205=>"000001000",
72206=>"111101011",
72207=>"000000000",
72208=>"110111000",
72209=>"011111011",
72210=>"111011101",
72211=>"010010110",
72212=>"111111111",
72213=>"100010100",
72214=>"110000000",
72215=>"110010111",
72216=>"000111000",
72217=>"110111111",
72218=>"101111111",
72219=>"000001000",
72220=>"111101001",
72221=>"111001111",
72222=>"111011000",
72223=>"010010000",
72224=>"000000000",
72225=>"000010001",
72226=>"101011000",
72227=>"011001000",
72228=>"000100110",
72229=>"001010010",
72230=>"110111100",
72231=>"000000111",
72232=>"110111111",
72233=>"111111111",
72234=>"001100000",
72235=>"111100000",
72236=>"100011011",
72237=>"111110111",
72238=>"101100101",
72239=>"011101001",
72240=>"111001100",
72241=>"000001001",
72242=>"000101110",
72243=>"111010000",
72244=>"110110111",
72245=>"101100110",
72246=>"011011110",
72247=>"000000000",
72248=>"010000000",
72249=>"000000000",
72250=>"101000101",
72251=>"000111001",
72252=>"010011001",
72253=>"011111110",
72254=>"000000000",
72255=>"100110111",
72256=>"110111100",
72257=>"000011111",
72258=>"101000000",
72259=>"100110111",
72260=>"111000000",
72261=>"101000000",
72262=>"111000101",
72263=>"111111001",
72264=>"110110111",
72265=>"000110110",
72266=>"001000000",
72267=>"011110010",
72268=>"000010010",
72269=>"010011001",
72270=>"000100110",
72271=>"010101000",
72272=>"111111111",
72273=>"010010000",
72274=>"001100101",
72275=>"111001000",
72276=>"110000000",
72277=>"010001111",
72278=>"100011000",
72279=>"000111100",
72280=>"111110110",
72281=>"001001001",
72282=>"001000111",
72283=>"111111111",
72284=>"000000000",
72285=>"000001001",
72286=>"111111010",
72287=>"001011110",
72288=>"100000010",
72289=>"110110011",
72290=>"101000100",
72291=>"110100000",
72292=>"011111101",
72293=>"011001001",
72294=>"110110110",
72295=>"111111100",
72296=>"010010111",
72297=>"000000000",
72298=>"110111100",
72299=>"111101110",
72300=>"101111111",
72301=>"000110011",
72302=>"111101101",
72303=>"111111111",
72304=>"000100100",
72305=>"000000001",
72306=>"110110010",
72307=>"000110010",
72308=>"010010000",
72309=>"000000000",
72310=>"000011010",
72311=>"101000000",
72312=>"100000000",
72313=>"110100010",
72314=>"011010011",
72315=>"011111010",
72316=>"110111011",
72317=>"111100000",
72318=>"010000000",
72319=>"111001001",
72320=>"001000011",
72321=>"111101100",
72322=>"111000010",
72323=>"011100101",
72324=>"111111101",
72325=>"111101010",
72326=>"000010010",
72327=>"000110110",
72328=>"101001011",
72329=>"000010110",
72330=>"010011000",
72331=>"111111010",
72332=>"000110010",
72333=>"111000010",
72334=>"000001011",
72335=>"000000000",
72336=>"100111110",
72337=>"010110101",
72338=>"000111111",
72339=>"110111110",
72340=>"001111100",
72341=>"001000101",
72342=>"111111010",
72343=>"100100011",
72344=>"111111111",
72345=>"110111111",
72346=>"000100111",
72347=>"111101000",
72348=>"110101000",
72349=>"000000000",
72350=>"001111111",
72351=>"110100100",
72352=>"001101101",
72353=>"111000000",
72354=>"001101111",
72355=>"010001111",
72356=>"110111100",
72357=>"100011010",
72358=>"111110110",
72359=>"001001000",
72360=>"001100111",
72361=>"000000111",
72362=>"000000111",
72363=>"111000000",
72364=>"111011010",
72365=>"100000100",
72366=>"111110110",
72367=>"011010100",
72368=>"101000000",
72369=>"010111011",
72370=>"011100111",
72371=>"011100100",
72372=>"100101111",
72373=>"111110001",
72374=>"000010011",
72375=>"000000010",
72376=>"010010111",
72377=>"000111111",
72378=>"010110011",
72379=>"000111110",
72380=>"110011011",
72381=>"111111111",
72382=>"101100100",
72383=>"010000000",
72384=>"111000000",
72385=>"010000010",
72386=>"111111111",
72387=>"100110100",
72388=>"111001000",
72389=>"111110110",
72390=>"100110100",
72391=>"010111010",
72392=>"010001010",
72393=>"100000000",
72394=>"110000111",
72395=>"000100111",
72396=>"010111011",
72397=>"011111110",
72398=>"111111111",
72399=>"000000000",
72400=>"100110000",
72401=>"000110110",
72402=>"000010001",
72403=>"000000010",
72404=>"000000100",
72405=>"010100100",
72406=>"000010000",
72407=>"000010110",
72408=>"110111111",
72409=>"010010000",
72410=>"101100100",
72411=>"010110110",
72412=>"111100101",
72413=>"101001011",
72414=>"010111110",
72415=>"000000000",
72416=>"101001000",
72417=>"111000000",
72418=>"101100100",
72419=>"000100100",
72420=>"000000000",
72421=>"111000101",
72422=>"111000000",
72423=>"100101110",
72424=>"010000000",
72425=>"000000000",
72426=>"110011011",
72427=>"011111111",
72428=>"100000000",
72429=>"000000000",
72430=>"000001111",
72431=>"110100000",
72432=>"110111101",
72433=>"111011001",
72434=>"000001000",
72435=>"111101110",
72436=>"001110100",
72437=>"000001111",
72438=>"100000010",
72439=>"111000111",
72440=>"111111111",
72441=>"111000111",
72442=>"010000001",
72443=>"000011010",
72444=>"000000000",
72445=>"101000000",
72446=>"010111111",
72447=>"100000000",
72448=>"101110010",
72449=>"000111111",
72450=>"010000110",
72451=>"000111111",
72452=>"101011000",
72453=>"000001000",
72454=>"000010000",
72455=>"101111010",
72456=>"100000000",
72457=>"010000110",
72458=>"000001000",
72459=>"111000000",
72460=>"111111000",
72461=>"000111111",
72462=>"011010000",
72463=>"000000100",
72464=>"000001000",
72465=>"000000101",
72466=>"011011000",
72467=>"000000010",
72468=>"101101111",
72469=>"010111111",
72470=>"011111111",
72471=>"111110110",
72472=>"011101001",
72473=>"000000101",
72474=>"000000101",
72475=>"111100000",
72476=>"111000011",
72477=>"001000001",
72478=>"010110001",
72479=>"000011111",
72480=>"111101111",
72481=>"000101001",
72482=>"111101000",
72483=>"101111000",
72484=>"001001011",
72485=>"011001000",
72486=>"011011000",
72487=>"001000000",
72488=>"000011111",
72489=>"111111001",
72490=>"000000111",
72491=>"000000111",
72492=>"111001001",
72493=>"111000010",
72494=>"100000100",
72495=>"000010000",
72496=>"000110111",
72497=>"110000000",
72498=>"101110111",
72499=>"101000011",
72500=>"111000000",
72501=>"100100000",
72502=>"110000011",
72503=>"111100000",
72504=>"111101000",
72505=>"101001000",
72506=>"001101111",
72507=>"111010010",
72508=>"111001000",
72509=>"010111011",
72510=>"000001100",
72511=>"100110011",
72512=>"001000000",
72513=>"100000000",
72514=>"110111000",
72515=>"001000000",
72516=>"100111001",
72517=>"000000100",
72518=>"000000111",
72519=>"000001000",
72520=>"101101000",
72521=>"000001000",
72522=>"000010001",
72523=>"000101111",
72524=>"111000000",
72525=>"000000000",
72526=>"001011000",
72527=>"111101000",
72528=>"010010000",
72529=>"011001010",
72530=>"010000001",
72531=>"000000000",
72532=>"000011010",
72533=>"110000100",
72534=>"000011110",
72535=>"000010011",
72536=>"101111111",
72537=>"010100100",
72538=>"000100111",
72539=>"110110000",
72540=>"000000000",
72541=>"000101111",
72542=>"111110000",
72543=>"010010000",
72544=>"111011000",
72545=>"000110111",
72546=>"000000111",
72547=>"111001001",
72548=>"101111000",
72549=>"110000000",
72550=>"111000000",
72551=>"111111111",
72552=>"100110000",
72553=>"000100000",
72554=>"111111000",
72555=>"000010000",
72556=>"011111111",
72557=>"000101111",
72558=>"111111000",
72559=>"011111110",
72560=>"011011011",
72561=>"001111111",
72562=>"011000010",
72563=>"111110010",
72564=>"111101000",
72565=>"000000000",
72566=>"010111001",
72567=>"111010000",
72568=>"111100101",
72569=>"110010011",
72570=>"100000000",
72571=>"000000000",
72572=>"111011100",
72573=>"000001001",
72574=>"110001111",
72575=>"000001111",
72576=>"000010001",
72577=>"000000000",
72578=>"000000100",
72579=>"000101000",
72580=>"101101000",
72581=>"111111010",
72582=>"110110100",
72583=>"110100100",
72584=>"010000111",
72585=>"000000101",
72586=>"100010111",
72587=>"000110000",
72588=>"000000111",
72589=>"010010101",
72590=>"000110110",
72591=>"000000000",
72592=>"111000000",
72593=>"111000000",
72594=>"101001110",
72595=>"000000110",
72596=>"100100100",
72597=>"000000100",
72598=>"011010000",
72599=>"101111011",
72600=>"010010000",
72601=>"000011111",
72602=>"000010111",
72603=>"111000000",
72604=>"100000111",
72605=>"111111011",
72606=>"100011111",
72607=>"000000000",
72608=>"010111101",
72609=>"101011111",
72610=>"000010011",
72611=>"011001000",
72612=>"000000000",
72613=>"011001000",
72614=>"111010000",
72615=>"000000011",
72616=>"100000100",
72617=>"110011111",
72618=>"011101111",
72619=>"001000000",
72620=>"001101101",
72621=>"000010110",
72622=>"101011111",
72623=>"111111000",
72624=>"100100000",
72625=>"001001111",
72626=>"000000101",
72627=>"010110100",
72628=>"110100000",
72629=>"001101101",
72630=>"000100100",
72631=>"111010111",
72632=>"111000000",
72633=>"101101001",
72634=>"111010010",
72635=>"011000011",
72636=>"111001010",
72637=>"111111111",
72638=>"000001110",
72639=>"010111111",
72640=>"000100101",
72641=>"000000000",
72642=>"111111000",
72643=>"110011111",
72644=>"101101111",
72645=>"000101100",
72646=>"000101111",
72647=>"101100111",
72648=>"001100000",
72649=>"111001000",
72650=>"000010001",
72651=>"010000000",
72652=>"011011000",
72653=>"111111000",
72654=>"000000000",
72655=>"000000111",
72656=>"110111000",
72657=>"011111100",
72658=>"101101100",
72659=>"010000000",
72660=>"111101000",
72661=>"000110111",
72662=>"111011010",
72663=>"000100111",
72664=>"111010000",
72665=>"111101000",
72666=>"010111110",
72667=>"001000111",
72668=>"011011110",
72669=>"000010011",
72670=>"111100011",
72671=>"000001000",
72672=>"000000100",
72673=>"000110111",
72674=>"111101000",
72675=>"100111011",
72676=>"110000010",
72677=>"010010000",
72678=>"011001000",
72679=>"101101111",
72680=>"111111000",
72681=>"011001111",
72682=>"001000100",
72683=>"111101101",
72684=>"001111000",
72685=>"001001000",
72686=>"010010010",
72687=>"011000001",
72688=>"101100011",
72689=>"110111110",
72690=>"011110100",
72691=>"000001100",
72692=>"110101001",
72693=>"000000000",
72694=>"011111000",
72695=>"111110000",
72696=>"000100000",
72697=>"111111011",
72698=>"101111111",
72699=>"111000000",
72700=>"111011000",
72701=>"000110110",
72702=>"001000000",
72703=>"000000000",
72704=>"001000110",
72705=>"001000110",
72706=>"100100111",
72707=>"001000001",
72708=>"110100100",
72709=>"011001000",
72710=>"001001000",
72711=>"001000001",
72712=>"110000100",
72713=>"000100110",
72714=>"110000000",
72715=>"110000100",
72716=>"001001000",
72717=>"001001000",
72718=>"110100100",
72719=>"110100100",
72720=>"111011001",
72721=>"111001001",
72722=>"011100011",
72723=>"010010000",
72724=>"001111100",
72725=>"100000000",
72726=>"100111000",
72727=>"110100010",
72728=>"000100000",
72729=>"100111101",
72730=>"001011000",
72731=>"000000011",
72732=>"000000110",
72733=>"011001011",
72734=>"111101011",
72735=>"000100000",
72736=>"010000111",
72737=>"011011000",
72738=>"000100111",
72739=>"000000011",
72740=>"000000000",
72741=>"001111110",
72742=>"100101111",
72743=>"010011000",
72744=>"001001111",
72745=>"000000100",
72746=>"100100000",
72747=>"000001000",
72748=>"100101101",
72749=>"110101011",
72750=>"011100110",
72751=>"000011000",
72752=>"010011011",
72753=>"111010010",
72754=>"000010011",
72755=>"011111111",
72756=>"100100110",
72757=>"100100101",
72758=>"111011110",
72759=>"010100010",
72760=>"011011000",
72761=>"111000111",
72762=>"110100110",
72763=>"010100110",
72764=>"000001000",
72765=>"111111110",
72766=>"100001111",
72767=>"111100000",
72768=>"100110111",
72769=>"001000000",
72770=>"011011000",
72771=>"110000010",
72772=>"000001011",
72773=>"111000100",
72774=>"001000011",
72775=>"111101111",
72776=>"110110010",
72777=>"111011011",
72778=>"110100111",
72779=>"110100100",
72780=>"110100110",
72781=>"001111111",
72782=>"010011111",
72783=>"100100111",
72784=>"001011011",
72785=>"111110111",
72786=>"111110010",
72787=>"000000000",
72788=>"100111111",
72789=>"111111111",
72790=>"011110011",
72791=>"100100001",
72792=>"111000010",
72793=>"111111111",
72794=>"101111001",
72795=>"010010100",
72796=>"001011000",
72797=>"001000000",
72798=>"000011111",
72799=>"100100110",
72800=>"000100010",
72801=>"010011011",
72802=>"111001100",
72803=>"100000000",
72804=>"000110111",
72805=>"001011011",
72806=>"000000111",
72807=>"110100100",
72808=>"110000001",
72809=>"011011001",
72810=>"011000000",
72811=>"100100110",
72812=>"000101111",
72813=>"111001011",
72814=>"011000000",
72815=>"010000110",
72816=>"101111101",
72817=>"111000000",
72818=>"000100111",
72819=>"100100111",
72820=>"001000000",
72821=>"110100010",
72822=>"001001001",
72823=>"011011011",
72824=>"000000000",
72825=>"011001000",
72826=>"100010100",
72827=>"010011100",
72828=>"111111011",
72829=>"111110000",
72830=>"001011011",
72831=>"000101111",
72832=>"100000110",
72833=>"001000000",
72834=>"011000010",
72835=>"000000010",
72836=>"100000110",
72837=>"110110101",
72838=>"000100100",
72839=>"000011111",
72840=>"000000000",
72841=>"011011111",
72842=>"010010011",
72843=>"011011000",
72844=>"000000011",
72845=>"000000000",
72846=>"100101001",
72847=>"110000001",
72848=>"100111111",
72849=>"100110110",
72850=>"000100010",
72851=>"001000111",
72852=>"100001011",
72853=>"000001000",
72854=>"111110111",
72855=>"001000000",
72856=>"000110111",
72857=>"111001001",
72858=>"100100110",
72859=>"000000110",
72860=>"001011011",
72861=>"100001001",
72862=>"111000000",
72863=>"110100110",
72864=>"001000100",
72865=>"111010000",
72866=>"001011000",
72867=>"110000100",
72868=>"001101101",
72869=>"100110111",
72870=>"111111000",
72871=>"011011001",
72872=>"011111011",
72873=>"011010100",
72874=>"001001000",
72875=>"100000100",
72876=>"010011000",
72877=>"101101111",
72878=>"101100110",
72879=>"001011010",
72880=>"000010101",
72881=>"000111111",
72882=>"010011000",
72883=>"000000000",
72884=>"011000011",
72885=>"100010100",
72886=>"011010111",
72887=>"001011010",
72888=>"111011010",
72889=>"100011001",
72890=>"001001010",
72891=>"111000111",
72892=>"001111001",
72893=>"001011011",
72894=>"000000000",
72895=>"001111001",
72896=>"110000000",
72897=>"000100000",
72898=>"110111011",
72899=>"010011010",
72900=>"000110111",
72901=>"100111111",
72902=>"001000001",
72903=>"100100100",
72904=>"000010001",
72905=>"100100100",
72906=>"110111001",
72907=>"101100111",
72908=>"111110110",
72909=>"010000110",
72910=>"110110011",
72911=>"100011111",
72912=>"000100010",
72913=>"110110110",
72914=>"100000101",
72915=>"101000100",
72916=>"110100111",
72917=>"011010011",
72918=>"101100110",
72919=>"111011000",
72920=>"100100010",
72921=>"000001011",
72922=>"110010100",
72923=>"101001001",
72924=>"110100110",
72925=>"001001100",
72926=>"101100100",
72927=>"111100000",
72928=>"100111111",
72929=>"000011000",
72930=>"000001100",
72931=>"101111011",
72932=>"100100100",
72933=>"000000000",
72934=>"011101011",
72935=>"011110010",
72936=>"001001001",
72937=>"100011010",
72938=>"110100000",
72939=>"001011011",
72940=>"001011011",
72941=>"111100101",
72942=>"000100010",
72943=>"001111110",
72944=>"110100110",
72945=>"010111100",
72946=>"010100000",
72947=>"111111101",
72948=>"111111011",
72949=>"001001000",
72950=>"100000000",
72951=>"011001000",
72952=>"000001001",
72953=>"011011000",
72954=>"110100000",
72955=>"000010110",
72956=>"100100110",
72957=>"001011000",
72958=>"001010011",
72959=>"100110110",
72960=>"000000100",
72961=>"110000000",
72962=>"000001001",
72963=>"111101101",
72964=>"000110110",
72965=>"001111111",
72966=>"000000000",
72967=>"000000111",
72968=>"110111111",
72969=>"000010000",
72970=>"001000110",
72971=>"000000000",
72972=>"110100000",
72973=>"000000010",
72974=>"111010010",
72975=>"111000000",
72976=>"100111111",
72977=>"101010111",
72978=>"000111111",
72979=>"101101000",
72980=>"111000000",
72981=>"111101101",
72982=>"000111111",
72983=>"101011111",
72984=>"110001000",
72985=>"111111111",
72986=>"101101111",
72987=>"001000000",
72988=>"000000011",
72989=>"001101000",
72990=>"111111001",
72991=>"111101100",
72992=>"000010011",
72993=>"111111100",
72994=>"100000110",
72995=>"000111111",
72996=>"110110110",
72997=>"000010000",
72998=>"101000000",
72999=>"100000001",
73000=>"110100110",
73001=>"010110100",
73002=>"101000011",
73003=>"110100010",
73004=>"100100001",
73005=>"111001000",
73006=>"000111111",
73007=>"000011000",
73008=>"000010111",
73009=>"011100100",
73010=>"000000000",
73011=>"000111111",
73012=>"000111011",
73013=>"000111001",
73014=>"000111010",
73015=>"100000000",
73016=>"111111111",
73017=>"111001001",
73018=>"011000000",
73019=>"111000000",
73020=>"100010001",
73021=>"000111011",
73022=>"111000010",
73023=>"000000000",
73024=>"111000000",
73025=>"011110100",
73026=>"110111110",
73027=>"000110011",
73028=>"111000000",
73029=>"111011000",
73030=>"111000000",
73031=>"101111000",
73032=>"111111011",
73033=>"110000000",
73034=>"111000000",
73035=>"001111100",
73036=>"111000000",
73037=>"000000110",
73038=>"110001001",
73039=>"110000000",
73040=>"000101010",
73041=>"101111010",
73042=>"100000001",
73043=>"100110000",
73044=>"111001001",
73045=>"000110100",
73046=>"000001011",
73047=>"000000101",
73048=>"111001001",
73049=>"011110110",
73050=>"010010000",
73051=>"111111110",
73052=>"000111111",
73053=>"010010001",
73054=>"111100000",
73055=>"000011000",
73056=>"000000111",
73057=>"000010000",
73058=>"110000101",
73059=>"011011000",
73060=>"011001100",
73061=>"011000111",
73062=>"101110010",
73063=>"000100111",
73064=>"110000101",
73065=>"111011001",
73066=>"000100111",
73067=>"111101111",
73068=>"000111111",
73069=>"111000010",
73070=>"100000000",
73071=>"000000000",
73072=>"001011011",
73073=>"100111111",
73074=>"000110010",
73075=>"111110010",
73076=>"000001010",
73077=>"110000000",
73078=>"001001000",
73079=>"111100000",
73080=>"111111001",
73081=>"000101001",
73082=>"000000000",
73083=>"000110000",
73084=>"000000110",
73085=>"101001100",
73086=>"111101000",
73087=>"010011000",
73088=>"111110110",
73089=>"001101010",
73090=>"000000101",
73091=>"111111110",
73092=>"000001011",
73093=>"111011110",
73094=>"100011011",
73095=>"101011110",
73096=>"000111110",
73097=>"000010010",
73098=>"111010000",
73099=>"101111000",
73100=>"000000000",
73101=>"111000011",
73102=>"001111111",
73103=>"111011111",
73104=>"100000000",
73105=>"111000000",
73106=>"101000101",
73107=>"101010001",
73108=>"000001111",
73109=>"000000111",
73110=>"111111111",
73111=>"010110100",
73112=>"111000010",
73113=>"010001111",
73114=>"001011010",
73115=>"111111001",
73116=>"110111110",
73117=>"000010110",
73118=>"111111111",
73119=>"000111110",
73120=>"110110001",
73121=>"011110000",
73122=>"100111010",
73123=>"110000001",
73124=>"001000000",
73125=>"111011000",
73126=>"000111110",
73127=>"111101011",
73128=>"000000110",
73129=>"000000111",
73130=>"000111100",
73131=>"000010110",
73132=>"110111110",
73133=>"000000000",
73134=>"001001011",
73135=>"111100000",
73136=>"110000000",
73137=>"110110010",
73138=>"111000000",
73139=>"110000000",
73140=>"001110110",
73141=>"100111110",
73142=>"010111111",
73143=>"101011110",
73144=>"001010011",
73145=>"000110010",
73146=>"000000111",
73147=>"111111001",
73148=>"101111111",
73149=>"011001111",
73150=>"011100110",
73151=>"010111111",
73152=>"111100000",
73153=>"001011011",
73154=>"111000000",
73155=>"000011000",
73156=>"010011010",
73157=>"001000110",
73158=>"000000100",
73159=>"010000111",
73160=>"111000110",
73161=>"111001000",
73162=>"000000000",
73163=>"111000100",
73164=>"010000000",
73165=>"001010011",
73166=>"001111110",
73167=>"000011001",
73168=>"011000000",
73169=>"100001011",
73170=>"001011000",
73171=>"101101101",
73172=>"101011000",
73173=>"001011110",
73174=>"111111101",
73175=>"000000001",
73176=>"110101000",
73177=>"110000101",
73178=>"111111100",
73179=>"111101001",
73180=>"001011011",
73181=>"000100111",
73182=>"111011010",
73183=>"101001100",
73184=>"010000000",
73185=>"000011101",
73186=>"011111001",
73187=>"111111011",
73188=>"001000111",
73189=>"011000101",
73190=>"000000001",
73191=>"000100110",
73192=>"000000000",
73193=>"101110011",
73194=>"110000010",
73195=>"001011111",
73196=>"111101000",
73197=>"101111111",
73198=>"000110000",
73199=>"000000010",
73200=>"111000000",
73201=>"100100110",
73202=>"100000010",
73203=>"110011011",
73204=>"000000101",
73205=>"110000000",
73206=>"100000011",
73207=>"010111111",
73208=>"000000001",
73209=>"111101000",
73210=>"100111100",
73211=>"111101100",
73212=>"111011111",
73213=>"001111111",
73214=>"000011011",
73215=>"010000010",
73216=>"110011000",
73217=>"001101111",
73218=>"000000000",
73219=>"111111111",
73220=>"011101111",
73221=>"111111001",
73222=>"000000000",
73223=>"111010111",
73224=>"111110111",
73225=>"000000000",
73226=>"000000000",
73227=>"111011111",
73228=>"000000110",
73229=>"001000000",
73230=>"111100100",
73231=>"111111100",
73232=>"000001001",
73233=>"111111110",
73234=>"111111110",
73235=>"011100000",
73236=>"101101110",
73237=>"000000000",
73238=>"000010100",
73239=>"001010010",
73240=>"000101000",
73241=>"011111000",
73242=>"111111111",
73243=>"110010010",
73244=>"000000000",
73245=>"000000000",
73246=>"111000000",
73247=>"111000111",
73248=>"000000111",
73249=>"000111111",
73250=>"111011110",
73251=>"111111111",
73252=>"001001011",
73253=>"000010001",
73254=>"111111000",
73255=>"110111110",
73256=>"111011000",
73257=>"111111111",
73258=>"000001000",
73259=>"111111000",
73260=>"000000000",
73261=>"000100010",
73262=>"101011101",
73263=>"001010000",
73264=>"000000010",
73265=>"011011011",
73266=>"001111111",
73267=>"111000000",
73268=>"000000000",
73269=>"000000000",
73270=>"010000000",
73271=>"111010111",
73272=>"111101111",
73273=>"000000000",
73274=>"001101111",
73275=>"000000111",
73276=>"110010011",
73277=>"000011010",
73278=>"001110110",
73279=>"111010011",
73280=>"010000100",
73281=>"000100111",
73282=>"111111111",
73283=>"111101110",
73284=>"111111011",
73285=>"000111111",
73286=>"000000110",
73287=>"110000000",
73288=>"010110101",
73289=>"000000000",
73290=>"000000111",
73291=>"000000000",
73292=>"010110110",
73293=>"110110111",
73294=>"101111101",
73295=>"111001000",
73296=>"011111110",
73297=>"011111000",
73298=>"010111010",
73299=>"011000000",
73300=>"001110000",
73301=>"000110110",
73302=>"010011000",
73303=>"100000000",
73304=>"101110110",
73305=>"100000010",
73306=>"000000001",
73307=>"000000000",
73308=>"011111011",
73309=>"001001111",
73310=>"111111111",
73311=>"011110011",
73312=>"111110111",
73313=>"111111111",
73314=>"000010001",
73315=>"001001000",
73316=>"010001101",
73317=>"000110111",
73318=>"000001001",
73319=>"111011010",
73320=>"111001101",
73321=>"000000000",
73322=>"001011000",
73323=>"010110111",
73324=>"111111111",
73325=>"000001001",
73326=>"111110011",
73327=>"000001111",
73328=>"000000001",
73329=>"000000110",
73330=>"000000000",
73331=>"000000000",
73332=>"111111111",
73333=>"000000000",
73334=>"000001001",
73335=>"111001001",
73336=>"111000000",
73337=>"000001111",
73338=>"001000111",
73339=>"101101111",
73340=>"110000000",
73341=>"110100000",
73342=>"110000001",
73343=>"100100000",
73344=>"111000000",
73345=>"000000001",
73346=>"111111111",
73347=>"111000100",
73348=>"111110000",
73349=>"000010000",
73350=>"000000000",
73351=>"000000111",
73352=>"000000100",
73353=>"010100001",
73354=>"001011000",
73355=>"111000000",
73356=>"111111111",
73357=>"011010010",
73358=>"100111111",
73359=>"011011001",
73360=>"000111011",
73361=>"000000000",
73362=>"000110000",
73363=>"111111010",
73364=>"000001000",
73365=>"111111111",
73366=>"011111111",
73367=>"111111111",
73368=>"001111011",
73369=>"011111111",
73370=>"011010010",
73371=>"100000101",
73372=>"111111110",
73373=>"000000100",
73374=>"111111110",
73375=>"000000000",
73376=>"000101011",
73377=>"000010000",
73378=>"001011010",
73379=>"001011110",
73380=>"111000010",
73381=>"011100001",
73382=>"111110110",
73383=>"000000111",
73384=>"000100011",
73385=>"110111111",
73386=>"110111111",
73387=>"000000000",
73388=>"110010011",
73389=>"111111010",
73390=>"001011010",
73391=>"111111101",
73392=>"100111111",
73393=>"111011011",
73394=>"001110000",
73395=>"100111111",
73396=>"000011111",
73397=>"000000000",
73398=>"111111011",
73399=>"111111100",
73400=>"111110010",
73401=>"100010000",
73402=>"000000000",
73403=>"001001111",
73404=>"000000101",
73405=>"111111011",
73406=>"111111111",
73407=>"000000000",
73408=>"000011010",
73409=>"111111010",
73410=>"000110111",
73411=>"100110111",
73412=>"000010010",
73413=>"110000000",
73414=>"000001000",
73415=>"000000001",
73416=>"010111011",
73417=>"110000000",
73418=>"010111000",
73419=>"000000001",
73420=>"111111100",
73421=>"110000000",
73422=>"000000000",
73423=>"110000101",
73424=>"011010000",
73425=>"101100111",
73426=>"111001000",
73427=>"111111101",
73428=>"110111111",
73429=>"000101111",
73430=>"110111000",
73431=>"001111110",
73432=>"000000000",
73433=>"110000100",
73434=>"000001000",
73435=>"000000000",
73436=>"000011011",
73437=>"111111111",
73438=>"111111000",
73439=>"111000000",
73440=>"111100000",
73441=>"000000000",
73442=>"000111110",
73443=>"111111011",
73444=>"111010000",
73445=>"111010110",
73446=>"101111111",
73447=>"000010000",
73448=>"101001000",
73449=>"110010111",
73450=>"000000000",
73451=>"110000000",
73452=>"111111111",
73453=>"111111111",
73454=>"000000000",
73455=>"101111111",
73456=>"000000000",
73457=>"011001000",
73458=>"111111111",
73459=>"001001000",
73460=>"111110100",
73461=>"000000100",
73462=>"010100110",
73463=>"000000000",
73464=>"000011111",
73465=>"011100111",
73466=>"000000000",
73467=>"001000000",
73468=>"000000101",
73469=>"111111001",
73470=>"111101101",
73471=>"000000000",
73472=>"110010110",
73473=>"110000000",
73474=>"001001111",
73475=>"111000101",
73476=>"011001011",
73477=>"010000001",
73478=>"001000110",
73479=>"101111111",
73480=>"010000001",
73481=>"001001001",
73482=>"000100011",
73483=>"000001000",
73484=>"111000100",
73485=>"000100000",
73486=>"000001001",
73487=>"111000110",
73488=>"000111000",
73489=>"000010110",
73490=>"110000110",
73491=>"011000000",
73492=>"111101001",
73493=>"111000100",
73494=>"100110001",
73495=>"101111110",
73496=>"101000001",
73497=>"011010101",
73498=>"111000000",
73499=>"001001011",
73500=>"101000000",
73501=>"110111000",
73502=>"111101111",
73503=>"111110000",
73504=>"101111010",
73505=>"001100100",
73506=>"100111111",
73507=>"110000000",
73508=>"111001001",
73509=>"100000011",
73510=>"100000000",
73511=>"001100110",
73512=>"000111111",
73513=>"110110110",
73514=>"000000111",
73515=>"000000010",
73516=>"001001001",
73517=>"100101101",
73518=>"110101111",
73519=>"111001110",
73520=>"111000000",
73521=>"111001001",
73522=>"111111110",
73523=>"001011111",
73524=>"011001011",
73525=>"110000111",
73526=>"110001011",
73527=>"111101000",
73528=>"000000111",
73529=>"000000000",
73530=>"100001000",
73531=>"111111111",
73532=>"100111001",
73533=>"110000000",
73534=>"000000000",
73535=>"010000000",
73536=>"001010111",
73537=>"101000001",
73538=>"111011101",
73539=>"100000001",
73540=>"111000000",
73541=>"111111101",
73542=>"001000011",
73543=>"101111101",
73544=>"010011000",
73545=>"000001000",
73546=>"001000000",
73547=>"001101111",
73548=>"001000001",
73549=>"011000101",
73550=>"111100100",
73551=>"111101100",
73552=>"111000000",
73553=>"100111010",
73554=>"010010101",
73555=>"001001000",
73556=>"001000000",
73557=>"110100000",
73558=>"111110000",
73559=>"001010011",
73560=>"111111001",
73561=>"101000000",
73562=>"111001000",
73563=>"000010100",
73564=>"000000000",
73565=>"011001000",
73566=>"010010111",
73567=>"010001000",
73568=>"000000000",
73569=>"001000000",
73570=>"000000111",
73571=>"100110001",
73572=>"111000000",
73573=>"000111000",
73574=>"000000111",
73575=>"010111000",
73576=>"101010111",
73577=>"000010000",
73578=>"000110110",
73579=>"011110000",
73580=>"111111100",
73581=>"001001101",
73582=>"001101110",
73583=>"000000000",
73584=>"011011010",
73585=>"000111111",
73586=>"001100110",
73587=>"000000100",
73588=>"110100000",
73589=>"011000101",
73590=>"000000111",
73591=>"000100101",
73592=>"101001101",
73593=>"010000010",
73594=>"001000000",
73595=>"010000000",
73596=>"000001000",
73597=>"101101011",
73598=>"000110010",
73599=>"101001000",
73600=>"100000111",
73601=>"111010010",
73602=>"001001001",
73603=>"110111000",
73604=>"000001000",
73605=>"000001110",
73606=>"011000000",
73607=>"001001101",
73608=>"010101100",
73609=>"110101101",
73610=>"101101111",
73611=>"110101111",
73612=>"000010111",
73613=>"000100011",
73614=>"000000110",
73615=>"000000101",
73616=>"111101000",
73617=>"101011000",
73618=>"001001111",
73619=>"111111001",
73620=>"000000100",
73621=>"000000111",
73622=>"010011001",
73623=>"001011000",
73624=>"000100101",
73625=>"000010001",
73626=>"000000111",
73627=>"100001111",
73628=>"011011000",
73629=>"101101111",
73630=>"100000000",
73631=>"000000010",
73632=>"011011111",
73633=>"101111111",
73634=>"111111001",
73635=>"101000000",
73636=>"010101111",
73637=>"001001001",
73638=>"011010000",
73639=>"110101000",
73640=>"111000111",
73641=>"110000000",
73642=>"100100111",
73643=>"001000111",
73644=>"110100101",
73645=>"000000001",
73646=>"101111001",
73647=>"000110111",
73648=>"000100111",
73649=>"111011100",
73650=>"111101000",
73651=>"000000000",
73652=>"110010000",
73653=>"011111111",
73654=>"011111111",
73655=>"000000100",
73656=>"011101100",
73657=>"010000000",
73658=>"111000000",
73659=>"011001000",
73660=>"001111000",
73661=>"100110111",
73662=>"000000011",
73663=>"101111110",
73664=>"000000000",
73665=>"000101111",
73666=>"000000010",
73667=>"010000100",
73668=>"001000001",
73669=>"100011110",
73670=>"101111111",
73671=>"000000011",
73672=>"010101111",
73673=>"111001101",
73674=>"010111111",
73675=>"000000101",
73676=>"010000001",
73677=>"000000001",
73678=>"101101110",
73679=>"110111110",
73680=>"000000110",
73681=>"110110100",
73682=>"111001111",
73683=>"011111000",
73684=>"000000001",
73685=>"111100000",
73686=>"111000000",
73687=>"001111000",
73688=>"111110010",
73689=>"010000000",
73690=>"000101111",
73691=>"001000111",
73692=>"111011000",
73693=>"000000111",
73694=>"010111111",
73695=>"111100111",
73696=>"111011101",
73697=>"101110000",
73698=>"101110010",
73699=>"011000001",
73700=>"000011111",
73701=>"000100101",
73702=>"110111111",
73703=>"011111000",
73704=>"000110110",
73705=>"101000000",
73706=>"101001000",
73707=>"000000111",
73708=>"000000001",
73709=>"011000000",
73710=>"000000000",
73711=>"111000000",
73712=>"011000000",
73713=>"011100111",
73714=>"100010010",
73715=>"111101000",
73716=>"110110001",
73717=>"110100101",
73718=>"001101011",
73719=>"000000111",
73720=>"000111111",
73721=>"111110000",
73722=>"110000000",
73723=>"010000001",
73724=>"000000111",
73725=>"000100111",
73726=>"000100100",
73727=>"101001100",
73728=>"101001000",
73729=>"110111001",
73730=>"111011001",
73731=>"101100110",
73732=>"111011011",
73733=>"111000000",
73734=>"000110111",
73735=>"010110010",
73736=>"001000100",
73737=>"110001001",
73738=>"011000100",
73739=>"000010100",
73740=>"111001000",
73741=>"000001100",
73742=>"111001001",
73743=>"100101101",
73744=>"110100001",
73745=>"111000111",
73746=>"110000000",
73747=>"110000000",
73748=>"011110000",
73749=>"111011000",
73750=>"001101111",
73751=>"111001000",
73752=>"111011000",
73753=>"011010011",
73754=>"111001011",
73755=>"100000001",
73756=>"000001001",
73757=>"000101101",
73758=>"001011111",
73759=>"000000111",
73760=>"110111100",
73761=>"001001001",
73762=>"000000101",
73763=>"111001000",
73764=>"000110010",
73765=>"001001001",
73766=>"100011001",
73767=>"000100110",
73768=>"001111110",
73769=>"000111011",
73770=>"110111111",
73771=>"111000000",
73772=>"100001001",
73773=>"100111111",
73774=>"000001100",
73775=>"000100100",
73776=>"001000110",
73777=>"101000111",
73778=>"001010010",
73779=>"001111111",
73780=>"000110100",
73781=>"101111100",
73782=>"111001001",
73783=>"101000001",
73784=>"100110110",
73785=>"111011011",
73786=>"111111100",
73787=>"011011011",
73788=>"111000001",
73789=>"111011001",
73790=>"101001000",
73791=>"010011001",
73792=>"111101001",
73793=>"101011011",
73794=>"001000101",
73795=>"110000011",
73796=>"111011111",
73797=>"011010000",
73798=>"000100010",
73799=>"000110111",
73800=>"100100011",
73801=>"110000000",
73802=>"110010010",
73803=>"111001101",
73804=>"110001001",
73805=>"010101111",
73806=>"111001111",
73807=>"110110110",
73808=>"111000000",
73809=>"100111001",
73810=>"010100100",
73811=>"000110100",
73812=>"001001000",
73813=>"001100100",
73814=>"000010101",
73815=>"011001001",
73816=>"011000111",
73817=>"000000111",
73818=>"111001001",
73819=>"001011110",
73820=>"001001001",
73821=>"100000001",
73822=>"000111111",
73823=>"111100011",
73824=>"111001011",
73825=>"000001000",
73826=>"110001001",
73827=>"111101111",
73828=>"111011110",
73829=>"000110110",
73830=>"010000000",
73831=>"000110100",
73832=>"111001101",
73833=>"110000110",
73834=>"000110000",
73835=>"001011111",
73836=>"001011000",
73837=>"101101100",
73838=>"000000000",
73839=>"111000110",
73840=>"000100101",
73841=>"001000100",
73842=>"110000001",
73843=>"011110100",
73844=>"111100000",
73845=>"010011011",
73846=>"111000011",
73847=>"000100011",
73848=>"000100000",
73849=>"000000011",
73850=>"011011100",
73851=>"000000101",
73852=>"111010001",
73853=>"110101000",
73854=>"000101101",
73855=>"110001001",
73856=>"000000000",
73857=>"110010000",
73858=>"000111111",
73859=>"000100100",
73860=>"000111110",
73861=>"000110100",
73862=>"001001101",
73863=>"111001001",
73864=>"101011111",
73865=>"110010100",
73866=>"001101111",
73867=>"001111001",
73868=>"001000001",
73869=>"110110000",
73870=>"100000000",
73871=>"110000001",
73872=>"010111111",
73873=>"111011010",
73874=>"111001001",
73875=>"111111011",
73876=>"111000001",
73877=>"001001001",
73878=>"111001001",
73879=>"000100100",
73880=>"100110010",
73881=>"000110111",
73882=>"101001111",
73883=>"000100000",
73884=>"110100000",
73885=>"111000010",
73886=>"000111111",
73887=>"010001000",
73888=>"011000000",
73889=>"001111111",
73890=>"000110000",
73891=>"100001110",
73892=>"111110110",
73893=>"000000100",
73894=>"000101100",
73895=>"011001110",
73896=>"001111001",
73897=>"111110000",
73898=>"111001000",
73899=>"110000000",
73900=>"000001000",
73901=>"100001001",
73902=>"111111011",
73903=>"110000110",
73904=>"100110110",
73905=>"100000001",
73906=>"001011111",
73907=>"010000100",
73908=>"001110110",
73909=>"101101101",
73910=>"001111111",
73911=>"100010000",
73912=>"100000001",
73913=>"100101001",
73914=>"000110101",
73915=>"000000011",
73916=>"101000100",
73917=>"110001001",
73918=>"011000011",
73919=>"100110111",
73920=>"110100100",
73921=>"111001000",
73922=>"101000111",
73923=>"000110110",
73924=>"001100100",
73925=>"000110001",
73926=>"001100111",
73927=>"001011011",
73928=>"000000000",
73929=>"010001011",
73930=>"101111110",
73931=>"010000100",
73932=>"100010110",
73933=>"111111001",
73934=>"010001000",
73935=>"111001110",
73936=>"111000001",
73937=>"001010010",
73938=>"011011010",
73939=>"001110111",
73940=>"000000100",
73941=>"111001000",
73942=>"111011001",
73943=>"100110100",
73944=>"000100110",
73945=>"110001000",
73946=>"100100000",
73947=>"100001000",
73948=>"010010001",
73949=>"100110110",
73950=>"000111111",
73951=>"001001111",
73952=>"111110010",
73953=>"101111011",
73954=>"000100110",
73955=>"011100100",
73956=>"111001000",
73957=>"001110011",
73958=>"110111111",
73959=>"100000000",
73960=>"001110110",
73961=>"111001101",
73962=>"111011010",
73963=>"000000001",
73964=>"011110000",
73965=>"001100000",
73966=>"000000000",
73967=>"101110010",
73968=>"010001000",
73969=>"000001011",
73970=>"000011011",
73971=>"000100100",
73972=>"111011111",
73973=>"111001001",
73974=>"011001001",
73975=>"000110110",
73976=>"111001001",
73977=>"100100100",
73978=>"001011001",
73979=>"100001011",
73980=>"000110111",
73981=>"001110110",
73982=>"000010011",
73983=>"010110010",
73984=>"011011000",
73985=>"101101100",
73986=>"100000101",
73987=>"000000100",
73988=>"100111001",
73989=>"110101101",
73990=>"010111111",
73991=>"010000001",
73992=>"000101111",
73993=>"000000101",
73994=>"010110110",
73995=>"010010000",
73996=>"101000110",
73997=>"111011101",
73998=>"100100010",
73999=>"111000000",
74000=>"101101110",
74001=>"000000111",
74002=>"101100110",
74003=>"000001000",
74004=>"111110100",
74005=>"001101111",
74006=>"101000100",
74007=>"001111000",
74008=>"000001101",
74009=>"011001000",
74010=>"011011011",
74011=>"000000101",
74012=>"100101100",
74013=>"111111011",
74014=>"000101101",
74015=>"000100000",
74016=>"000000000",
74017=>"111001110",
74018=>"100111101",
74019=>"000000100",
74020=>"101000001",
74021=>"011001011",
74022=>"000010110",
74023=>"111010000",
74024=>"111111010",
74025=>"011000011",
74026=>"101101000",
74027=>"001000000",
74028=>"000100000",
74029=>"000110111",
74030=>"111111101",
74031=>"101111111",
74032=>"000001111",
74033=>"100101111",
74034=>"011110101",
74035=>"101101111",
74036=>"111010000",
74037=>"100100000",
74038=>"001001001",
74039=>"000010011",
74040=>"111100110",
74041=>"000000000",
74042=>"001111111",
74043=>"000000100",
74044=>"110001000",
74045=>"111111000",
74046=>"000000000",
74047=>"011011101",
74048=>"000110111",
74049=>"001111111",
74050=>"010000111",
74051=>"110111011",
74052=>"111101110",
74053=>"100110111",
74054=>"111100000",
74055=>"000000110",
74056=>"001100000",
74057=>"010011000",
74058=>"000000000",
74059=>"110110011",
74060=>"100100101",
74061=>"100000010",
74062=>"000100111",
74063=>"000000111",
74064=>"000001010",
74065=>"111111111",
74066=>"010010100",
74067=>"101001000",
74068=>"000010100",
74069=>"110000100",
74070=>"111111110",
74071=>"000000001",
74072=>"100111000",
74073=>"000001000",
74074=>"100000001",
74075=>"100001100",
74076=>"111101101",
74077=>"001000000",
74078=>"111000000",
74079=>"011110111",
74080=>"000000111",
74081=>"111111000",
74082=>"000000101",
74083=>"110101000",
74084=>"110000010",
74085=>"101011110",
74086=>"110111000",
74087=>"001100010",
74088=>"111000000",
74089=>"110111101",
74090=>"000011100",
74091=>"110111001",
74092=>"010000111",
74093=>"110111101",
74094=>"110000100",
74095=>"100001010",
74096=>"100110011",
74097=>"000110111",
74098=>"100100000",
74099=>"001000000",
74100=>"011010000",
74101=>"000000000",
74102=>"101010010",
74103=>"010111000",
74104=>"000000000",
74105=>"100111011",
74106=>"100010111",
74107=>"000100001",
74108=>"000011110",
74109=>"000000000",
74110=>"000000101",
74111=>"110110000",
74112=>"111111111",
74113=>"101101111",
74114=>"110000000",
74115=>"100111010",
74116=>"001101001",
74117=>"111010001",
74118=>"100101101",
74119=>"000000000",
74120=>"001010010",
74121=>"110000000",
74122=>"011011010",
74123=>"000000111",
74124=>"111111010",
74125=>"000001011",
74126=>"000101011",
74127=>"000000000",
74128=>"111111011",
74129=>"100111010",
74130=>"010010000",
74131=>"111111111",
74132=>"101110011",
74133=>"001101101",
74134=>"110011010",
74135=>"001111111",
74136=>"010001111",
74137=>"000001000",
74138=>"111110100",
74139=>"101101101",
74140=>"101100111",
74141=>"001000000",
74142=>"101101101",
74143=>"000000000",
74144=>"001000001",
74145=>"001111111",
74146=>"111010011",
74147=>"000100111",
74148=>"101111111",
74149=>"110110011",
74150=>"000100100",
74151=>"000000000",
74152=>"000000101",
74153=>"100100111",
74154=>"101101111",
74155=>"000100010",
74156=>"000111011",
74157=>"000000100",
74158=>"110111000",
74159=>"011101010",
74160=>"101101000",
74161=>"101101001",
74162=>"001111110",
74163=>"000010010",
74164=>"001011011",
74165=>"100111000",
74166=>"000111011",
74167=>"110010111",
74168=>"101100000",
74169=>"111011010",
74170=>"110011100",
74171=>"000011110",
74172=>"110100010",
74173=>"101001000",
74174=>"000000000",
74175=>"000110101",
74176=>"000101000",
74177=>"111111011",
74178=>"001000010",
74179=>"101101101",
74180=>"110010111",
74181=>"101001111",
74182=>"000101011",
74183=>"001000000",
74184=>"110010010",
74185=>"111111111",
74186=>"000111110",
74187=>"000100110",
74188=>"110111000",
74189=>"101110001",
74190=>"101111010",
74191=>"101101101",
74192=>"000000000",
74193=>"111111110",
74194=>"111110110",
74195=>"010010111",
74196=>"101001101",
74197=>"100100110",
74198=>"100000000",
74199=>"110000110",
74200=>"111000000",
74201=>"010011111",
74202=>"010010111",
74203=>"101111101",
74204=>"111001011",
74205=>"000001111",
74206=>"111111111",
74207=>"010011110",
74208=>"000010000",
74209=>"100000100",
74210=>"100111110",
74211=>"001000011",
74212=>"001101001",
74213=>"110110010",
74214=>"100000010",
74215=>"011100010",
74216=>"111110110",
74217=>"000000000",
74218=>"110011001",
74219=>"000000111",
74220=>"010010011",
74221=>"110101100",
74222=>"000000000",
74223=>"011100100",
74224=>"111110000",
74225=>"100000101",
74226=>"000000101",
74227=>"101110010",
74228=>"110001010",
74229=>"001011000",
74230=>"000000000",
74231=>"000100000",
74232=>"000000000",
74233=>"000100100",
74234=>"110010000",
74235=>"101111100",
74236=>"001101111",
74237=>"111000000",
74238=>"101100100",
74239=>"001000000",
74240=>"000001011",
74241=>"100010011",
74242=>"111001000",
74243=>"111000000",
74244=>"011010001",
74245=>"111101000",
74246=>"010101000",
74247=>"000000010",
74248=>"000000000",
74249=>"111000000",
74250=>"111101100",
74251=>"001001111",
74252=>"100000010",
74253=>"000111111",
74254=>"100100100",
74255=>"100000101",
74256=>"011000001",
74257=>"111111000",
74258=>"000000000",
74259=>"100001000",
74260=>"000111111",
74261=>"000010000",
74262=>"000010111",
74263=>"000110110",
74264=>"111001101",
74265=>"100111110",
74266=>"000110111",
74267=>"000000001",
74268=>"000001100",
74269=>"001000000",
74270=>"000000000",
74271=>"001000010",
74272=>"111100101",
74273=>"101000001",
74274=>"000010010",
74275=>"101000000",
74276=>"011110110",
74277=>"010000010",
74278=>"010010010",
74279=>"000100100",
74280=>"110110010",
74281=>"010011111",
74282=>"011001001",
74283=>"000001000",
74284=>"000111011",
74285=>"111111110",
74286=>"110110101",
74287=>"001011001",
74288=>"111000111",
74289=>"000110111",
74290=>"001001000",
74291=>"111000011",
74292=>"111101001",
74293=>"110010010",
74294=>"111110011",
74295=>"000001001",
74296=>"111000000",
74297=>"001001101",
74298=>"000111111",
74299=>"000000110",
74300=>"000011110",
74301=>"010000011",
74302=>"111001000",
74303=>"100101000",
74304=>"111000000",
74305=>"111010001",
74306=>"010111001",
74307=>"000000001",
74308=>"000000111",
74309=>"101001001",
74310=>"000001101",
74311=>"111111110",
74312=>"100000111",
74313=>"110110111",
74314=>"000000000",
74315=>"001000001",
74316=>"110001000",
74317=>"011001111",
74318=>"000000100",
74319=>"000110111",
74320=>"101111100",
74321=>"111010000",
74322=>"100110110",
74323=>"001110011",
74324=>"100000001",
74325=>"111100011",
74326=>"001011011",
74327=>"001001000",
74328=>"000101110",
74329=>"000111111",
74330=>"000111101",
74331=>"000011010",
74332=>"111001001",
74333=>"000110000",
74334=>"111010111",
74335=>"010000101",
74336=>"110111000",
74337=>"000000111",
74338=>"111001001",
74339=>"000011011",
74340=>"001001110",
74341=>"010110110",
74342=>"000010110",
74343=>"111111001",
74344=>"110111100",
74345=>"010111000",
74346=>"001000000",
74347=>"000000111",
74348=>"111111010",
74349=>"111111001",
74350=>"000000001",
74351=>"000000111",
74352=>"000111011",
74353=>"010111110",
74354=>"111111111",
74355=>"111101000",
74356=>"000001010",
74357=>"000000000",
74358=>"011000000",
74359=>"011001000",
74360=>"001111000",
74361=>"000000110",
74362=>"000111101",
74363=>"000001010",
74364=>"011000010",
74365=>"000001110",
74366=>"010001111",
74367=>"001101000",
74368=>"000010010",
74369=>"111110000",
74370=>"111001000",
74371=>"001001110",
74372=>"101000000",
74373=>"001000110",
74374=>"100110100",
74375=>"000000010",
74376=>"001010111",
74377=>"000000111",
74378=>"011111000",
74379=>"000111111",
74380=>"111001001",
74381=>"111101111",
74382=>"001111100",
74383=>"000000000",
74384=>"011111000",
74385=>"010111111",
74386=>"111101101",
74387=>"000110110",
74388=>"001100110",
74389=>"111000000",
74390=>"111100100",
74391=>"000100100",
74392=>"000000000",
74393=>"000000000",
74394=>"110100000",
74395=>"101010010",
74396=>"110001000",
74397=>"111101101",
74398=>"111001000",
74399=>"000000010",
74400=>"000011110",
74401=>"111101001",
74402=>"000000110",
74403=>"101110110",
74404=>"000000100",
74405=>"000111110",
74406=>"001001001",
74407=>"000111101",
74408=>"111111000",
74409=>"010011000",
74410=>"111100001",
74411=>"000001001",
74412=>"001110110",
74413=>"010100101",
74414=>"100110100",
74415=>"011110110",
74416=>"000010110",
74417=>"000101011",
74418=>"000001100",
74419=>"000010011",
74420=>"000110111",
74421=>"101110100",
74422=>"100100111",
74423=>"001111011",
74424=>"000000111",
74425=>"000000110",
74426=>"000001000",
74427=>"100010010",
74428=>"000000001",
74429=>"111111001",
74430=>"011001000",
74431=>"111011001",
74432=>"000010110",
74433=>"010000000",
74434=>"110110111",
74435=>"000100110",
74436=>"000000000",
74437=>"101111011",
74438=>"111110111",
74439=>"000111001",
74440=>"000100101",
74441=>"001000110",
74442=>"001111110",
74443=>"111110000",
74444=>"000001111",
74445=>"100000010",
74446=>"000101101",
74447=>"111111000",
74448=>"011111110",
74449=>"001001111",
74450=>"010000110",
74451=>"001000011",
74452=>"000000111",
74453=>"101101101",
74454=>"101001001",
74455=>"110111001",
74456=>"000110110",
74457=>"010000000",
74458=>"000110110",
74459=>"111101000",
74460=>"000100111",
74461=>"000111001",
74462=>"010000011",
74463=>"000010000",
74464=>"000110110",
74465=>"101100011",
74466=>"001111111",
74467=>"011011011",
74468=>"010111001",
74469=>"110000011",
74470=>"000000101",
74471=>"000011101",
74472=>"101111111",
74473=>"111101001",
74474=>"111001001",
74475=>"111101001",
74476=>"111010110",
74477=>"001111000",
74478=>"000000000",
74479=>"000000110",
74480=>"000001011",
74481=>"101010000",
74482=>"111000000",
74483=>"000110110",
74484=>"111001011",
74485=>"111111001",
74486=>"001001000",
74487=>"010101000",
74488=>"000000110",
74489=>"100110111",
74490=>"000000100",
74491=>"000111111",
74492=>"011010010",
74493=>"000101101",
74494=>"110100001",
74495=>"010110110",
74496=>"011011001",
74497=>"010000111",
74498=>"111101101",
74499=>"000000010",
74500=>"000001001",
74501=>"111111110",
74502=>"100110111",
74503=>"000100111",
74504=>"000000000",
74505=>"001100010",
74506=>"111100000",
74507=>"101000000",
74508=>"000010010",
74509=>"111000100",
74510=>"101001011",
74511=>"000011100",
74512=>"100100010",
74513=>"100001011",
74514=>"111101000",
74515=>"111010000",
74516=>"101101101",
74517=>"111010000",
74518=>"001101111",
74519=>"000000111",
74520=>"111111011",
74521=>"000110110",
74522=>"010111111",
74523=>"000000001",
74524=>"011011000",
74525=>"111000000",
74526=>"001101101",
74527=>"000111000",
74528=>"000010010",
74529=>"010010011",
74530=>"100000000",
74531=>"000000000",
74532=>"011101001",
74533=>"110110111",
74534=>"000000011",
74535=>"000000101",
74536=>"000000111",
74537=>"000001011",
74538=>"000101000",
74539=>"000111111",
74540=>"001000001",
74541=>"101110000",
74542=>"111111111",
74543=>"001101010",
74544=>"110111000",
74545=>"010011011",
74546=>"000111101",
74547=>"111110111",
74548=>"111111001",
74549=>"010000000",
74550=>"100001000",
74551=>"100110010",
74552=>"111010111",
74553=>"111000000",
74554=>"000000000",
74555=>"000100010",
74556=>"000110100",
74557=>"111111000",
74558=>"111101101",
74559=>"110111001",
74560=>"001101101",
74561=>"100010111",
74562=>"111100111",
74563=>"111101000",
74564=>"010010000",
74565=>"100100000",
74566=>"111101110",
74567=>"000001010",
74568=>"010000000",
74569=>"010010000",
74570=>"000000000",
74571=>"010000000",
74572=>"111101100",
74573=>"001111101",
74574=>"000111110",
74575=>"110111000",
74576=>"111000100",
74577=>"111111110",
74578=>"111011000",
74579=>"010011100",
74580=>"101101101",
74581=>"001001110",
74582=>"011011011",
74583=>"111000010",
74584=>"001110011",
74585=>"000011011",
74586=>"011001101",
74587=>"000100100",
74588=>"000110000",
74589=>"010001001",
74590=>"111101111",
74591=>"011100001",
74592=>"000101111",
74593=>"100000010",
74594=>"001000111",
74595=>"100101101",
74596=>"000000000",
74597=>"100100100",
74598=>"000000010",
74599=>"011111100",
74600=>"111011011",
74601=>"111100111",
74602=>"010101101",
74603=>"001010000",
74604=>"000011111",
74605=>"101101111",
74606=>"000110111",
74607=>"101101100",
74608=>"001001000",
74609=>"000000010",
74610=>"000000000",
74611=>"000111110",
74612=>"011010000",
74613=>"101000000",
74614=>"001101101",
74615=>"000100101",
74616=>"111000111",
74617=>"000110111",
74618=>"100000110",
74619=>"100111000",
74620=>"100100110",
74621=>"011110100",
74622=>"011111100",
74623=>"101101001",
74624=>"111000101",
74625=>"111101000",
74626=>"011000000",
74627=>"101111011",
74628=>"011010000",
74629=>"001000010",
74630=>"010011110",
74631=>"000001011",
74632=>"000110100",
74633=>"110110011",
74634=>"100100101",
74635=>"011010000",
74636=>"111101000",
74637=>"111111111",
74638=>"010011000",
74639=>"100000100",
74640=>"011101101",
74641=>"000000000",
74642=>"000000111",
74643=>"111101111",
74644=>"011001111",
74645=>"000100101",
74646=>"111011101",
74647=>"001110111",
74648=>"111001000",
74649=>"010000001",
74650=>"111000000",
74651=>"110000001",
74652=>"010100001",
74653=>"101001000",
74654=>"101111000",
74655=>"000000010",
74656=>"000110111",
74657=>"101001001",
74658=>"000011101",
74659=>"000011111",
74660=>"000111011",
74661=>"000100101",
74662=>"000000000",
74663=>"000000000",
74664=>"011111101",
74665=>"000111111",
74666=>"001011001",
74667=>"111001101",
74668=>"001111111",
74669=>"111000111",
74670=>"110101100",
74671=>"000111111",
74672=>"010111101",
74673=>"000011111",
74674=>"110000111",
74675=>"001000100",
74676=>"100011000",
74677=>"101111101",
74678=>"000011000",
74679=>"000000001",
74680=>"000011011",
74681=>"010011111",
74682=>"000000001",
74683=>"010010010",
74684=>"100010000",
74685=>"010111110",
74686=>"100111110",
74687=>"000011000",
74688=>"111000000",
74689=>"000101111",
74690=>"010010000",
74691=>"110000000",
74692=>"000011101",
74693=>"010011101",
74694=>"000000110",
74695=>"101111111",
74696=>"000010010",
74697=>"001000000",
74698=>"111111110",
74699=>"111000000",
74700=>"001100101",
74701=>"001001110",
74702=>"101101101",
74703=>"000010010",
74704=>"111100000",
74705=>"101111111",
74706=>"000010111",
74707=>"011010000",
74708=>"011101011",
74709=>"000100111",
74710=>"000000000",
74711=>"000111111",
74712=>"111000101",
74713=>"111110010",
74714=>"000000111",
74715=>"111100110",
74716=>"100101000",
74717=>"010000011",
74718=>"101101010",
74719=>"001101111",
74720=>"110000010",
74721=>"111111000",
74722=>"111000000",
74723=>"010011001",
74724=>"000001001",
74725=>"100011010",
74726=>"110110110",
74727=>"001111011",
74728=>"111000101",
74729=>"000010000",
74730=>"111001001",
74731=>"000010010",
74732=>"000000000",
74733=>"110000000",
74734=>"110010110",
74735=>"001000000",
74736=>"000010000",
74737=>"000100001",
74738=>"000111011",
74739=>"000110001",
74740=>"010110111",
74741=>"011111111",
74742=>"000010000",
74743=>"000000101",
74744=>"000111000",
74745=>"110010001",
74746=>"011101100",
74747=>"100101010",
74748=>"011101101",
74749=>"100100000",
74750=>"111100100",
74751=>"110100111",
74752=>"001000100",
74753=>"100101100",
74754=>"000000111",
74755=>"000101111",
74756=>"011110110",
74757=>"000001111",
74758=>"011111101",
74759=>"101010111",
74760=>"000101010",
74761=>"000101010",
74762=>"110100100",
74763=>"000011011",
74764=>"010001001",
74765=>"000000101",
74766=>"100001011",
74767=>"011111100",
74768=>"000000011",
74769=>"000101101",
74770=>"000000001",
74771=>"100000100",
74772=>"011101111",
74773=>"110001010",
74774=>"101101111",
74775=>"010110111",
74776=>"010000100",
74777=>"111101001",
74778=>"001101010",
74779=>"101100011",
74780=>"110100100",
74781=>"000000000",
74782=>"001000000",
74783=>"000101100",
74784=>"110000001",
74785=>"010101111",
74786=>"010010010",
74787=>"111100101",
74788=>"101100000",
74789=>"111010111",
74790=>"000111000",
74791=>"011111111",
74792=>"100111111",
74793=>"111111000",
74794=>"101101111",
74795=>"111000000",
74796=>"101100011",
74797=>"101111000",
74798=>"001110110",
74799=>"000011101",
74800=>"000010010",
74801=>"101101000",
74802=>"001000000",
74803=>"001010010",
74804=>"111101001",
74805=>"001111111",
74806=>"001001001",
74807=>"010010111",
74808=>"111111010",
74809=>"000000100",
74810=>"000000101",
74811=>"101101111",
74812=>"011000000",
74813=>"111111111",
74814=>"000000000",
74815=>"001000100",
74816=>"100111101",
74817=>"110000001",
74818=>"101100100",
74819=>"100100100",
74820=>"010000000",
74821=>"000000000",
74822=>"111110101",
74823=>"000101111",
74824=>"000000001",
74825=>"101010010",
74826=>"000000000",
74827=>"101000110",
74828=>"111001000",
74829=>"001000000",
74830=>"110011001",
74831=>"110111111",
74832=>"111000110",
74833=>"000111111",
74834=>"000000111",
74835=>"100100100",
74836=>"101111011",
74837=>"100101000",
74838=>"101100001",
74839=>"100100100",
74840=>"110010011",
74841=>"001001001",
74842=>"000010011",
74843=>"010011010",
74844=>"111000000",
74845=>"000000101",
74846=>"100001110",
74847=>"001001001",
74848=>"011011000",
74849=>"010010011",
74850=>"100100001",
74851=>"010111110",
74852=>"000001100",
74853=>"101001000",
74854=>"100111111",
74855=>"101100111",
74856=>"010001000",
74857=>"111101101",
74858=>"111111111",
74859=>"000000011",
74860=>"010001010",
74861=>"000011110",
74862=>"111011011",
74863=>"001000011",
74864=>"000000001",
74865=>"111111111",
74866=>"100100100",
74867=>"111011000",
74868=>"111101000",
74869=>"010000000",
74870=>"101010110",
74871=>"000010000",
74872=>"000000000",
74873=>"101001101",
74874=>"110010110",
74875=>"010000111",
74876=>"011110100",
74877=>"001000001",
74878=>"111000000",
74879=>"000000110",
74880=>"110000101",
74881=>"000000011",
74882=>"111010110",
74883=>"111011110",
74884=>"100000001",
74885=>"111010010",
74886=>"111110110",
74887=>"110010000",
74888=>"000001011",
74889=>"100110010",
74890=>"100010001",
74891=>"011101110",
74892=>"010111100",
74893=>"110010000",
74894=>"101101100",
74895=>"001000010",
74896=>"000100100",
74897=>"111111111",
74898=>"010010100",
74899=>"110110110",
74900=>"010011111",
74901=>"101101101",
74902=>"101101111",
74903=>"001001001",
74904=>"111111011",
74905=>"011000001",
74906=>"001011000",
74907=>"000101001",
74908=>"011111011",
74909=>"011010010",
74910=>"111101111",
74911=>"111111011",
74912=>"001100100",
74913=>"001000000",
74914=>"100001101",
74915=>"111010111",
74916=>"101011100",
74917=>"011010000",
74918=>"001110111",
74919=>"110100100",
74920=>"000111111",
74921=>"111111111",
74922=>"000000100",
74923=>"101101101",
74924=>"000100110",
74925=>"000000001",
74926=>"011011001",
74927=>"010011010",
74928=>"010000110",
74929=>"011010100",
74930=>"100101100",
74931=>"111100100",
74932=>"010011011",
74933=>"100111010",
74934=>"000010001",
74935=>"100000001",
74936=>"000000000",
74937=>"001011000",
74938=>"111010111",
74939=>"011101100",
74940=>"000000000",
74941=>"111111000",
74942=>"110100011",
74943=>"100010000",
74944=>"000101101",
74945=>"010010010",
74946=>"000101111",
74947=>"100101110",
74948=>"111101100",
74949=>"110111011",
74950=>"011011111",
74951=>"010100101",
74952=>"101100101",
74953=>"000011010",
74954=>"010101101",
74955=>"001000001",
74956=>"011101001",
74957=>"110011001",
74958=>"111100100",
74959=>"001101111",
74960=>"010111111",
74961=>"110111100",
74962=>"001010011",
74963=>"011010010",
74964=>"111101101",
74965=>"110010111",
74966=>"111101101",
74967=>"001011001",
74968=>"010010000",
74969=>"000101111",
74970=>"111001011",
74971=>"011010010",
74972=>"101101001",
74973=>"101000000",
74974=>"111000010",
74975=>"000000010",
74976=>"001100000",
74977=>"000000010",
74978=>"100110111",
74979=>"011011110",
74980=>"000000000",
74981=>"010111110",
74982=>"011000000",
74983=>"100100000",
74984=>"000000000",
74985=>"111000000",
74986=>"011011001",
74987=>"001110100",
74988=>"011001000",
74989=>"011001001",
74990=>"000000110",
74991=>"000000011",
74992=>"011000000",
74993=>"101110100",
74994=>"001010000",
74995=>"100100000",
74996=>"110101000",
74997=>"111110110",
74998=>"100000010",
74999=>"101001011",
75000=>"111000000",
75001=>"101010000",
75002=>"111100000",
75003=>"001101101",
75004=>"101101000",
75005=>"001000101",
75006=>"111111011",
75007=>"110100110",
75008=>"111100101",
75009=>"000111000",
75010=>"000001111",
75011=>"101110110",
75012=>"001001000",
75013=>"111011000",
75014=>"100001111",
75015=>"110110000",
75016=>"000101101",
75017=>"000111000",
75018=>"110111111",
75019=>"001101111",
75020=>"101111011",
75021=>"000000010",
75022=>"101111001",
75023=>"000111110",
75024=>"100001111",
75025=>"001001111",
75026=>"000001111",
75027=>"100000010",
75028=>"111001111",
75029=>"010110100",
75030=>"011000001",
75031=>"111010000",
75032=>"101000111",
75033=>"011001111",
75034=>"100100111",
75035=>"000000000",
75036=>"011110111",
75037=>"110111111",
75038=>"101001011",
75039=>"000111111",
75040=>"001010110",
75041=>"000000001",
75042=>"000110111",
75043=>"110110000",
75044=>"001000100",
75045=>"010101111",
75046=>"010111000",
75047=>"011111000",
75048=>"000101111",
75049=>"111110000",
75050=>"010000000",
75051=>"000000111",
75052=>"001001011",
75053=>"000111111",
75054=>"001111010",
75055=>"100001101",
75056=>"000000101",
75057=>"111011111",
75058=>"000000101",
75059=>"001101111",
75060=>"001000000",
75061=>"111001011",
75062=>"110010011",
75063=>"010000000",
75064=>"000000110",
75065=>"101111101",
75066=>"000101010",
75067=>"100000111",
75068=>"010001111",
75069=>"111111000",
75070=>"000000111",
75071=>"111011100",
75072=>"011111101",
75073=>"101111010",
75074=>"111111100",
75075=>"011100000",
75076=>"010011011",
75077=>"010010000",
75078=>"000101111",
75079=>"110101001",
75080=>"101111100",
75081=>"101111111",
75082=>"111000000",
75083=>"000000111",
75084=>"110010000",
75085=>"100110000",
75086=>"001110100",
75087=>"101011111",
75088=>"111000001",
75089=>"011000000",
75090=>"000011101",
75091=>"001001000",
75092=>"000001001",
75093=>"101111111",
75094=>"001000000",
75095=>"001001111",
75096=>"111111111",
75097=>"000001011",
75098=>"011111110",
75099=>"000000101",
75100=>"111000000",
75101=>"000001011",
75102=>"000001101",
75103=>"001000100",
75104=>"111110000",
75105=>"010111010",
75106=>"111011011",
75107=>"001111001",
75108=>"100100000",
75109=>"100000000",
75110=>"110110110",
75111=>"001111110",
75112=>"011101001",
75113=>"110000000",
75114=>"001000000",
75115=>"101101000",
75116=>"110111011",
75117=>"000111001",
75118=>"101111010",
75119=>"010011111",
75120=>"000011000",
75121=>"000000110",
75122=>"000100110",
75123=>"111010000",
75124=>"000001110",
75125=>"000000000",
75126=>"000000111",
75127=>"001111010",
75128=>"000000000",
75129=>"010000000",
75130=>"000000001",
75131=>"101001011",
75132=>"001011110",
75133=>"100100100",
75134=>"000011111",
75135=>"111001011",
75136=>"110010000",
75137=>"100111111",
75138=>"110100010",
75139=>"010100101",
75140=>"010111111",
75141=>"101001000",
75142=>"100100110",
75143=>"100000000",
75144=>"100101100",
75145=>"000000011",
75146=>"111100111",
75147=>"111000000",
75148=>"000000010",
75149=>"011001000",
75150=>"000000001",
75151=>"000100001",
75152=>"011111100",
75153=>"111001000",
75154=>"000010111",
75155=>"110000000",
75156=>"100101000",
75157=>"001001000",
75158=>"000010111",
75159=>"011011000",
75160=>"111111101",
75161=>"000111111",
75162=>"101110111",
75163=>"111111000",
75164=>"000000010",
75165=>"111000000",
75166=>"110000000",
75167=>"110111000",
75168=>"101111111",
75169=>"000000100",
75170=>"111110000",
75171=>"101011111",
75172=>"000110000",
75173=>"010000011",
75174=>"110010001",
75175=>"110010000",
75176=>"001100101",
75177=>"000000000",
75178=>"101111111",
75179=>"111111010",
75180=>"101010000",
75181=>"011001111",
75182=>"110011111",
75183=>"001001011",
75184=>"110000100",
75185=>"001000001",
75186=>"101111111",
75187=>"000111111",
75188=>"001100100",
75189=>"000111111",
75190=>"100111000",
75191=>"000101110",
75192=>"100100111",
75193=>"111111011",
75194=>"110101000",
75195=>"101000000",
75196=>"000101111",
75197=>"111111111",
75198=>"111110110",
75199=>"000000010",
75200=>"000000111",
75201=>"000000111",
75202=>"000111010",
75203=>"000100100",
75204=>"000000000",
75205=>"100000000",
75206=>"000110110",
75207=>"110010000",
75208=>"000000110",
75209=>"000000000",
75210=>"101000100",
75211=>"001001111",
75212=>"110100100",
75213=>"001100110",
75214=>"000010111",
75215=>"111000010",
75216=>"000010111",
75217=>"110110010",
75218=>"101010000",
75219=>"010000001",
75220=>"001011110",
75221=>"100000000",
75222=>"111111100",
75223=>"000010100",
75224=>"111100000",
75225=>"100000111",
75226=>"001001111",
75227=>"101001000",
75228=>"001100111",
75229=>"001111111",
75230=>"111110000",
75231=>"000000101",
75232=>"111001011",
75233=>"000101101",
75234=>"100111000",
75235=>"011101010",
75236=>"000000011",
75237=>"000000000",
75238=>"111110111",
75239=>"111001100",
75240=>"111111110",
75241=>"001000110",
75242=>"011011111",
75243=>"000000001",
75244=>"111000000",
75245=>"111110010",
75246=>"000000000",
75247=>"001000010",
75248=>"111010000",
75249=>"001000000",
75250=>"111000000",
75251=>"000000000",
75252=>"001001011",
75253=>"100000011",
75254=>"000000000",
75255=>"100000000",
75256=>"001000110",
75257=>"101110101",
75258=>"100100111",
75259=>"010000000",
75260=>"000000000",
75261=>"101100111",
75262=>"001001000",
75263=>"111001000",
75264=>"110010000",
75265=>"110001110",
75266=>"001001101",
75267=>"110100100",
75268=>"011010001",
75269=>"110110000",
75270=>"111001010",
75271=>"100000111",
75272=>"110110110",
75273=>"000001111",
75274=>"101001011",
75275=>"110111001",
75276=>"110100000",
75277=>"100100110",
75278=>"000100110",
75279=>"000001000",
75280=>"111000000",
75281=>"001001111",
75282=>"010000111",
75283=>"011110110",
75284=>"101111110",
75285=>"110111011",
75286=>"110110110",
75287=>"000111111",
75288=>"011001001",
75289=>"111001001",
75290=>"110110000",
75291=>"011001001",
75292=>"000001111",
75293=>"000001111",
75294=>"110110001",
75295=>"000110110",
75296=>"000000011",
75297=>"110110111",
75298=>"110001111",
75299=>"100110110",
75300=>"001001010",
75301=>"011000000",
75302=>"110110100",
75303=>"110110110",
75304=>"001001111",
75305=>"100110100",
75306=>"001001111",
75307=>"100000011",
75308=>"001011111",
75309=>"001000001",
75310=>"110110010",
75311=>"000011111",
75312=>"001000110",
75313=>"111111011",
75314=>"101001000",
75315=>"001001011",
75316=>"001001111",
75317=>"111111101",
75318=>"000110011",
75319=>"000001001",
75320=>"000110111",
75321=>"001001001",
75322=>"000101000",
75323=>"000101111",
75324=>"001010000",
75325=>"110111000",
75326=>"000000001",
75327=>"110111000",
75328=>"101111111",
75329=>"110111011",
75330=>"001000111",
75331=>"100111000",
75332=>"110110100",
75333=>"000000101",
75334=>"000000110",
75335=>"010111001",
75336=>"111010111",
75337=>"000000000",
75338=>"001001111",
75339=>"100111111",
75340=>"100110000",
75341=>"111111100",
75342=>"100100000",
75343=>"000001111",
75344=>"111111001",
75345=>"100001000",
75346=>"110110000",
75347=>"110011101",
75348=>"111001001",
75349=>"111111111",
75350=>"011000001",
75351=>"001111111",
75352=>"000110100",
75353=>"001011111",
75354=>"101001010",
75355=>"110111000",
75356=>"001000111",
75357=>"000010010",
75358=>"111001001",
75359=>"111110000",
75360=>"100110000",
75361=>"110111111",
75362=>"101000101",
75363=>"011011111",
75364=>"011001011",
75365=>"110001000",
75366=>"000001111",
75367=>"000000110",
75368=>"001100010",
75369=>"110000000",
75370=>"010000001",
75371=>"110110001",
75372=>"011001001",
75373=>"001001001",
75374=>"110110110",
75375=>"101000000",
75376=>"111111011",
75377=>"000000111",
75378=>"000000100",
75379=>"110111000",
75380=>"000000001",
75381=>"001000000",
75382=>"100000001",
75383=>"110111100",
75384=>"001001001",
75385=>"110000000",
75386=>"110100000",
75387=>"100110110",
75388=>"010000000",
75389=>"111001000",
75390=>"011011111",
75391=>"110000000",
75392=>"000001110",
75393=>"110111000",
75394=>"110110110",
75395=>"110100000",
75396=>"110110110",
75397=>"001011111",
75398=>"000010011",
75399=>"000100000",
75400=>"100101100",
75401=>"000000100",
75402=>"000000000",
75403=>"110011000",
75404=>"111001001",
75405=>"010000100",
75406=>"000000000",
75407=>"000000111",
75408=>"111101001",
75409=>"011011111",
75410=>"001001110",
75411=>"110000000",
75412=>"000000000",
75413=>"100100111",
75414=>"110110101",
75415=>"110111000",
75416=>"001000001",
75417=>"001011110",
75418=>"001001111",
75419=>"100001101",
75420=>"000010000",
75421=>"000100100",
75422=>"111111111",
75423=>"000000000",
75424=>"000011101",
75425=>"000011011",
75426=>"011001111",
75427=>"000110001",
75428=>"110110100",
75429=>"111111101",
75430=>"100110000",
75431=>"001001111",
75432=>"011000001",
75433=>"101000000",
75434=>"000000110",
75435=>"010000110",
75436=>"110000001",
75437=>"110110000",
75438=>"101111111",
75439=>"100111100",
75440=>"000000000",
75441=>"110010011",
75442=>"111001001",
75443=>"111001000",
75444=>"011110111",
75445=>"000011111",
75446=>"000011001",
75447=>"000001000",
75448=>"010110100",
75449=>"010010001",
75450=>"110110111",
75451=>"111001001",
75452=>"001011000",
75453=>"111111010",
75454=>"110110000",
75455=>"000110110",
75456=>"000000111",
75457=>"001001001",
75458=>"110110110",
75459=>"000000000",
75460=>"001001111",
75461=>"111001110",
75462=>"000101111",
75463=>"000001111",
75464=>"011111101",
75465=>"000000000",
75466=>"000011111",
75467=>"110000110",
75468=>"100000111",
75469=>"000001001",
75470=>"001001001",
75471=>"110000011",
75472=>"110110110",
75473=>"110110110",
75474=>"110000001",
75475=>"110001000",
75476=>"111001000",
75477=>"101011001",
75478=>"011110110",
75479=>"001111111",
75480=>"001001011",
75481=>"110100001",
75482=>"110100000",
75483=>"001001011",
75484=>"111111111",
75485=>"110110110",
75486=>"111110010",
75487=>"011001011",
75488=>"000001010",
75489=>"011000000",
75490=>"111000000",
75491=>"011111001",
75492=>"001001011",
75493=>"110110000",
75494=>"110110110",
75495=>"100110010",
75496=>"110001000",
75497=>"010000000",
75498=>"001001000",
75499=>"000111111",
75500=>"000000000",
75501=>"110010000",
75502=>"010010000",
75503=>"000000000",
75504=>"000000000",
75505=>"001001111",
75506=>"010000100",
75507=>"000110100",
75508=>"111111001",
75509=>"001001001",
75510=>"000011000",
75511=>"111101101",
75512=>"001001111",
75513=>"000010110",
75514=>"100001000",
75515=>"010001101",
75516=>"011001001",
75517=>"000001000",
75518=>"111100000",
75519=>"001001101",
75520=>"001000111",
75521=>"111001000",
75522=>"000000000",
75523=>"111000001",
75524=>"110100101",
75525=>"111000101",
75526=>"111111111",
75527=>"000101000",
75528=>"101101100",
75529=>"111101111",
75530=>"001100001",
75531=>"001101110",
75532=>"000011100",
75533=>"111111000",
75534=>"011011000",
75535=>"110111111",
75536=>"111000101",
75537=>"010111000",
75538=>"010100110",
75539=>"000000111",
75540=>"111001111",
75541=>"111111001",
75542=>"000111101",
75543=>"010000000",
75544=>"101000000",
75545=>"011000011",
75546=>"111101111",
75547=>"001001101",
75548=>"000000000",
75549=>"000011011",
75550=>"110000110",
75551=>"000111111",
75552=>"111100000",
75553=>"101100011",
75554=>"000001010",
75555=>"000000000",
75556=>"101000001",
75557=>"100000111",
75558=>"010001011",
75559=>"110001001",
75560=>"101111010",
75561=>"000011011",
75562=>"010101100",
75563=>"100100000",
75564=>"001011101",
75565=>"110010111",
75566=>"111101011",
75567=>"011111010",
75568=>"111101000",
75569=>"100100101",
75570=>"000010011",
75571=>"110110110",
75572=>"000000000",
75573=>"010111110",
75574=>"111111111",
75575=>"011000001",
75576=>"100001111",
75577=>"101101111",
75578=>"001111111",
75579=>"000000101",
75580=>"001100110",
75581=>"110111000",
75582=>"101101100",
75583=>"101101000",
75584=>"111111010",
75585=>"100101111",
75586=>"111010000",
75587=>"011000100",
75588=>"010111010",
75589=>"101000101",
75590=>"110000100",
75591=>"100111011",
75592=>"011111000",
75593=>"110101000",
75594=>"000000000",
75595=>"000000111",
75596=>"110000001",
75597=>"100000101",
75598=>"111001001",
75599=>"100000101",
75600=>"000110000",
75601=>"111111010",
75602=>"000111010",
75603=>"000011011",
75604=>"000010011",
75605=>"100101101",
75606=>"001101100",
75607=>"101000111",
75608=>"001111110",
75609=>"000010101",
75610=>"110011001",
75611=>"101111011",
75612=>"100000111",
75613=>"100000100",
75614=>"010111101",
75615=>"111001001",
75616=>"111101101",
75617=>"001110010",
75618=>"101101001",
75619=>"011110100",
75620=>"100000101",
75621=>"101111010",
75622=>"111010000",
75623=>"000110111",
75624=>"001111010",
75625=>"110101010",
75626=>"000000011",
75627=>"111000001",
75628=>"110001000",
75629=>"000011110",
75630=>"101101010",
75631=>"111111011",
75632=>"100000111",
75633=>"000101001",
75634=>"110111111",
75635=>"101111010",
75636=>"100111111",
75637=>"111011101",
75638=>"111011001",
75639=>"111111001",
75640=>"110110110",
75641=>"000000111",
75642=>"000000001",
75643=>"101110000",
75644=>"011100001",
75645=>"000000110",
75646=>"000010010",
75647=>"001111111",
75648=>"011001001",
75649=>"111101000",
75650=>"000000000",
75651=>"000010000",
75652=>"000100111",
75653=>"111110000",
75654=>"001001111",
75655=>"011000000",
75656=>"001001001",
75657=>"111000011",
75658=>"000010010",
75659=>"010110100",
75660=>"101000000",
75661=>"001100001",
75662=>"000111111",
75663=>"110000010",
75664=>"001000001",
75665=>"111101100",
75666=>"110000100",
75667=>"011000000",
75668=>"000001110",
75669=>"101001000",
75670=>"101001001",
75671=>"001100100",
75672=>"101000000",
75673=>"001010010",
75674=>"000111111",
75675=>"010010000",
75676=>"000001001",
75677=>"111000100",
75678=>"011111111",
75679=>"100001001",
75680=>"101000100",
75681=>"111111101",
75682=>"000110000",
75683=>"000010010",
75684=>"111111111",
75685=>"000001001",
75686=>"111111111",
75687=>"101101011",
75688=>"011111001",
75689=>"110110111",
75690=>"101101101",
75691=>"001000000",
75692=>"010010000",
75693=>"111101001",
75694=>"000000001",
75695=>"101011000",
75696=>"011000000",
75697=>"110001001",
75698=>"000000000",
75699=>"000001000",
75700=>"010111111",
75701=>"011111011",
75702=>"101101101",
75703=>"000000011",
75704=>"100000001",
75705=>"010010000",
75706=>"110010111",
75707=>"000000101",
75708=>"101111111",
75709=>"011111101",
75710=>"111000101",
75711=>"000101110",
75712=>"111000010",
75713=>"001000111",
75714=>"000110001",
75715=>"100000111",
75716=>"000010110",
75717=>"001000101",
75718=>"011111000",
75719=>"111111101",
75720=>"010000010",
75721=>"001011001",
75722=>"110111101",
75723=>"111001001",
75724=>"001100000",
75725=>"111101101",
75726=>"000000101",
75727=>"111111101",
75728=>"111110110",
75729=>"000001001",
75730=>"010010010",
75731=>"110011010",
75732=>"101101101",
75733=>"100000000",
75734=>"101101101",
75735=>"000110011",
75736=>"101101101",
75737=>"111010010",
75738=>"110011010",
75739=>"111101000",
75740=>"000111001",
75741=>"111000000",
75742=>"000101111",
75743=>"101001000",
75744=>"000010010",
75745=>"111011101",
75746=>"000010011",
75747=>"110000000",
75748=>"101000000",
75749=>"111001010",
75750=>"111001110",
75751=>"000000000",
75752=>"100111101",
75753=>"100001000",
75754=>"101001000",
75755=>"101111101",
75756=>"101001000",
75757=>"000001101",
75758=>"100101110",
75759=>"101000000",
75760=>"101100100",
75761=>"100000111",
75762=>"101101001",
75763=>"011110110",
75764=>"100010110",
75765=>"101010011",
75766=>"000000001",
75767=>"011111010",
75768=>"101101101",
75769=>"010010000",
75770=>"000000111",
75771=>"111011110",
75772=>"100101101",
75773=>"000100000",
75774=>"001100101",
75775=>"001000010",
75776=>"101001001",
75777=>"000000000",
75778=>"101100101",
75779=>"000000110",
75780=>"101111110",
75781=>"011000000",
75782=>"111110000",
75783=>"110000111",
75784=>"101011010",
75785=>"000001000",
75786=>"001100110",
75787=>"110010000",
75788=>"000100101",
75789=>"100111110",
75790=>"100001001",
75791=>"000001111",
75792=>"110111010",
75793=>"100111000",
75794=>"111010101",
75795=>"000000011",
75796=>"001001000",
75797=>"010000100",
75798=>"000111111",
75799=>"111100111",
75800=>"111100111",
75801=>"011011001",
75802=>"010000000",
75803=>"011000000",
75804=>"111110100",
75805=>"111101010",
75806=>"101111111",
75807=>"100000000",
75808=>"111111111",
75809=>"111010010",
75810=>"101101100",
75811=>"010100110",
75812=>"111100100",
75813=>"001100000",
75814=>"110010000",
75815=>"000111110",
75816=>"111000000",
75817=>"110000001",
75818=>"000111111",
75819=>"010111111",
75820=>"010001001",
75821=>"100000111",
75822=>"100000000",
75823=>"101001111",
75824=>"000000010",
75825=>"111111111",
75826=>"100001001",
75827=>"000000001",
75828=>"111110000",
75829=>"000010101",
75830=>"100011011",
75831=>"110101101",
75832=>"110000101",
75833=>"000000000",
75834=>"111010010",
75835=>"111000000",
75836=>"010111110",
75837=>"111101101",
75838=>"000000000",
75839=>"001011111",
75840=>"110010111",
75841=>"111000000",
75842=>"011100111",
75843=>"000100110",
75844=>"111111010",
75845=>"111001101",
75846=>"000111010",
75847=>"000000000",
75848=>"111110000",
75849=>"000111010",
75850=>"100001101",
75851=>"010110110",
75852=>"111011000",
75853=>"000001000",
75854=>"111111111",
75855=>"000101111",
75856=>"111111100",
75857=>"100010001",
75858=>"100000010",
75859=>"111101101",
75860=>"101101111",
75861=>"010111111",
75862=>"110110010",
75863=>"000111111",
75864=>"111111111",
75865=>"011000010",
75866=>"010110110",
75867=>"011110000",
75868=>"010000000",
75869=>"001001011",
75870=>"010000111",
75871=>"000011011",
75872=>"000000000",
75873=>"010110000",
75874=>"001101111",
75875=>"001011000",
75876=>"100101000",
75877=>"101011011",
75878=>"110000000",
75879=>"000001111",
75880=>"110010111",
75881=>"010111101",
75882=>"000000111",
75883=>"111001000",
75884=>"111100101",
75885=>"000010111",
75886=>"011010011",
75887=>"010000000",
75888=>"011100000",
75889=>"111000000",
75890=>"110110110",
75891=>"000000111",
75892=>"000000111",
75893=>"001000000",
75894=>"010000010",
75895=>"000101000",
75896=>"000000111",
75897=>"000000111",
75898=>"100000010",
75899=>"001001000",
75900=>"000110110",
75901=>"101100110",
75902=>"000001111",
75903=>"101101000",
75904=>"000000010",
75905=>"111100100",
75906=>"000000000",
75907=>"001000111",
75908=>"101000100",
75909=>"100000000",
75910=>"001001000",
75911=>"010011000",
75912=>"101001001",
75913=>"110111000",
75914=>"000001000",
75915=>"001100111",
75916=>"111100101",
75917=>"000000100",
75918=>"111111111",
75919=>"000000001",
75920=>"101101111",
75921=>"111001000",
75922=>"111011000",
75923=>"110010110",
75924=>"110111111",
75925=>"000111111",
75926=>"110111111",
75927=>"000000000",
75928=>"111111110",
75929=>"000111111",
75930=>"010100100",
75931=>"100000110",
75932=>"000011011",
75933=>"101000000",
75934=>"000000110",
75935=>"001001000",
75936=>"101011101",
75937=>"010010011",
75938=>"000101111",
75939=>"111010111",
75940=>"000000010",
75941=>"110001000",
75942=>"101001000",
75943=>"010010100",
75944=>"000000110",
75945=>"010111111",
75946=>"101000001",
75947=>"110010000",
75948=>"010011111",
75949=>"100000000",
75950=>"101111000",
75951=>"000011000",
75952=>"010010001",
75953=>"011111110",
75954=>"000000010",
75955=>"001101100",
75956=>"110100100",
75957=>"000100111",
75958=>"010100111",
75959=>"000110111",
75960=>"000001011",
75961=>"111111111",
75962=>"001010010",
75963=>"000000111",
75964=>"000000101",
75965=>"111101111",
75966=>"100100000",
75967=>"110110101",
75968=>"000000000",
75969=>"111000000",
75970=>"010000110",
75971=>"111101100",
75972=>"001000111",
75973=>"111111010",
75974=>"011000011",
75975=>"111001000",
75976=>"101111111",
75977=>"111010000",
75978=>"100101111",
75979=>"111101011",
75980=>"111011001",
75981=>"010011011",
75982=>"001111111",
75983=>"001000010",
75984=>"010000000",
75985=>"101100000",
75986=>"110010110",
75987=>"101111101",
75988=>"110000000",
75989=>"111111001",
75990=>"001000000",
75991=>"111000011",
75992=>"000000111",
75993=>"100000000",
75994=>"101011000",
75995=>"111010111",
75996=>"011111101",
75997=>"000011111",
75998=>"010000101",
75999=>"000000000",
76000=>"000000000",
76001=>"101000010",
76002=>"000000000",
76003=>"011111100",
76004=>"111100000",
76005=>"111000101",
76006=>"101101111",
76007=>"101110010",
76008=>"100000000",
76009=>"010000100",
76010=>"000100000",
76011=>"010110111",
76012=>"011001000",
76013=>"100000000",
76014=>"000000000",
76015=>"000010000",
76016=>"111011100",
76017=>"111111100",
76018=>"011000100",
76019=>"111101100",
76020=>"100110000",
76021=>"100100100",
76022=>"000000000",
76023=>"111001011",
76024=>"011110111",
76025=>"000111111",
76026=>"001000000",
76027=>"111111000",
76028=>"000000001",
76029=>"000000110",
76030=>"010010001",
76031=>"000000000",
76032=>"110011000",
76033=>"000100111",
76034=>"101000001",
76035=>"000000110",
76036=>"001001010",
76037=>"100000000",
76038=>"110111010",
76039=>"010100000",
76040=>"110110110",
76041=>"001000100",
76042=>"000000100",
76043=>"000000000",
76044=>"001000000",
76045=>"111110110",
76046=>"001011011",
76047=>"110000000",
76048=>"011001111",
76049=>"000000001",
76050=>"000000000",
76051=>"000111111",
76052=>"111001101",
76053=>"000000000",
76054=>"001111111",
76055=>"100100111",
76056=>"101000100",
76057=>"000111001",
76058=>"011000000",
76059=>"111101000",
76060=>"000001110",
76061=>"000000101",
76062=>"111001000",
76063=>"010000000",
76064=>"110101100",
76065=>"011101000",
76066=>"001100010",
76067=>"000000000",
76068=>"001011111",
76069=>"111111111",
76070=>"000000001",
76071=>"000000111",
76072=>"111111110",
76073=>"111111100",
76074=>"000000000",
76075=>"110101111",
76076=>"010111011",
76077=>"000000111",
76078=>"101111001",
76079=>"000100000",
76080=>"000000111",
76081=>"001001001",
76082=>"001100000",
76083=>"111111111",
76084=>"110000111",
76085=>"111110111",
76086=>"010100101",
76087=>"000000000",
76088=>"110000000",
76089=>"000001101",
76090=>"101000101",
76091=>"000100100",
76092=>"100010101",
76093=>"111111111",
76094=>"100000001",
76095=>"110111010",
76096=>"110001000",
76097=>"001101000",
76098=>"000001010",
76099=>"110010100",
76100=>"000110111",
76101=>"110001111",
76102=>"111000111",
76103=>"011110000",
76104=>"000000011",
76105=>"010001000",
76106=>"111001111",
76107=>"110000000",
76108=>"000100110",
76109=>"011100011",
76110=>"000111100",
76111=>"011011011",
76112=>"111111010",
76113=>"010011010",
76114=>"001110111",
76115=>"011001001",
76116=>"000000000",
76117=>"111011111",
76118=>"100100100",
76119=>"000000000",
76120=>"111100000",
76121=>"000011010",
76122=>"000000000",
76123=>"110110000",
76124=>"000010000",
76125=>"011001001",
76126=>"000010010",
76127=>"000001001",
76128=>"010111110",
76129=>"111111101",
76130=>"101000101",
76131=>"000000000",
76132=>"000001000",
76133=>"111011011",
76134=>"111110000",
76135=>"000100000",
76136=>"110000111",
76137=>"000000000",
76138=>"110000001",
76139=>"100001000",
76140=>"101111111",
76141=>"000100001",
76142=>"111011011",
76143=>"110000000",
76144=>"111111111",
76145=>"010000111",
76146=>"110100101",
76147=>"100111111",
76148=>"100110111",
76149=>"000000100",
76150=>"110110110",
76151=>"111110010",
76152=>"000000000",
76153=>"111111010",
76154=>"111111100",
76155=>"001000001",
76156=>"100100110",
76157=>"111101001",
76158=>"000001110",
76159=>"011000000",
76160=>"111111001",
76161=>"110100000",
76162=>"011011110",
76163=>"001000011",
76164=>"000000101",
76165=>"111111111",
76166=>"100111110",
76167=>"011100000",
76168=>"110111111",
76169=>"101111111",
76170=>"000000111",
76171=>"010000000",
76172=>"110110000",
76173=>"110110000",
76174=>"001000000",
76175=>"000000100",
76176=>"110100100",
76177=>"000001101",
76178=>"000000000",
76179=>"111001000",
76180=>"000001001",
76181=>"000000000",
76182=>"000001000",
76183=>"110011011",
76184=>"001110000",
76185=>"000000111",
76186=>"000000000",
76187=>"101000000",
76188=>"010111010",
76189=>"111111111",
76190=>"111000010",
76191=>"000000000",
76192=>"001101101",
76193=>"111001111",
76194=>"110111111",
76195=>"000111111",
76196=>"101001110",
76197=>"110111000",
76198=>"111111011",
76199=>"110111111",
76200=>"000111001",
76201=>"110001110",
76202=>"001000000",
76203=>"000000001",
76204=>"111100111",
76205=>"110111011",
76206=>"110101111",
76207=>"010111010",
76208=>"100010000",
76209=>"100100000",
76210=>"000000000",
76211=>"011101010",
76212=>"110110111",
76213=>"111001000",
76214=>"010111010",
76215=>"111111001",
76216=>"011110111",
76217=>"110110001",
76218=>"010010000",
76219=>"110111010",
76220=>"101111001",
76221=>"111111111",
76222=>"010011111",
76223=>"110111011",
76224=>"011000000",
76225=>"111000001",
76226=>"000000111",
76227=>"011011001",
76228=>"101110000",
76229=>"001111111",
76230=>"000000010",
76231=>"000000000",
76232=>"100101111",
76233=>"010010000",
76234=>"100110111",
76235=>"001000000",
76236=>"011000000",
76237=>"001011110",
76238=>"111000000",
76239=>"111101111",
76240=>"110101110",
76241=>"111111111",
76242=>"000110111",
76243=>"110111111",
76244=>"001000000",
76245=>"011000100",
76246=>"110110011",
76247=>"110100000",
76248=>"000000111",
76249=>"000000010",
76250=>"000000100",
76251=>"001000000",
76252=>"100111101",
76253=>"000100000",
76254=>"110111000",
76255=>"110001000",
76256=>"001000000",
76257=>"111001101",
76258=>"000000000",
76259=>"110111111",
76260=>"101011010",
76261=>"000111010",
76262=>"000110110",
76263=>"010011001",
76264=>"100111111",
76265=>"010010111",
76266=>"001000001",
76267=>"110110110",
76268=>"010010000",
76269=>"000101010",
76270=>"011000010",
76271=>"001000010",
76272=>"101100101",
76273=>"100001111",
76274=>"000001001",
76275=>"011000010",
76276=>"111100000",
76277=>"010110111",
76278=>"000000000",
76279=>"100000000",
76280=>"010000000",
76281=>"000010010",
76282=>"000000000",
76283=>"001110000",
76284=>"000000000",
76285=>"011001000",
76286=>"100100100",
76287=>"001000000",
76288=>"000100110",
76289=>"000010001",
76290=>"100000010",
76291=>"000000000",
76292=>"000010000",
76293=>"100000110",
76294=>"001001111",
76295=>"000010010",
76296=>"010011000",
76297=>"001000111",
76298=>"001001000",
76299=>"000001000",
76300=>"001000001",
76301=>"111111101",
76302=>"000011100",
76303=>"000000000",
76304=>"111000000",
76305=>"110100010",
76306=>"100000001",
76307=>"110101111",
76308=>"110011000",
76309=>"111100110",
76310=>"001000000",
76311=>"101001000",
76312=>"101000111",
76313=>"011111011",
76314=>"000000000",
76315=>"111000101",
76316=>"111000010",
76317=>"100000001",
76318=>"110111111",
76319=>"001110000",
76320=>"000010010",
76321=>"100001101",
76322=>"110101000",
76323=>"111010000",
76324=>"111000000",
76325=>"000011111",
76326=>"010110000",
76327=>"011110000",
76328=>"010110001",
76329=>"010010001",
76330=>"100110101",
76331=>"111110111",
76332=>"000000100",
76333=>"111101111",
76334=>"010010000",
76335=>"000000000",
76336=>"101111101",
76337=>"000000111",
76338=>"100010010",
76339=>"000101111",
76340=>"001000111",
76341=>"001011000",
76342=>"000001111",
76343=>"111001101",
76344=>"010000011",
76345=>"001101111",
76346=>"111101010",
76347=>"011000110",
76348=>"000011011",
76349=>"110111111",
76350=>"011000100",
76351=>"110110010",
76352=>"000010011",
76353=>"000010111",
76354=>"111010101",
76355=>"010000110",
76356=>"100101000",
76357=>"001001101",
76358=>"000001111",
76359=>"111111101",
76360=>"110000111",
76361=>"111110000",
76362=>"001001011",
76363=>"011011000",
76364=>"100000111",
76365=>"100100100",
76366=>"001000001",
76367=>"010100101",
76368=>"101101000",
76369=>"111111111",
76370=>"111111101",
76371=>"010111010",
76372=>"001100110",
76373=>"000000000",
76374=>"011000000",
76375=>"000000011",
76376=>"100000000",
76377=>"111111000",
76378=>"111011111",
76379=>"111111000",
76380=>"000000000",
76381=>"000011110",
76382=>"111111111",
76383=>"110000011",
76384=>"000010000",
76385=>"100000100",
76386=>"101001111",
76387=>"001100111",
76388=>"111111001",
76389=>"000000100",
76390=>"101111111",
76391=>"010010000",
76392=>"101001111",
76393=>"101101011",
76394=>"111010010",
76395=>"001111111",
76396=>"110110101",
76397=>"111111111",
76398=>"010000000",
76399=>"000000100",
76400=>"011011010",
76401=>"000000001",
76402=>"000000111",
76403=>"001010000",
76404=>"011000000",
76405=>"001101110",
76406=>"000000100",
76407=>"110000111",
76408=>"100001111",
76409=>"010000110",
76410=>"000001001",
76411=>"101111101",
76412=>"000000111",
76413=>"011101010",
76414=>"001010111",
76415=>"101101100",
76416=>"011001010",
76417=>"111010011",
76418=>"111101100",
76419=>"111111100",
76420=>"001001001",
76421=>"111011011",
76422=>"000111111",
76423=>"100000100",
76424=>"100101110",
76425=>"011001101",
76426=>"100000111",
76427=>"111110010",
76428=>"101101111",
76429=>"000000010",
76430=>"000000100",
76431=>"001001000",
76432=>"101101001",
76433=>"101111111",
76434=>"101000010",
76435=>"000111010",
76436=>"000000001",
76437=>"010000111",
76438=>"000100111",
76439=>"001111100",
76440=>"011010101",
76441=>"101111110",
76442=>"001000111",
76443=>"000000101",
76444=>"101111000",
76445=>"111001011",
76446=>"011000000",
76447=>"110110000",
76448=>"001001110",
76449=>"001000001",
76450=>"111011100",
76451=>"000010000",
76452=>"110111111",
76453=>"110101000",
76454=>"110110001",
76455=>"111010111",
76456=>"101000111",
76457=>"000010000",
76458=>"101100111",
76459=>"000000111",
76460=>"111111111",
76461=>"000000000",
76462=>"100001001",
76463=>"010111101",
76464=>"101000111",
76465=>"001000100",
76466=>"101101110",
76467=>"000110001",
76468=>"110111010",
76469=>"111111111",
76470=>"011100100",
76471=>"000011101",
76472=>"000100100",
76473=>"011000010",
76474=>"111010000",
76475=>"111101000",
76476=>"001011110",
76477=>"010010101",
76478=>"111111001",
76479=>"101011010",
76480=>"101001111",
76481=>"101000111",
76482=>"010010000",
76483=>"000000011",
76484=>"000000001",
76485=>"110000110",
76486=>"000011100",
76487=>"101000000",
76488=>"001111100",
76489=>"001001001",
76490=>"011011111",
76491=>"000000111",
76492=>"000000100",
76493=>"000000001",
76494=>"101101000",
76495=>"101101010",
76496=>"111101101",
76497=>"110110001",
76498=>"010000000",
76499=>"000000000",
76500=>"110000000",
76501=>"100000000",
76502=>"010000111",
76503=>"001011011",
76504=>"111010000",
76505=>"011111111",
76506=>"100101001",
76507=>"111001111",
76508=>"000000100",
76509=>"101111010",
76510=>"000100111",
76511=>"001000101",
76512=>"111101101",
76513=>"101100111",
76514=>"001010000",
76515=>"000100000",
76516=>"101000010",
76517=>"000000000",
76518=>"000000000",
76519=>"000000000",
76520=>"100100100",
76521=>"000111111",
76522=>"100000100",
76523=>"000101101",
76524=>"000000101",
76525=>"010001001",
76526=>"010000010",
76527=>"101000001",
76528=>"111001000",
76529=>"011010001",
76530=>"010111111",
76531=>"000110100",
76532=>"000011000",
76533=>"101001100",
76534=>"000100000",
76535=>"000110110",
76536=>"001101010",
76537=>"010101010",
76538=>"000000000",
76539=>"011000000",
76540=>"101001101",
76541=>"010010010",
76542=>"001111000",
76543=>"001010111",
76544=>"101100101",
76545=>"011000010",
76546=>"000010010",
76547=>"011000000",
76548=>"000001001",
76549=>"001011010",
76550=>"111111111",
76551=>"010111000",
76552=>"001001001",
76553=>"101000010",
76554=>"000000000",
76555=>"000100110",
76556=>"011010000",
76557=>"000000011",
76558=>"110101000",
76559=>"101011100",
76560=>"111111011",
76561=>"111111010",
76562=>"111110011",
76563=>"000000000",
76564=>"001000110",
76565=>"111001001",
76566=>"111100110",
76567=>"010000000",
76568=>"010000100",
76569=>"011010010",
76570=>"000000111",
76571=>"001000110",
76572=>"000000011",
76573=>"001111100",
76574=>"000010010",
76575=>"101111101",
76576=>"000000101",
76577=>"000000000",
76578=>"011101111",
76579=>"000001000",
76580=>"000000000",
76581=>"000001111",
76582=>"000010011",
76583=>"001001101",
76584=>"011111001",
76585=>"000100011",
76586=>"010000001",
76587=>"001011011",
76588=>"001100101",
76589=>"100101110",
76590=>"111001111",
76591=>"111111111",
76592=>"111111111",
76593=>"000000001",
76594=>"010111100",
76595=>"000100110",
76596=>"101001111",
76597=>"111111110",
76598=>"010000011",
76599=>"001001101",
76600=>"101000000",
76601=>"000110000",
76602=>"000011110",
76603=>"011011111",
76604=>"000111011",
76605=>"011111011",
76606=>"000000000",
76607=>"100100110",
76608=>"001000110",
76609=>"000000011",
76610=>"000100000",
76611=>"101001011",
76612=>"101001011",
76613=>"111111011",
76614=>"011000111",
76615=>"111111011",
76616=>"000001000",
76617=>"111111111",
76618=>"000000000",
76619=>"001001101",
76620=>"111011111",
76621=>"000000001",
76622=>"000000000",
76623=>"101111111",
76624=>"000000000",
76625=>"111111000",
76626=>"000101111",
76627=>"000010011",
76628=>"000000110",
76629=>"001001111",
76630=>"000000010",
76631=>"000110101",
76632=>"000111111",
76633=>"000000011",
76634=>"101011001",
76635=>"000000011",
76636=>"000000010",
76637=>"001110100",
76638=>"111111100",
76639=>"111101000",
76640=>"111000000",
76641=>"000000010",
76642=>"000000000",
76643=>"111000100",
76644=>"011111011",
76645=>"000111000",
76646=>"100011000",
76647=>"111111111",
76648=>"111010111",
76649=>"111010111",
76650=>"010111001",
76651=>"111111011",
76652=>"000111011",
76653=>"110110000",
76654=>"000000001",
76655=>"000000011",
76656=>"000000100",
76657=>"000000000",
76658=>"101000100",
76659=>"010110100",
76660=>"111001001",
76661=>"001000010",
76662=>"111111011",
76663=>"111101101",
76664=>"000110010",
76665=>"000011101",
76666=>"000100101",
76667=>"101010110",
76668=>"001001000",
76669=>"000000100",
76670=>"001111101",
76671=>"000010001",
76672=>"001000000",
76673=>"001111011",
76674=>"100000000",
76675=>"111111011",
76676=>"010010001",
76677=>"101101101",
76678=>"000000110",
76679=>"000000101",
76680=>"000000001",
76681=>"000111111",
76682=>"000011010",
76683=>"111011010",
76684=>"001001000",
76685=>"001000011",
76686=>"011000001",
76687=>"101001001",
76688=>"100100000",
76689=>"111100000",
76690=>"001000000",
76691=>"000000000",
76692=>"000000000",
76693=>"110111100",
76694=>"101000110",
76695=>"000000001",
76696=>"000000110",
76697=>"000111111",
76698=>"000011000",
76699=>"000111001",
76700=>"000101100",
76701=>"111000101",
76702=>"001000010",
76703=>"000011011",
76704=>"000000101",
76705=>"111110000",
76706=>"111111101",
76707=>"001000000",
76708=>"010000000",
76709=>"000000111",
76710=>"000000000",
76711=>"111001111",
76712=>"000000111",
76713=>"000001000",
76714=>"111000010",
76715=>"000000000",
76716=>"111111111",
76717=>"111111111",
76718=>"000101011",
76719=>"011111000",
76720=>"001111101",
76721=>"001001100",
76722=>"001110000",
76723=>"000011011",
76724=>"111111011",
76725=>"111000101",
76726=>"000000001",
76727=>"000011111",
76728=>"000100100",
76729=>"001000001",
76730=>"010111101",
76731=>"100000111",
76732=>"111010111",
76733=>"001000000",
76734=>"100111011",
76735=>"000111111",
76736=>"011001010",
76737=>"000000111",
76738=>"111101101",
76739=>"000010010",
76740=>"000111000",
76741=>"000000100",
76742=>"000000000",
76743=>"000000101",
76744=>"001101101",
76745=>"001101001",
76746=>"111001001",
76747=>"000101000",
76748=>"000100000",
76749=>"100000001",
76750=>"110101000",
76751=>"001111111",
76752=>"111111110",
76753=>"000000111",
76754=>"001000000",
76755=>"111111010",
76756=>"000000000",
76757=>"111001001",
76758=>"001000000",
76759=>"100111111",
76760=>"000111111",
76761=>"000100111",
76762=>"000001001",
76763=>"000000000",
76764=>"111010111",
76765=>"111111111",
76766=>"111011111",
76767=>"111111010",
76768=>"000000110",
76769=>"110111010",
76770=>"111111000",
76771=>"100101111",
76772=>"010000000",
76773=>"011001000",
76774=>"001000101",
76775=>"000000001",
76776=>"110000000",
76777=>"000000001",
76778=>"100100111",
76779=>"110000000",
76780=>"111111111",
76781=>"100111011",
76782=>"000001000",
76783=>"111011011",
76784=>"001111111",
76785=>"000000011",
76786=>"001000010",
76787=>"100101101",
76788=>"011001011",
76789=>"000000000",
76790=>"010000010",
76791=>"111001001",
76792=>"010000001",
76793=>"111101101",
76794=>"000000000",
76795=>"001001001",
76796=>"000010010",
76797=>"000010000",
76798=>"001000000",
76799=>"111001011",
76800=>"111011101",
76801=>"111111111",
76802=>"000010010",
76803=>"100000000",
76804=>"110111111",
76805=>"111000111",
76806=>"110010111",
76807=>"000111011",
76808=>"100100000",
76809=>"000000000",
76810=>"100100100",
76811=>"001101111",
76812=>"111010000",
76813=>"110100101",
76814=>"100101100",
76815=>"111111101",
76816=>"000000000",
76817=>"000000100",
76818=>"011001000",
76819=>"011101111",
76820=>"000000100",
76821=>"000111111",
76822=>"011011001",
76823=>"101001100",
76824=>"000000000",
76825=>"000000010",
76826=>"100100101",
76827=>"111100000",
76828=>"100001111",
76829=>"001111111",
76830=>"001000000",
76831=>"000010111",
76832=>"000111011",
76833=>"100100000",
76834=>"000010110",
76835=>"100000010",
76836=>"000100111",
76837=>"011011101",
76838=>"001011111",
76839=>"111010000",
76840=>"111111111",
76841=>"111111110",
76842=>"100000100",
76843=>"011111010",
76844=>"111110011",
76845=>"100000110",
76846=>"111001000",
76847=>"111000000",
76848=>"000000111",
76849=>"010101111",
76850=>"101111100",
76851=>"000111110",
76852=>"011011001",
76853=>"111111000",
76854=>"011011001",
76855=>"000111011",
76856=>"111001000",
76857=>"000000000",
76858=>"101100100",
76859=>"000000111",
76860=>"100000000",
76861=>"010111011",
76862=>"001001111",
76863=>"010111110",
76864=>"111010000",
76865=>"000100000",
76866=>"111000000",
76867=>"111110000",
76868=>"000100011",
76869=>"101000100",
76870=>"100111011",
76871=>"100010111",
76872=>"000000011",
76873=>"101001011",
76874=>"101000000",
76875=>"000000000",
76876=>"111111011",
76877=>"000100110",
76878=>"000010110",
76879=>"000110111",
76880=>"000011111",
76881=>"110101000",
76882=>"011111111",
76883=>"111111111",
76884=>"111110010",
76885=>"011011011",
76886=>"000110101",
76887=>"101111111",
76888=>"100111110",
76889=>"000111000",
76890=>"100111111",
76891=>"101111110",
76892=>"100000000",
76893=>"000000001",
76894=>"111111111",
76895=>"111111100",
76896=>"111111111",
76897=>"000000001",
76898=>"111110011",
76899=>"000001101",
76900=>"000100000",
76901=>"010011100",
76902=>"111010010",
76903=>"000111111",
76904=>"001000100",
76905=>"010100100",
76906=>"011000000",
76907=>"010011111",
76908=>"000100000",
76909=>"000100111",
76910=>"000000010",
76911=>"111000111",
76912=>"000001011",
76913=>"000000000",
76914=>"110110110",
76915=>"001011000",
76916=>"000111011",
76917=>"011000111",
76918=>"111010000",
76919=>"111111111",
76920=>"000000000",
76921=>"000000111",
76922=>"111100000",
76923=>"101111000",
76924=>"000000000",
76925=>"101100111",
76926=>"001001001",
76927=>"000000000",
76928=>"101100000",
76929=>"010000000",
76930=>"111100000",
76931=>"011001000",
76932=>"000100011",
76933=>"101111010",
76934=>"110110110",
76935=>"000000110",
76936=>"010110110",
76937=>"000001001",
76938=>"000100110",
76939=>"111000100",
76940=>"101101101",
76941=>"100111111",
76942=>"111000000",
76943=>"111101001",
76944=>"101011111",
76945=>"111111000",
76946=>"000000001",
76947=>"000000000",
76948=>"001001111",
76949=>"101000000",
76950=>"111100000",
76951=>"000001001",
76952=>"111101101",
76953=>"101100000",
76954=>"000101110",
76955=>"111101111",
76956=>"001011101",
76957=>"000000000",
76958=>"000000110",
76959=>"001101111",
76960=>"100010011",
76961=>"011111111",
76962=>"100000110",
76963=>"000110000",
76964=>"111000000",
76965=>"001111111",
76966=>"001000101",
76967=>"111111010",
76968=>"000000101",
76969=>"011001101",
76970=>"010000100",
76971=>"010011101",
76972=>"100010000",
76973=>"111111110",
76974=>"110110110",
76975=>"100000010",
76976=>"111010000",
76977=>"000001011",
76978=>"110000101",
76979=>"000000100",
76980=>"101101010",
76981=>"111010110",
76982=>"001000000",
76983=>"000000110",
76984=>"001000000",
76985=>"000000111",
76986=>"111011111",
76987=>"101000111",
76988=>"000100110",
76989=>"111000010",
76990=>"000000000",
76991=>"000111000",
76992=>"000010010",
76993=>"101000100",
76994=>"111100010",
76995=>"000100000",
76996=>"101101100",
76997=>"000001111",
76998=>"111101010",
76999=>"001000101",
77000=>"011010111",
77001=>"111100000",
77002=>"010101110",
77003=>"101100000",
77004=>"100111111",
77005=>"000000000",
77006=>"101101101",
77007=>"000000101",
77008=>"010100000",
77009=>"110110111",
77010=>"011000100",
77011=>"110111101",
77012=>"010111001",
77013=>"000101111",
77014=>"010101000",
77015=>"000011101",
77016=>"011111010",
77017=>"000110110",
77018=>"010111100",
77019=>"000000111",
77020=>"110110010",
77021=>"100101000",
77022=>"010010100",
77023=>"111111111",
77024=>"100000000",
77025=>"010000000",
77026=>"111001110",
77027=>"000111101",
77028=>"000101101",
77029=>"000000000",
77030=>"010001000",
77031=>"001011111",
77032=>"111101001",
77033=>"000001001",
77034=>"001001001",
77035=>"111000100",
77036=>"110000000",
77037=>"000100100",
77038=>"000000000",
77039=>"110100000",
77040=>"000100011",
77041=>"000100111",
77042=>"011111011",
77043=>"000111111",
77044=>"111110011",
77045=>"000000111",
77046=>"000110111",
77047=>"001010000",
77048=>"100000000",
77049=>"111111101",
77050=>"000100100",
77051=>"000000010",
77052=>"100111000",
77053=>"000100101",
77054=>"010010111",
77055=>"111110000",
77056=>"111100110",
77057=>"010110011",
77058=>"101001101",
77059=>"100101111",
77060=>"100110110",
77061=>"100100101",
77062=>"111111011",
77063=>"111011010",
77064=>"110100000",
77065=>"100000000",
77066=>"101011101",
77067=>"100110100",
77068=>"110100100",
77069=>"110111001",
77070=>"100110000",
77071=>"010100111",
77072=>"100000100",
77073=>"111100111",
77074=>"000100111",
77075=>"000000001",
77076=>"111001111",
77077=>"110110011",
77078=>"111001000",
77079=>"001110000",
77080=>"100110110",
77081=>"000101011",
77082=>"110100110",
77083=>"100100000",
77084=>"011110110",
77085=>"011011001",
77086=>"110100011",
77087=>"101001000",
77088=>"110001101",
77089=>"100100110",
77090=>"000100110",
77091=>"110000010",
77092=>"000110111",
77093=>"110100110",
77094=>"000010111",
77095=>"100000100",
77096=>"010011100",
77097=>"000111100",
77098=>"111110110",
77099=>"001001000",
77100=>"001110110",
77101=>"001110111",
77102=>"001110110",
77103=>"110111111",
77104=>"011001001",
77105=>"110001000",
77106=>"000100100",
77107=>"111100011",
77108=>"100011011",
77109=>"110010000",
77110=>"000001011",
77111=>"110110100",
77112=>"011010110",
77113=>"100100100",
77114=>"111110010",
77115=>"101001000",
77116=>"000100100",
77117=>"110011011",
77118=>"100100000",
77119=>"000010011",
77120=>"101011100",
77121=>"010100110",
77122=>"011110000",
77123=>"100100100",
77124=>"011000000",
77125=>"110110000",
77126=>"000001010",
77127=>"001011101",
77128=>"101111110",
77129=>"110100100",
77130=>"110000011",
77131=>"100111111",
77132=>"000100000",
77133=>"111111111",
77134=>"101011001",
77135=>"011100000",
77136=>"100010010",
77137=>"101011111",
77138=>"111110001",
77139=>"001000000",
77140=>"111110111",
77141=>"110000110",
77142=>"111001001",
77143=>"101001001",
77144=>"001111111",
77145=>"000000001",
77146=>"100001001",
77147=>"101001001",
77148=>"101100100",
77149=>"100000000",
77150=>"000011011",
77151=>"100100111",
77152=>"100100100",
77153=>"000000000",
77154=>"100100100",
77155=>"111110110",
77156=>"011000000",
77157=>"101001100",
77158=>"100100100",
77159=>"001011011",
77160=>"110100010",
77161=>"100100000",
77162=>"000100110",
77163=>"011111010",
77164=>"111100100",
77165=>"001011000",
77166=>"010100100",
77167=>"101110110",
77168=>"111111011",
77169=>"100110110",
77170=>"111111101",
77171=>"001001000",
77172=>"011110111",
77173=>"100100000",
77174=>"100100001",
77175=>"000010111",
77176=>"011010111",
77177=>"001100111",
77178=>"000100010",
77179=>"011011000",
77180=>"011000000",
77181=>"001010010",
77182=>"011011011",
77183=>"100001000",
77184=>"101100111",
77185=>"101000100",
77186=>"001111011",
77187=>"111100100",
77188=>"111011011",
77189=>"011011111",
77190=>"000100100",
77191=>"100100100",
77192=>"100101111",
77193=>"111111100",
77194=>"001011000",
77195=>"010000000",
77196=>"100011011",
77197=>"100100000",
77198=>"000100100",
77199=>"100100100",
77200=>"010010000",
77201=>"100101100",
77202=>"100100110",
77203=>"111110110",
77204=>"011000000",
77205=>"101100100",
77206=>"110100100",
77207=>"100110010",
77208=>"011001000",
77209=>"001011011",
77210=>"100101011",
77211=>"011011001",
77212=>"111110110",
77213=>"100001100",
77214=>"011110011",
77215=>"110110110",
77216=>"101011101",
77217=>"000110000",
77218=>"011000001",
77219=>"100100111",
77220=>"011110110",
77221=>"111111110",
77222=>"010010010",
77223=>"011100100",
77224=>"001011111",
77225=>"111111111",
77226=>"100100100",
77227=>"100100100",
77228=>"000000111",
77229=>"100000000",
77230=>"000101010",
77231=>"001001011",
77232=>"100100110",
77233=>"111100100",
77234=>"101110000",
77235=>"110110011",
77236=>"001001001",
77237=>"110111111",
77238=>"110110110",
77239=>"001000000",
77240=>"110100110",
77241=>"111100100",
77242=>"100110100",
77243=>"011111111",
77244=>"111111111",
77245=>"011001000",
77246=>"110110110",
77247=>"011001001",
77248=>"101110101",
77249=>"110010000",
77250=>"100110001",
77251=>"100000101",
77252=>"100100110",
77253=>"000101100",
77254=>"110010000",
77255=>"111111110",
77256=>"011011110",
77257=>"011001000",
77258=>"010000100",
77259=>"011011001",
77260=>"000011001",
77261=>"001010100",
77262=>"011011001",
77263=>"100101111",
77264=>"000011000",
77265=>"000000010",
77266=>"111110010",
77267=>"110100100",
77268=>"110000100",
77269=>"111110110",
77270=>"111100100",
77271=>"000100100",
77272=>"001001001",
77273=>"000000010",
77274=>"110110110",
77275=>"011011011",
77276=>"001110000",
77277=>"111011111",
77278=>"100100011",
77279=>"110110100",
77280=>"011111011",
77281=>"101111110",
77282=>"011011011",
77283=>"110111110",
77284=>"000001010",
77285=>"111101100",
77286=>"001110100",
77287=>"001010111",
77288=>"000110100",
77289=>"001000111",
77290=>"100001001",
77291=>"111100000",
77292=>"111100100",
77293=>"100000000",
77294=>"000000000",
77295=>"100000111",
77296=>"010111111",
77297=>"000100100",
77298=>"000110000",
77299=>"011011010",
77300=>"011100100",
77301=>"000001011",
77302=>"000100010",
77303=>"001011011",
77304=>"110100111",
77305=>"011011111",
77306=>"010010110",
77307=>"000000000",
77308=>"011101111",
77309=>"001011110",
77310=>"000000010",
77311=>"000000000",
77312=>"000000100",
77313=>"000000000",
77314=>"101101101",
77315=>"111000111",
77316=>"111011110",
77317=>"101111000",
77318=>"100100010",
77319=>"111110111",
77320=>"111101101",
77321=>"010000000",
77322=>"011011000",
77323=>"101101100",
77324=>"000100000",
77325=>"111000000",
77326=>"001111110",
77327=>"010111100",
77328=>"111011001",
77329=>"100101101",
77330=>"000000011",
77331=>"000000000",
77332=>"000000000",
77333=>"011111000",
77334=>"110101111",
77335=>"001011111",
77336=>"000000111",
77337=>"011111111",
77338=>"100000101",
77339=>"111001101",
77340=>"010111000",
77341=>"010000000",
77342=>"111000001",
77343=>"011111000",
77344=>"010101111",
77345=>"111000111",
77346=>"011011111",
77347=>"010010000",
77348=>"111111010",
77349=>"000100000",
77350=>"111111111",
77351=>"100110000",
77352=>"000001101",
77353=>"101100111",
77354=>"001111000",
77355=>"011000001",
77356=>"110010011",
77357=>"010011101",
77358=>"111111011",
77359=>"000010100",
77360=>"100000000",
77361=>"110011001",
77362=>"001000111",
77363=>"111110111",
77364=>"110000000",
77365=>"111111111",
77366=>"110110100",
77367=>"010001111",
77368=>"000100000",
77369=>"101000000",
77370=>"000000000",
77371=>"111111111",
77372=>"111111110",
77373=>"001011011",
77374=>"101000000",
77375=>"101111011",
77376=>"111001011",
77377=>"111110010",
77378=>"000000000",
77379=>"110111110",
77380=>"011001000",
77381=>"000010010",
77382=>"000111100",
77383=>"101100110",
77384=>"101110010",
77385=>"000000001",
77386=>"100100111",
77387=>"110000111",
77388=>"111000111",
77389=>"001001000",
77390=>"111110111",
77391=>"010101111",
77392=>"110111111",
77393=>"000100111",
77394=>"111111111",
77395=>"110010010",
77396=>"101111100",
77397=>"110100111",
77398=>"111110111",
77399=>"111101101",
77400=>"000000001",
77401=>"111111111",
77402=>"011111110",
77403=>"111111010",
77404=>"011100111",
77405=>"001011000",
77406=>"000100101",
77407=>"111111011",
77408=>"111111000",
77409=>"111111111",
77410=>"101000111",
77411=>"110111000",
77412=>"111111100",
77413=>"010010010",
77414=>"001000010",
77415=>"000000000",
77416=>"000011000",
77417=>"000000000",
77418=>"000000000",
77419=>"110111000",
77420=>"011111111",
77421=>"000111000",
77422=>"011111111",
77423=>"010111010",
77424=>"110111111",
77425=>"000000000",
77426=>"111111001",
77427=>"000110000",
77428=>"111100000",
77429=>"000101000",
77430=>"000000011",
77431=>"101000000",
77432=>"111101000",
77433=>"010011111",
77434=>"000100001",
77435=>"001001001",
77436=>"001000111",
77437=>"100100000",
77438=>"000001001",
77439=>"110111000",
77440=>"111010010",
77441=>"100000000",
77442=>"111000111",
77443=>"111000101",
77444=>"011111111",
77445=>"000000010",
77446=>"011011000",
77447=>"010110110",
77448=>"111111111",
77449=>"111111100",
77450=>"000111011",
77451=>"110010111",
77452=>"111101001",
77453=>"100111111",
77454=>"000110111",
77455=>"110110000",
77456=>"000011110",
77457=>"111111010",
77458=>"100111111",
77459=>"001001011",
77460=>"111011111",
77461=>"111111111",
77462=>"101111000",
77463=>"111000001",
77464=>"000000000",
77465=>"000100111",
77466=>"111011111",
77467=>"100111000",
77468=>"010101111",
77469=>"110100111",
77470=>"000000000",
77471=>"111001111",
77472=>"000010001",
77473=>"111000111",
77474=>"100001000",
77475=>"000000111",
77476=>"000000010",
77477=>"111111110",
77478=>"000001011",
77479=>"000000000",
77480=>"111101111",
77481=>"111100111",
77482=>"000000000",
77483=>"101101101",
77484=>"001010110",
77485=>"111111111",
77486=>"000111011",
77487=>"011111110",
77488=>"100101111",
77489=>"000101010",
77490=>"111101111",
77491=>"001001111",
77492=>"000010000",
77493=>"000011000",
77494=>"010000100",
77495=>"011000110",
77496=>"100110110",
77497=>"011010111",
77498=>"000000111",
77499=>"111000111",
77500=>"101100111",
77501=>"111000000",
77502=>"010111100",
77503=>"000000101",
77504=>"011111000",
77505=>"010000111",
77506=>"100101000",
77507=>"111111010",
77508=>"101111111",
77509=>"000101101",
77510=>"100101111",
77511=>"111111111",
77512=>"110110000",
77513=>"111111111",
77514=>"011010101",
77515=>"010111110",
77516=>"010111011",
77517=>"000000111",
77518=>"100101100",
77519=>"111111111",
77520=>"111111000",
77521=>"001111100",
77522=>"111111111",
77523=>"101011111",
77524=>"000000000",
77525=>"000110000",
77526=>"101001000",
77527=>"100101010",
77528=>"111111011",
77529=>"110001000",
77530=>"000000010",
77531=>"101000101",
77532=>"111101011",
77533=>"000111111",
77534=>"111110111",
77535=>"011100010",
77536=>"010011111",
77537=>"001000111",
77538=>"110111111",
77539=>"011111011",
77540=>"011111001",
77541=>"111011101",
77542=>"110111000",
77543=>"111111101",
77544=>"101100000",
77545=>"000000100",
77546=>"001011100",
77547=>"111001111",
77548=>"101001001",
77549=>"110101111",
77550=>"000000111",
77551=>"000100011",
77552=>"111100000",
77553=>"010011111",
77554=>"111111111",
77555=>"110111000",
77556=>"110100011",
77557=>"010110111",
77558=>"111000000",
77559=>"111001111",
77560=>"111111111",
77561=>"111011000",
77562=>"011010111",
77563=>"101110000",
77564=>"111111101",
77565=>"010110111",
77566=>"110110000",
77567=>"001111110",
77568=>"011011001",
77569=>"000100111",
77570=>"101000000",
77571=>"000101110",
77572=>"100111001",
77573=>"111110010",
77574=>"100111111",
77575=>"010000000",
77576=>"000110100",
77577=>"110010110",
77578=>"011111011",
77579=>"000000011",
77580=>"101100000",
77581=>"011101111",
77582=>"111111111",
77583=>"000001001",
77584=>"110110111",
77585=>"110111110",
77586=>"111111000",
77587=>"011011111",
77588=>"101000000",
77589=>"011111010",
77590=>"011001000",
77591=>"000000111",
77592=>"111111100",
77593=>"111111101",
77594=>"000111000",
77595=>"000000010",
77596=>"101000111",
77597=>"000000100",
77598=>"111111000",
77599=>"110010010",
77600=>"010010000",
77601=>"010011011",
77602=>"011000111",
77603=>"000000000",
77604=>"100101111",
77605=>"111101001",
77606=>"000011011",
77607=>"000011010",
77608=>"101000100",
77609=>"001000100",
77610=>"001111111",
77611=>"111100100",
77612=>"000100001",
77613=>"000001010",
77614=>"011111001",
77615=>"110111111",
77616=>"000110000",
77617=>"111001000",
77618=>"001000011",
77619=>"111110111",
77620=>"111111101",
77621=>"111111010",
77622=>"111100110",
77623=>"000011111",
77624=>"111111000",
77625=>"111111111",
77626=>"000000100",
77627=>"100011000",
77628=>"111111001",
77629=>"001101111",
77630=>"010000100",
77631=>"111111111",
77632=>"111101101",
77633=>"000110110",
77634=>"111100000",
77635=>"011011110",
77636=>"000110110",
77637=>"111001001",
77638=>"010110000",
77639=>"000110101",
77640=>"000000000",
77641=>"110111111",
77642=>"111101110",
77643=>"001110111",
77644=>"111111111",
77645=>"000111111",
77646=>"011101110",
77647=>"000000000",
77648=>"111110111",
77649=>"011011111",
77650=>"010111100",
77651=>"011001000",
77652=>"000000000",
77653=>"111111100",
77654=>"001001001",
77655=>"111111111",
77656=>"000100101",
77657=>"001111111",
77658=>"111111101",
77659=>"111111111",
77660=>"010111110",
77661=>"000001001",
77662=>"000000000",
77663=>"111110110",
77664=>"000010010",
77665=>"001111000",
77666=>"110000000",
77667=>"110100000",
77668=>"111111111",
77669=>"111001000",
77670=>"000100101",
77671=>"110111111",
77672=>"111111010",
77673=>"000111111",
77674=>"000010110",
77675=>"000000101",
77676=>"010100010",
77677=>"010110111",
77678=>"010011000",
77679=>"010010111",
77680=>"010110110",
77681=>"000001000",
77682=>"111011011",
77683=>"000110111",
77684=>"110000111",
77685=>"000000001",
77686=>"101111111",
77687=>"111111000",
77688=>"000000000",
77689=>"101010110",
77690=>"010111111",
77691=>"001001001",
77692=>"000110111",
77693=>"110100000",
77694=>"000101000",
77695=>"111111111",
77696=>"110111000",
77697=>"111101111",
77698=>"010111111",
77699=>"000100111",
77700=>"010111111",
77701=>"101110101",
77702=>"111101101",
77703=>"011111111",
77704=>"111111001",
77705=>"100000010",
77706=>"000000011",
77707=>"000000000",
77708=>"000000000",
77709=>"110111111",
77710=>"111111010",
77711=>"101001111",
77712=>"100001011",
77713=>"110010001",
77714=>"111111101",
77715=>"000000001",
77716=>"111011001",
77717=>"111111110",
77718=>"011110011",
77719=>"101101011",
77720=>"000110111",
77721=>"000000001",
77722=>"010111111",
77723=>"000000000",
77724=>"111011001",
77725=>"110110010",
77726=>"000000111",
77727=>"000000000",
77728=>"001001001",
77729=>"111111000",
77730=>"001101100",
77731=>"010000101",
77732=>"110110000",
77733=>"100110100",
77734=>"001111111",
77735=>"010001010",
77736=>"010111111",
77737=>"111111111",
77738=>"000000000",
77739=>"111101110",
77740=>"001001000",
77741=>"111111111",
77742=>"111100000",
77743=>"001000010",
77744=>"000001010",
77745=>"000110110",
77746=>"010001000",
77747=>"000100110",
77748=>"000110111",
77749=>"010111000",
77750=>"111111111",
77751=>"101111011",
77752=>"011110001",
77753=>"010111100",
77754=>"111110110",
77755=>"010110110",
77756=>"001000100",
77757=>"111111111",
77758=>"010010001",
77759=>"111111000",
77760=>"010111000",
77761=>"010111110",
77762=>"110111111",
77763=>"001101111",
77764=>"000000000",
77765=>"100100100",
77766=>"111111101",
77767=>"010111111",
77768=>"000000101",
77769=>"111111000",
77770=>"111111111",
77771=>"000111010",
77772=>"000011011",
77773=>"000010111",
77774=>"001010110",
77775=>"000010111",
77776=>"010010110",
77777=>"001101100",
77778=>"111001000",
77779=>"000110001",
77780=>"111001111",
77781=>"011100100",
77782=>"110000111",
77783=>"110111111",
77784=>"000000000",
77785=>"110110000",
77786=>"111100100",
77787=>"110000010",
77788=>"111101000",
77789=>"000011111",
77790=>"000111111",
77791=>"111110110",
77792=>"010000000",
77793=>"110000000",
77794=>"101100001",
77795=>"000100100",
77796=>"000010111",
77797=>"010100010",
77798=>"000000111",
77799=>"010001100",
77800=>"110100101",
77801=>"000110100",
77802=>"101110111",
77803=>"000111110",
77804=>"111000000",
77805=>"101010110",
77806=>"011001001",
77807=>"010000101",
77808=>"000000000",
77809=>"011011001",
77810=>"000010010",
77811=>"010011011",
77812=>"111111100",
77813=>"101001000",
77814=>"111111110",
77815=>"000110011",
77816=>"111000000",
77817=>"111000010",
77818=>"011111111",
77819=>"111111111",
77820=>"010111111",
77821=>"000110101",
77822=>"001101111",
77823=>"000000111",
77824=>"011011000",
77825=>"001011011",
77826=>"100100100",
77827=>"100100001",
77828=>"110110110",
77829=>"000100100",
77830=>"101100100",
77831=>"000000000",
77832=>"000000000",
77833=>"100000110",
77834=>"001010010",
77835=>"100100100",
77836=>"000000100",
77837=>"100011111",
77838=>"111100110",
77839=>"011100111",
77840=>"111101111",
77841=>"111100110",
77842=>"100100110",
77843=>"001011011",
77844=>"111111101",
77845=>"111100000",
77846=>"000101001",
77847=>"100010110",
77848=>"100100100",
77849=>"101011011",
77850=>"111011111",
77851=>"000001111",
77852=>"011011001",
77853=>"011011000",
77854=>"111100100",
77855=>"000011011",
77856=>"011011001",
77857=>"100000100",
77858=>"000111110",
77859=>"011011000",
77860=>"100010100",
77861=>"001011011",
77862=>"000011011",
77863=>"000000000",
77864=>"110011011",
77865=>"000011111",
77866=>"100000000",
77867=>"011000000",
77868=>"010011011",
77869=>"111110111",
77870=>"110111100",
77871=>"110000000",
77872=>"010011000",
77873=>"111101000",
77874=>"010000000",
77875=>"011011001",
77876=>"000011011",
77877=>"001000111",
77878=>"001011011",
77879=>"000000000",
77880=>"111100011",
77881=>"111100000",
77882=>"010000000",
77883=>"010010011",
77884=>"010010010",
77885=>"111011110",
77886=>"001100000",
77887=>"100111101",
77888=>"111111010",
77889=>"001001000",
77890=>"011100100",
77891=>"111000000",
77892=>"011101101",
77893=>"000100100",
77894=>"011111111",
77895=>"000011011",
77896=>"001111101",
77897=>"111100111",
77898=>"111100100",
77899=>"011110111",
77900=>"000000000",
77901=>"100000000",
77902=>"011110111",
77903=>"010011011",
77904=>"101000100",
77905=>"111111111",
77906=>"001000000",
77907=>"011101000",
77908=>"000000001",
77909=>"011011010",
77910=>"000001000",
77911=>"111000100",
77912=>"011110111",
77913=>"011011001",
77914=>"000101001",
77915=>"100101111",
77916=>"010100000",
77917=>"111101100",
77918=>"111011010",
77919=>"110100100",
77920=>"011001000",
77921=>"010000000",
77922=>"111100100",
77923=>"000110010",
77924=>"100000100",
77925=>"111111111",
77926=>"000111111",
77927=>"100011011",
77928=>"100010101",
77929=>"011000100",
77930=>"100111011",
77931=>"000011000",
77932=>"000101010",
77933=>"111101001",
77934=>"111100101",
77935=>"000101111",
77936=>"110011111",
77937=>"111000000",
77938=>"110100000",
77939=>"000100000",
77940=>"000101011",
77941=>"100100001",
77942=>"100000000",
77943=>"000100000",
77944=>"011011000",
77945=>"100110011",
77946=>"100000011",
77947=>"000000000",
77948=>"010110011",
77949=>"010110000",
77950=>"010000101",
77951=>"100100100",
77952=>"011011000",
77953=>"101100110",
77954=>"100000000",
77955=>"000111110",
77956=>"100000100",
77957=>"011011111",
77958=>"110011000",
77959=>"000001001",
77960=>"001101101",
77961=>"111100000",
77962=>"111100100",
77963=>"100000000",
77964=>"100100001",
77965=>"000000100",
77966=>"111100000",
77967=>"001000000",
77968=>"100101101",
77969=>"000000011",
77970=>"000011001",
77971=>"000101101",
77972=>"000011011",
77973=>"111100101",
77974=>"111011000",
77975=>"110100000",
77976=>"000000000",
77977=>"011011111",
77978=>"010011011",
77979=>"100000000",
77980=>"011010100",
77981=>"100000000",
77982=>"111100000",
77983=>"111100100",
77984=>"011011000",
77985=>"111000011",
77986=>"110011000",
77987=>"000010111",
77988=>"101100000",
77989=>"100110000",
77990=>"000111011",
77991=>"100111010",
77992=>"111000000",
77993=>"100100101",
77994=>"111100101",
77995=>"111100100",
77996=>"000010010",
77997=>"000000100",
77998=>"011110010",
77999=>"100101111",
78000=>"101000000",
78001=>"111110110",
78002=>"011100100",
78003=>"001110110",
78004=>"000011111",
78005=>"000010001",
78006=>"000101100",
78007=>"000000001",
78008=>"000001001",
78009=>"010001001",
78010=>"000011111",
78011=>"011111111",
78012=>"001011110",
78013=>"111111100",
78014=>"000000000",
78015=>"000000000",
78016=>"110000100",
78017=>"100100100",
78018=>"111111000",
78019=>"111000111",
78020=>"000000100",
78021=>"011011100",
78022=>"011011110",
78023=>"111111111",
78024=>"000100100",
78025=>"000000011",
78026=>"110101100",
78027=>"000000000",
78028=>"000011011",
78029=>"100001000",
78030=>"000111001",
78031=>"100000010",
78032=>"000000011",
78033=>"001111101",
78034=>"100001011",
78035=>"111100111",
78036=>"100000101",
78037=>"000100000",
78038=>"100100000",
78039=>"100100011",
78040=>"010011000",
78041=>"000100011",
78042=>"000111110",
78043=>"100100100",
78044=>"001011110",
78045=>"100100111",
78046=>"101110111",
78047=>"000000011",
78048=>"111000000",
78049=>"111100100",
78050=>"011000100",
78051=>"011000011",
78052=>"111100001",
78053=>"100100100",
78054=>"101000011",
78055=>"000011011",
78056=>"111100101",
78057=>"010011011",
78058=>"110101101",
78059=>"011100110",
78060=>"111100100",
78061=>"001000001",
78062=>"111100001",
78063=>"110100110",
78064=>"011011011",
78065=>"111111000",
78066=>"000100000",
78067=>"010111000",
78068=>"000100000",
78069=>"101100100",
78070=>"100000011",
78071=>"000001011",
78072=>"010110010",
78073=>"100101111",
78074=>"000011000",
78075=>"101111101",
78076=>"111011000",
78077=>"110100100",
78078=>"001011011",
78079=>"111100100",
78080=>"011001000",
78081=>"100110110",
78082=>"000000000",
78083=>"000111101",
78084=>"100000101",
78085=>"000000101",
78086=>"000000100",
78087=>"110000111",
78088=>"101100001",
78089=>"000000000",
78090=>"100000101",
78091=>"100110000",
78092=>"110110000",
78093=>"010011111",
78094=>"010011101",
78095=>"101111111",
78096=>"111111000",
78097=>"100000001",
78098=>"001101001",
78099=>"101111111",
78100=>"111001000",
78101=>"101111010",
78102=>"111101010",
78103=>"111110111",
78104=>"000001101",
78105=>"111111001",
78106=>"000000101",
78107=>"000000111",
78108=>"101101111",
78109=>"000111111",
78110=>"111000000",
78111=>"000110111",
78112=>"000000001",
78113=>"011111000",
78114=>"000110010",
78115=>"100110000",
78116=>"000001000",
78117=>"111001001",
78118=>"001111111",
78119=>"000000000",
78120=>"111111010",
78121=>"011110001",
78122=>"111101101",
78123=>"101001111",
78124=>"111111100",
78125=>"000101111",
78126=>"000000100",
78127=>"010000100",
78128=>"000001101",
78129=>"101001001",
78130=>"000000000",
78131=>"101001001",
78132=>"000110101",
78133=>"110000000",
78134=>"011111110",
78135=>"000000001",
78136=>"111001000",
78137=>"000000111",
78138=>"101100101",
78139=>"000001110",
78140=>"100100100",
78141=>"110111101",
78142=>"000100111",
78143=>"011001010",
78144=>"101101001",
78145=>"111001001",
78146=>"000010000",
78147=>"100110101",
78148=>"011000001",
78149=>"000001000",
78150=>"111111101",
78151=>"111111111",
78152=>"110110011",
78153=>"111110001",
78154=>"000000111",
78155=>"010101000",
78156=>"000000111",
78157=>"001101110",
78158=>"011001000",
78159=>"101010111",
78160=>"010010110",
78161=>"111000000",
78162=>"111111110",
78163=>"001001011",
78164=>"010010000",
78165=>"100010011",
78166=>"000000100",
78167=>"110001001",
78168=>"000000000",
78169=>"100100000",
78170=>"000110111",
78171=>"101100001",
78172=>"101000101",
78173=>"000001011",
78174=>"111011000",
78175=>"010000000",
78176=>"010110111",
78177=>"010000100",
78178=>"010010000",
78179=>"100001111",
78180=>"100101001",
78181=>"011001101",
78182=>"111001000",
78183=>"001111111",
78184=>"000000000",
78185=>"101000000",
78186=>"111110111",
78187=>"111101000",
78188=>"001000000",
78189=>"010011111",
78190=>"000000101",
78191=>"110000001",
78192=>"110110101",
78193=>"111001000",
78194=>"111111010",
78195=>"001001111",
78196=>"100000000",
78197=>"000001001",
78198=>"000100111",
78199=>"111110000",
78200=>"011001000",
78201=>"010000111",
78202=>"000001111",
78203=>"111000010",
78204=>"100110110",
78205=>"100000100",
78206=>"010111010",
78207=>"000000010",
78208=>"001000000",
78209=>"111000000",
78210=>"111111000",
78211=>"001111000",
78212=>"111110000",
78213=>"001000111",
78214=>"110001000",
78215=>"000000100",
78216=>"011011011",
78217=>"010010000",
78218=>"000001111",
78219=>"100001000",
78220=>"010110000",
78221=>"101010000",
78222=>"111111101",
78223=>"000000001",
78224=>"110110111",
78225=>"011111011",
78226=>"101101101",
78227=>"101100000",
78228=>"001111101",
78229=>"000000000",
78230=>"111101000",
78231=>"000011110",
78232=>"111111001",
78233=>"000110110",
78234=>"011111001",
78235=>"000010000",
78236=>"001111010",
78237=>"010000001",
78238=>"000100111",
78239=>"000000101",
78240=>"000100110",
78241=>"100000000",
78242=>"010101111",
78243=>"111000000",
78244=>"010000011",
78245=>"001001010",
78246=>"011110100",
78247=>"000101111",
78248=>"000111111",
78249=>"000110110",
78250=>"000110011",
78251=>"010000000",
78252=>"111010000",
78253=>"000000111",
78254=>"100100101",
78255=>"110110111",
78256=>"000000010",
78257=>"010011001",
78258=>"111000000",
78259=>"000100110",
78260=>"111111011",
78261=>"111000000",
78262=>"111111011",
78263=>"111111000",
78264=>"001001001",
78265=>"000010010",
78266=>"111111111",
78267=>"111100111",
78268=>"000000100",
78269=>"110110111",
78270=>"011000000",
78271=>"110110000",
78272=>"001011000",
78273=>"001000111",
78274=>"101111111",
78275=>"101001010",
78276=>"011011001",
78277=>"000001101",
78278=>"000000011",
78279=>"111100110",
78280=>"111101000",
78281=>"010110110",
78282=>"101111000",
78283=>"111000000",
78284=>"000000111",
78285=>"001011111",
78286=>"000000111",
78287=>"000000111",
78288=>"000000000",
78289=>"011000011",
78290=>"101000011",
78291=>"000000101",
78292=>"110110000",
78293=>"110100111",
78294=>"001000111",
78295=>"110000111",
78296=>"111111010",
78297=>"000101001",
78298=>"111010001",
78299=>"000010000",
78300=>"101100111",
78301=>"101111000",
78302=>"111110000",
78303=>"111111000",
78304=>"000000100",
78305=>"000000101",
78306=>"111110010",
78307=>"000111011",
78308=>"101001111",
78309=>"000010000",
78310=>"000000101",
78311=>"001000000",
78312=>"000000000",
78313=>"000010111",
78314=>"001000101",
78315=>"111111110",
78316=>"000010111",
78317=>"000001001",
78318=>"000000000",
78319=>"111000000",
78320=>"100100011",
78321=>"000011111",
78322=>"011000101",
78323=>"111000100",
78324=>"100110101",
78325=>"000000010",
78326=>"000001000",
78327=>"001000101",
78328=>"111111000",
78329=>"110000010",
78330=>"101000110",
78331=>"001011001",
78332=>"111101000",
78333=>"111010001",
78334=>"100100111",
78335=>"111111001",
78336=>"111011000",
78337=>"110011111",
78338=>"100000000",
78339=>"000000111",
78340=>"001011011",
78341=>"000001001",
78342=>"000010000",
78343=>"011011111",
78344=>"001011110",
78345=>"011010000",
78346=>"011011000",
78347=>"000100111",
78348=>"000000111",
78349=>"000000101",
78350=>"100011001",
78351=>"000001111",
78352=>"011010000",
78353=>"011111000",
78354=>"101111100",
78355=>"000111101",
78356=>"111011000",
78357=>"111110000",
78358=>"010011001",
78359=>"111111010",
78360=>"010010110",
78361=>"111111111",
78362=>"111011000",
78363=>"011010000",
78364=>"100100101",
78365=>"111010000",
78366=>"000011011",
78367=>"000000010",
78368=>"000000101",
78369=>"011000111",
78370=>"111011010",
78371=>"111011011",
78372=>"001001000",
78373=>"000110001",
78374=>"110010000",
78375=>"111000000",
78376=>"111011000",
78377=>"011000001",
78378=>"011000000",
78379=>"000000010",
78380=>"110100000",
78381=>"111011011",
78382=>"111011000",
78383=>"010000000",
78384=>"000111111",
78385=>"001001001",
78386=>"111111011",
78387=>"000010111",
78388=>"111011000",
78389=>"111111111",
78390=>"010011100",
78391=>"000110000",
78392=>"011111110",
78393=>"001101111",
78394=>"000100101",
78395=>"100000000",
78396=>"000100101",
78397=>"111111010",
78398=>"000000000",
78399=>"111111000",
78400=>"001000111",
78401=>"010011000",
78402=>"000010000",
78403=>"111111010",
78404=>"101100101",
78405=>"010000100",
78406=>"000000101",
78407=>"000000100",
78408=>"001111111",
78409=>"010111000",
78410=>"010000101",
78411=>"000000101",
78412=>"111111000",
78413=>"100100110",
78414=>"100100100",
78415=>"001000101",
78416=>"101011011",
78417=>"000111010",
78418=>"000010011",
78419=>"011111000",
78420=>"000011010",
78421=>"110110011",
78422=>"000100110",
78423=>"011111000",
78424=>"111001010",
78425=>"111001001",
78426=>"100100000",
78427=>"000000000",
78428=>"010011000",
78429=>"001001001",
78430=>"010000011",
78431=>"111001000",
78432=>"100010000",
78433=>"111111000",
78434=>"100000100",
78435=>"100100110",
78436=>"000100001",
78437=>"111010100",
78438=>"111010000",
78439=>"011111000",
78440=>"000011111",
78441=>"000010011",
78442=>"000000000",
78443=>"000000111",
78444=>"100111110",
78445=>"111111010",
78446=>"101100100",
78447=>"111101111",
78448=>"000001101",
78449=>"000000010",
78450=>"011010000",
78451=>"010000000",
78452=>"010000000",
78453=>"000000111",
78454=>"111111101",
78455=>"000000000",
78456=>"111001010",
78457=>"000100111",
78458=>"010000000",
78459=>"100101100",
78460=>"110000000",
78461=>"111100000",
78462=>"111110000",
78463=>"111111001",
78464=>"011010000",
78465=>"000111111",
78466=>"010010000",
78467=>"111001011",
78468=>"001010010",
78469=>"000000100",
78470=>"000010100",
78471=>"000001001",
78472=>"101111111",
78473=>"100101010",
78474=>"011001100",
78475=>"000010000",
78476=>"111011000",
78477=>"101100101",
78478=>"010011000",
78479=>"000000001",
78480=>"011011000",
78481=>"000111001",
78482=>"010010000",
78483=>"000000011",
78484=>"100000011",
78485=>"011011000",
78486=>"000000001",
78487=>"011001100",
78488=>"000000000",
78489=>"000000111",
78490=>"000000000",
78491=>"000000110",
78492=>"111110000",
78493=>"101000100",
78494=>"011000000",
78495=>"010010000",
78496=>"111111001",
78497=>"010111010",
78498=>"010011000",
78499=>"000111111",
78500=>"001101111",
78501=>"111101100",
78502=>"111110000",
78503=>"001111010",
78504=>"010010010",
78505=>"001111111",
78506=>"000100100",
78507=>"111010000",
78508=>"011010111",
78509=>"111010000",
78510=>"100111000",
78511=>"000100111",
78512=>"001010100",
78513=>"001111111",
78514=>"000000110",
78515=>"110100010",
78516=>"111110011",
78517=>"010111000",
78518=>"111011001",
78519=>"100000101",
78520=>"100100100",
78521=>"100000010",
78522=>"000000100",
78523=>"001111001",
78524=>"000000000",
78525=>"100111111",
78526=>"110011001",
78527=>"011010000",
78528=>"111000001",
78529=>"101101011",
78530=>"010110011",
78531=>"101100100",
78532=>"100101000",
78533=>"100000001",
78534=>"000001011",
78535=>"111000100",
78536=>"111111111",
78537=>"010011010",
78538=>"000000000",
78539=>"100000101",
78540=>"000011000",
78541=>"011110100",
78542=>"000000000",
78543=>"010010000",
78544=>"000000000",
78545=>"111100100",
78546=>"000100111",
78547=>"111111011",
78548=>"100101111",
78549=>"100111110",
78550=>"000000000",
78551=>"100111111",
78552=>"000011010",
78553=>"010011111",
78554=>"010000100",
78555=>"000000000",
78556=>"000111101",
78557=>"000111111",
78558=>"111101111",
78559=>"000000111",
78560=>"111111010",
78561=>"000100110",
78562=>"111100010",
78563=>"111110000",
78564=>"000000000",
78565=>"000000110",
78566=>"010000111",
78567=>"100100111",
78568=>"000111111",
78569=>"011011111",
78570=>"110011001",
78571=>"111101011",
78572=>"011111010",
78573=>"100000011",
78574=>"000110000",
78575=>"110000000",
78576=>"000000010",
78577=>"001000101",
78578=>"001001010",
78579=>"011011000",
78580=>"111110001",
78581=>"110001010",
78582=>"000000000",
78583=>"000011111",
78584=>"000000010",
78585=>"001111111",
78586=>"111101111",
78587=>"011111111",
78588=>"000000101",
78589=>"000100000",
78590=>"100111111",
78591=>"000000000",
78592=>"100000000",
78593=>"000100000",
78594=>"110000000",
78595=>"000000111",
78596=>"000001011",
78597=>"110000001",
78598=>"111101010",
78599=>"111000001",
78600=>"000101101",
78601=>"010110000",
78602=>"111111010",
78603=>"000110000",
78604=>"000111101",
78605=>"000010000",
78606=>"111011010",
78607=>"000111111",
78608=>"000010110",
78609=>"000111111",
78610=>"000000000",
78611=>"110111111",
78612=>"101000010",
78613=>"001111111",
78614=>"011100000",
78615=>"000111111",
78616=>"001001000",
78617=>"000100111",
78618=>"000000111",
78619=>"001000000",
78620=>"000111111",
78621=>"000100000",
78622=>"111110000",
78623=>"101000000",
78624=>"001100001",
78625=>"000000000",
78626=>"111010010",
78627=>"000000111",
78628=>"111000001",
78629=>"000000001",
78630=>"000000111",
78631=>"111111111",
78632=>"000111010",
78633=>"000000000",
78634=>"111011111",
78635=>"000111000",
78636=>"111011111",
78637=>"000111111",
78638=>"101001001",
78639=>"000001110",
78640=>"000101111",
78641=>"010000001",
78642=>"000000101",
78643=>"110011111",
78644=>"001000000",
78645=>"000110101",
78646=>"100111011",
78647=>"111000100",
78648=>"110000000",
78649=>"111000100",
78650=>"001101011",
78651=>"001000000",
78652=>"000010011",
78653=>"011001010",
78654=>"110100000",
78655=>"111110000",
78656=>"000000111",
78657=>"111010000",
78658=>"111111101",
78659=>"011100110",
78660=>"111111001",
78661=>"001111101",
78662=>"100000000",
78663=>"011000000",
78664=>"100111100",
78665=>"110111000",
78666=>"111111010",
78667=>"111010000",
78668=>"010000000",
78669=>"010010110",
78670=>"111101100",
78671=>"110110111",
78672=>"111000000",
78673=>"101000000",
78674=>"011111111",
78675=>"011000000",
78676=>"000000010",
78677=>"011000000",
78678=>"111011000",
78679=>"111111110",
78680=>"111111011",
78681=>"010011001",
78682=>"111110000",
78683=>"111010001",
78684=>"000000000",
78685=>"111100000",
78686=>"001111111",
78687=>"100001111",
78688=>"101111101",
78689=>"111110000",
78690=>"000000000",
78691=>"011101000",
78692=>"010000000",
78693=>"110000000",
78694=>"000001111",
78695=>"111101111",
78696=>"111101000",
78697=>"101110111",
78698=>"011000000",
78699=>"001001001",
78700=>"000000000",
78701=>"111111111",
78702=>"010111011",
78703=>"111111100",
78704=>"101000001",
78705=>"000000111",
78706=>"001111111",
78707=>"000000111",
78708=>"100111010",
78709=>"000000100",
78710=>"111111000",
78711=>"000001000",
78712=>"000101100",
78713=>"110010111",
78714=>"111110011",
78715=>"000000100",
78716=>"111111100",
78717=>"100000001",
78718=>"001111010",
78719=>"111000000",
78720=>"010011000",
78721=>"010010000",
78722=>"000000111",
78723=>"000111000",
78724=>"000000111",
78725=>"111000000",
78726=>"000000100",
78727=>"110000100",
78728=>"110111010",
78729=>"111100111",
78730=>"111011111",
78731=>"000000100",
78732=>"111101000",
78733=>"101101111",
78734=>"111000000",
78735=>"000010000",
78736=>"101101011",
78737=>"010011000",
78738=>"111010010",
78739=>"001100000",
78740=>"000000010",
78741=>"001011000",
78742=>"111110101",
78743=>"000000001",
78744=>"001101111",
78745=>"101000110",
78746=>"000000111",
78747=>"010000000",
78748=>"111010001",
78749=>"000000000",
78750=>"000000110",
78751=>"111000000",
78752=>"011001101",
78753=>"010111000",
78754=>"000101111",
78755=>"111000000",
78756=>"001111100",
78757=>"111110110",
78758=>"111001001",
78759=>"110010111",
78760=>"010111111",
78761=>"010000000",
78762=>"000000000",
78763=>"111001000",
78764=>"000110010",
78765=>"111000000",
78766=>"010100000",
78767=>"111110101",
78768=>"000110111",
78769=>"111110001",
78770=>"010000101",
78771=>"011011100",
78772=>"100110111",
78773=>"001111101",
78774=>"000111111",
78775=>"000101101",
78776=>"100000110",
78777=>"110000100",
78778=>"000000110",
78779=>"001111110",
78780=>"000001111",
78781=>"111111111",
78782=>"001011010",
78783=>"101000111",
78784=>"110000011",
78785=>"111000000",
78786=>"000111111",
78787=>"011001000",
78788=>"001000100",
78789=>"101000000",
78790=>"100111111",
78791=>"101001000",
78792=>"110000000",
78793=>"000111010",
78794=>"000110010",
78795=>"000000111",
78796=>"000111000",
78797=>"001001110",
78798=>"111001000",
78799=>"000000110",
78800=>"000011111",
78801=>"110000001",
78802=>"111000110",
78803=>"000110111",
78804=>"101000000",
78805=>"111000000",
78806=>"000000000",
78807=>"000000000",
78808=>"000111111",
78809=>"000111110",
78810=>"010100000",
78811=>"111111000",
78812=>"000010001",
78813=>"100111111",
78814=>"100110010",
78815=>"000000101",
78816=>"010111000",
78817=>"111000000",
78818=>"001000100",
78819=>"111000000",
78820=>"011000000",
78821=>"110000000",
78822=>"010000000",
78823=>"110000100",
78824=>"000010110",
78825=>"001111100",
78826=>"111110010",
78827=>"000111111",
78828=>"000111111",
78829=>"000100111",
78830=>"111000000",
78831=>"000000100",
78832=>"000010010",
78833=>"111110010",
78834=>"001011000",
78835=>"111111000",
78836=>"011010000",
78837=>"111101000",
78838=>"010000011",
78839=>"011100110",
78840=>"000000001",
78841=>"001111111",
78842=>"000000111",
78843=>"111000000",
78844=>"010010001",
78845=>"000000000",
78846=>"111101111",
78847=>"000101101",
78848=>"100100111",
78849=>"111100110",
78850=>"010111111",
78851=>"111000000",
78852=>"110011111",
78853=>"100001000",
78854=>"100111111",
78855=>"000000010",
78856=>"000011011",
78857=>"000111000",
78858=>"111101111",
78859=>"010011010",
78860=>"000010000",
78861=>"000000000",
78862=>"110110100",
78863=>"111000100",
78864=>"000001011",
78865=>"000100101",
78866=>"001111111",
78867=>"111100111",
78868=>"100011000",
78869=>"010000101",
78870=>"111011101",
78871=>"111000000",
78872=>"000011011",
78873=>"000010010",
78874=>"000001000",
78875=>"110111111",
78876=>"011011111",
78877=>"000100000",
78878=>"000000111",
78879=>"000101000",
78880=>"110001000",
78881=>"000000000",
78882=>"111100111",
78883=>"111001010",
78884=>"111010100",
78885=>"000001011",
78886=>"110110010",
78887=>"001000000",
78888=>"000000000",
78889=>"100000111",
78890=>"111111111",
78891=>"111011111",
78892=>"111011000",
78893=>"000000000",
78894=>"100000111",
78895=>"000000101",
78896=>"000000100",
78897=>"110110110",
78898=>"111011111",
78899=>"111100100",
78900=>"111100111",
78901=>"000110110",
78902=>"110111011",
78903=>"110100100",
78904=>"100100110",
78905=>"000100000",
78906=>"011111011",
78907=>"100101100",
78908=>"000000001",
78909=>"000100111",
78910=>"000111010",
78911=>"011000100",
78912=>"000111111",
78913=>"000000110",
78914=>"000111010",
78915=>"001110111",
78916=>"010111011",
78917=>"000000010",
78918=>"110010010",
78919=>"010011110",
78920=>"010110010",
78921=>"110010001",
78922=>"100100111",
78923=>"101101101",
78924=>"010010000",
78925=>"011011011",
78926=>"011011001",
78927=>"000100000",
78928=>"101000000",
78929=>"011111111",
78930=>"110000010",
78931=>"100010011",
78932=>"000000000",
78933=>"000011011",
78934=>"011110010",
78935=>"110000000",
78936=>"000110000",
78937=>"010011000",
78938=>"010000000",
78939=>"011010110",
78940=>"000000000",
78941=>"111010000",
78942=>"000000000",
78943=>"111111111",
78944=>"000010000",
78945=>"010010000",
78946=>"011111010",
78947=>"011000000",
78948=>"001010011",
78949=>"000001000",
78950=>"010110000",
78951=>"010011011",
78952=>"000100000",
78953=>"000000000",
78954=>"111011000",
78955=>"000011000",
78956=>"000101011",
78957=>"101111111",
78958=>"111000100",
78959=>"111111000",
78960=>"011000000",
78961=>"100100100",
78962=>"011111110",
78963=>"110011010",
78964=>"010100000",
78965=>"000000010",
78966=>"000000101",
78967=>"000010000",
78968=>"111000110",
78969=>"011011000",
78970=>"111111111",
78971=>"111010111",
78972=>"010000100",
78973=>"011011011",
78974=>"011101111",
78975=>"010110111",
78976=>"010111010",
78977=>"011101100",
78978=>"000101111",
78979=>"000111100",
78980=>"100111111",
78981=>"011111010",
78982=>"000100010",
78983=>"011110110",
78984=>"011010010",
78985=>"000111011",
78986=>"001000000",
78987=>"000000110",
78988=>"000000000",
78989=>"010010000",
78990=>"101000001",
78991=>"011010110",
78992=>"011010010",
78993=>"110000000",
78994=>"101000000",
78995=>"010111011",
78996=>"010110000",
78997=>"000111011",
78998=>"111111100",
78999=>"010110011",
79000=>"011101110",
79001=>"000000000",
79002=>"110100110",
79003=>"111111111",
79004=>"011011010",
79005=>"010011011",
79006=>"011101111",
79007=>"000011010",
79008=>"011011011",
79009=>"000000000",
79010=>"111010000",
79011=>"111111000",
79012=>"101100000",
79013=>"011010010",
79014=>"011000111",
79015=>"000000100",
79016=>"100100101",
79017=>"111110110",
79018=>"000000000",
79019=>"101101111",
79020=>"001001000",
79021=>"010111011",
79022=>"001000000",
79023=>"101111010",
79024=>"000001111",
79025=>"010011111",
79026=>"000011010",
79027=>"111111000",
79028=>"001000000",
79029=>"111100110",
79030=>"000001011",
79031=>"111000010",
79032=>"001110000",
79033=>"001001001",
79034=>"000000010",
79035=>"111111110",
79036=>"000000000",
79037=>"111111111",
79038=>"110010010",
79039=>"000110000",
79040=>"010111010",
79041=>"001000000",
79042=>"000000100",
79043=>"111000011",
79044=>"111111111",
79045=>"011000111",
79046=>"011110000",
79047=>"001011111",
79048=>"111000000",
79049=>"000011111",
79050=>"101111100",
79051=>"000010000",
79052=>"010011010",
79053=>"010100100",
79054=>"111010111",
79055=>"000000001",
79056=>"100011001",
79057=>"011010000",
79058=>"111111000",
79059=>"000010011",
79060=>"000000101",
79061=>"000000010",
79062=>"000010000",
79063=>"010000100",
79064=>"011000000",
79065=>"111100000",
79066=>"011011011",
79067=>"000111111",
79068=>"001111110",
79069=>"000101100",
79070=>"111111010",
79071=>"111101110",
79072=>"100111110",
79073=>"000000111",
79074=>"000000010",
79075=>"011011111",
79076=>"101100000",
79077=>"010111011",
79078=>"111110100",
79079=>"100000000",
79080=>"011000000",
79081=>"111100101",
79082=>"101101100",
79083=>"101000100",
79084=>"100100111",
79085=>"100111111",
79086=>"001111111",
79087=>"101000000",
79088=>"010100000",
79089=>"010111111",
79090=>"111111100",
79091=>"110000000",
79092=>"101011011",
79093=>"000000000",
79094=>"000010000",
79095=>"011011111",
79096=>"111111000",
79097=>"101100100",
79098=>"111110111",
79099=>"001000000",
79100=>"011111111",
79101=>"100000000",
79102=>"011011111",
79103=>"100000000",
79104=>"000001110",
79105=>"001000111",
79106=>"000001111",
79107=>"011000101",
79108=>"100100111",
79109=>"001000001",
79110=>"010000010",
79111=>"111100111",
79112=>"100111110",
79113=>"000010000",
79114=>"110001000",
79115=>"001001101",
79116=>"000000011",
79117=>"000001000",
79118=>"000100000",
79119=>"101101111",
79120=>"010100001",
79121=>"111000111",
79122=>"101000010",
79123=>"110000000",
79124=>"111111110",
79125=>"001101111",
79126=>"111011000",
79127=>"111111101",
79128=>"010001101",
79129=>"000000111",
79130=>"111110100",
79131=>"001000000",
79132=>"101101010",
79133=>"101000000",
79134=>"000010111",
79135=>"110101101",
79136=>"000000001",
79137=>"001001001",
79138=>"000000001",
79139=>"100100110",
79140=>"100000111",
79141=>"001000100",
79142=>"001111110",
79143=>"110010000",
79144=>"100111000",
79145=>"001110100",
79146=>"001101100",
79147=>"001101111",
79148=>"010000000",
79149=>"111000111",
79150=>"101000000",
79151=>"011111011",
79152=>"110000000",
79153=>"000110111",
79154=>"111111001",
79155=>"111110100",
79156=>"111010000",
79157=>"111000000",
79158=>"011000001",
79159=>"101111111",
79160=>"000001101",
79161=>"100000000",
79162=>"111011000",
79163=>"111010100",
79164=>"010011001",
79165=>"011000000",
79166=>"111001000",
79167=>"111001110",
79168=>"001010100",
79169=>"001111111",
79170=>"000010011",
79171=>"100000001",
79172=>"000111111",
79173=>"100101001",
79174=>"001000111",
79175=>"111001000",
79176=>"011101101",
79177=>"111001001",
79178=>"001011111",
79179=>"111111100",
79180=>"001001010",
79181=>"001001011",
79182=>"011111110",
79183=>"111000110",
79184=>"011011111",
79185=>"110000011",
79186=>"110000001",
79187=>"010000000",
79188=>"001001000",
79189=>"011000011",
79190=>"100110110",
79191=>"101101011",
79192=>"001111111",
79193=>"011101100",
79194=>"011011111",
79195=>"011001000",
79196=>"110110111",
79197=>"010110110",
79198=>"110111000",
79199=>"111100011",
79200=>"000111000",
79201=>"111111001",
79202=>"000101111",
79203=>"001100100",
79204=>"101101111",
79205=>"111010000",
79206=>"111000000",
79207=>"011111110",
79208=>"000110110",
79209=>"001010000",
79210=>"110110110",
79211=>"001101111",
79212=>"001001111",
79213=>"000000011",
79214=>"001011111",
79215=>"011001000",
79216=>"101111001",
79217=>"110111100",
79218=>"110110000",
79219=>"010000001",
79220=>"001111111",
79221=>"101111100",
79222=>"100011010",
79223=>"001001111",
79224=>"110110001",
79225=>"110110000",
79226=>"000101111",
79227=>"010111111",
79228=>"110000011",
79229=>"101010110",
79230=>"111001001",
79231=>"000000000",
79232=>"001000000",
79233=>"000000111",
79234=>"100100100",
79235=>"000100001",
79236=>"000100111",
79237=>"110100001",
79238=>"000110010",
79239=>"000001010",
79240=>"001011111",
79241=>"110110000",
79242=>"111111000",
79243=>"000101011",
79244=>"001111111",
79245=>"001101111",
79246=>"001100000",
79247=>"001100100",
79248=>"100000011",
79249=>"111110011",
79250=>"001000000",
79251=>"001000000",
79252=>"101001000",
79253=>"101110000",
79254=>"110000000",
79255=>"100100111",
79256=>"000000001",
79257=>"000111111",
79258=>"100111111",
79259=>"111000010",
79260=>"110010000",
79261=>"101100000",
79262=>"000000000",
79263=>"011000100",
79264=>"111011110",
79265=>"111000101",
79266=>"111000011",
79267=>"110010000",
79268=>"110111011",
79269=>"100100100",
79270=>"011111001",
79271=>"000101011",
79272=>"111110010",
79273=>"111111111",
79274=>"001111111",
79275=>"111001101",
79276=>"110011011",
79277=>"101111111",
79278=>"110100111",
79279=>"000000000",
79280=>"001000001",
79281=>"000010111",
79282=>"111000000",
79283=>"001101110",
79284=>"111010110",
79285=>"010010000",
79286=>"010101100",
79287=>"000001001",
79288=>"110110100",
79289=>"010000100",
79290=>"110110000",
79291=>"110000000",
79292=>"011010000",
79293=>"101001111",
79294=>"000010010",
79295=>"011110000",
79296=>"001000010",
79297=>"111010100",
79298=>"001000000",
79299=>"000110100",
79300=>"010110000",
79301=>"100101110",
79302=>"001111101",
79303=>"111101000",
79304=>"110101000",
79305=>"011011011",
79306=>"001001001",
79307=>"001111111",
79308=>"000000100",
79309=>"111001101",
79310=>"000001001",
79311=>"011111101",
79312=>"110001001",
79313=>"010111110",
79314=>"110100110",
79315=>"110100000",
79316=>"000000000",
79317=>"001001111",
79318=>"101000000",
79319=>"110000000",
79320=>"101111111",
79321=>"110100000",
79322=>"010010000",
79323=>"101110111",
79324=>"010010000",
79325=>"001101111",
79326=>"000110000",
79327=>"110001001",
79328=>"000010010",
79329=>"111101101",
79330=>"110110010",
79331=>"111100100",
79332=>"111010000",
79333=>"001000100",
79334=>"100000000",
79335=>"000111111",
79336=>"001001001",
79337=>"000011001",
79338=>"011000000",
79339=>"111101001",
79340=>"001111011",
79341=>"000001101",
79342=>"001000010",
79343=>"111111110",
79344=>"000001100",
79345=>"011011001",
79346=>"110111000",
79347=>"100000000",
79348=>"000000011",
79349=>"010110110",
79350=>"000000000",
79351=>"000010000",
79352=>"000000110",
79353=>"000000000",
79354=>"000001110",
79355=>"111001000",
79356=>"111110010",
79357=>"000110010",
79358=>"011101001",
79359=>"000000011",
79360=>"011111100",
79361=>"111000010",
79362=>"000000001",
79363=>"000000000",
79364=>"000111000",
79365=>"011001111",
79366=>"000001111",
79367=>"011000010",
79368=>"001000010",
79369=>"000000001",
79370=>"100110011",
79371=>"100001100",
79372=>"000000101",
79373=>"010111101",
79374=>"100011110",
79375=>"111110100",
79376=>"001000001",
79377=>"010010000",
79378=>"000000010",
79379=>"010110111",
79380=>"000001000",
79381=>"000000101",
79382=>"010111001",
79383=>"111111110",
79384=>"000000000",
79385=>"111011111",
79386=>"110011111",
79387=>"111011001",
79388=>"111000001",
79389=>"111000000",
79390=>"000101101",
79391=>"000001011",
79392=>"001111111",
79393=>"000011111",
79394=>"111000001",
79395=>"000000000",
79396=>"110100100",
79397=>"111111011",
79398=>"011010111",
79399=>"101100000",
79400=>"110010111",
79401=>"100000011",
79402=>"000111110",
79403=>"111011000",
79404=>"011000000",
79405=>"000000000",
79406=>"010001110",
79407=>"111001111",
79408=>"111001000",
79409=>"110101001",
79410=>"100000000",
79411=>"111000111",
79412=>"101000111",
79413=>"111111011",
79414=>"110011011",
79415=>"111001000",
79416=>"001001111",
79417=>"000101010",
79418=>"001001000",
79419=>"010000101",
79420=>"111011010",
79421=>"011010000",
79422=>"000001011",
79423=>"100001000",
79424=>"111111111",
79425=>"111111001",
79426=>"101001011",
79427=>"000000011",
79428=>"110110000",
79429=>"101110110",
79430=>"011111010",
79431=>"101100111",
79432=>"000000110",
79433=>"111000111",
79434=>"101001001",
79435=>"001100111",
79436=>"000000111",
79437=>"011111001",
79438=>"001001101",
79439=>"111000011",
79440=>"101111001",
79441=>"000111011",
79442=>"000111111",
79443=>"001001000",
79444=>"101100000",
79445=>"111110011",
79446=>"001001100",
79447=>"100000000",
79448=>"111011111",
79449=>"000000011",
79450=>"110101000",
79451=>"000010110",
79452=>"111111010",
79453=>"100100100",
79454=>"110110000",
79455=>"001010100",
79456=>"111111111",
79457=>"000000000",
79458=>"001111111",
79459=>"111110010",
79460=>"000001011",
79461=>"000000111",
79462=>"001111111",
79463=>"000000111",
79464=>"001101000",
79465=>"111000111",
79466=>"000110110",
79467=>"001111111",
79468=>"111001001",
79469=>"111111100",
79470=>"101101000",
79471=>"101001001",
79472=>"000010000",
79473=>"000111111",
79474=>"000110110",
79475=>"000000100",
79476=>"000000110",
79477=>"000000000",
79478=>"001001000",
79479=>"000000101",
79480=>"000100110",
79481=>"111000000",
79482=>"000000111",
79483=>"000101000",
79484=>"111001000",
79485=>"101000011",
79486=>"000000111",
79487=>"001001001",
79488=>"111101101",
79489=>"001011001",
79490=>"000110111",
79491=>"000000011",
79492=>"000000000",
79493=>"000111010",
79494=>"111100100",
79495=>"110000011",
79496=>"000000111",
79497=>"000000001",
79498=>"010010011",
79499=>"000110101",
79500=>"010110000",
79501=>"111111101",
79502=>"000111111",
79503=>"000000001",
79504=>"111100111",
79505=>"101000000",
79506=>"000000101",
79507=>"001000101",
79508=>"000000100",
79509=>"000001010",
79510=>"111010110",
79511=>"000110110",
79512=>"000001101",
79513=>"111001000",
79514=>"011011000",
79515=>"000000010",
79516=>"000000111",
79517=>"000111000",
79518=>"000111010",
79519=>"000001000",
79520=>"000011011",
79521=>"010111111",
79522=>"001111010",
79523=>"000011111",
79524=>"000110010",
79525=>"001001110",
79526=>"000010111",
79527=>"101101101",
79528=>"110010001",
79529=>"101101011",
79530=>"110111111",
79531=>"000000001",
79532=>"011000101",
79533=>"001000011",
79534=>"111111010",
79535=>"000111101",
79536=>"111101000",
79537=>"111110100",
79538=>"010000000",
79539=>"011100000",
79540=>"100111110",
79541=>"100110000",
79542=>"010000111",
79543=>"111111000",
79544=>"111110110",
79545=>"001001000",
79546=>"111001110",
79547=>"111001101",
79548=>"001000001",
79549=>"000110000",
79550=>"101110101",
79551=>"111000110",
79552=>"110000000",
79553=>"000010010",
79554=>"000100100",
79555=>"111011110",
79556=>"000111000",
79557=>"110001011",
79558=>"101001001",
79559=>"000111100",
79560=>"000000100",
79561=>"110001000",
79562=>"000111100",
79563=>"000000111",
79564=>"101111010",
79565=>"110101000",
79566=>"111101000",
79567=>"110111101",
79568=>"011111111",
79569=>"000111011",
79570=>"000000100",
79571=>"101111010",
79572=>"000000100",
79573=>"111110000",
79574=>"000000101",
79575=>"110101000",
79576=>"010110000",
79577=>"000001111",
79578=>"001000101",
79579=>"001000111",
79580=>"110010110",
79581=>"000001000",
79582=>"000011100",
79583=>"011001011",
79584=>"000000001",
79585=>"000000011",
79586=>"000100110",
79587=>"111000101",
79588=>"000000111",
79589=>"111111000",
79590=>"001101010",
79591=>"111111000",
79592=>"101000111",
79593=>"111000000",
79594=>"011010110",
79595=>"111001101",
79596=>"000010111",
79597=>"000010000",
79598=>"100000000",
79599=>"000111000",
79600=>"000110101",
79601=>"010001100",
79602=>"000000000",
79603=>"010111111",
79604=>"100111001",
79605=>"000001111",
79606=>"010000110",
79607=>"110011011",
79608=>"011111000",
79609=>"001000000",
79610=>"111111111",
79611=>"000000101",
79612=>"111111001",
79613=>"001010011",
79614=>"101001000",
79615=>"000110110",
79616=>"011111011",
79617=>"000000001",
79618=>"101101101",
79619=>"000000000",
79620=>"011101100",
79621=>"011111000",
79622=>"111001001",
79623=>"111111111",
79624=>"111111000",
79625=>"001000111",
79626=>"000100110",
79627=>"000000000",
79628=>"110111000",
79629=>"000000000",
79630=>"111111011",
79631=>"000000111",
79632=>"010010000",
79633=>"100111111",
79634=>"100100111",
79635=>"111101111",
79636=>"000000111",
79637=>"000000101",
79638=>"100000000",
79639=>"101100001",
79640=>"111111011",
79641=>"000111110",
79642=>"110000000",
79643=>"000000000",
79644=>"101000000",
79645=>"000111110",
79646=>"111000000",
79647=>"010100000",
79648=>"001100100",
79649=>"101000000",
79650=>"000000000",
79651=>"111110000",
79652=>"000001000",
79653=>"110111111",
79654=>"010010000",
79655=>"111000000",
79656=>"100100000",
79657=>"101111110",
79658=>"100100100",
79659=>"111000111",
79660=>"101101001",
79661=>"111010011",
79662=>"111001000",
79663=>"011001011",
79664=>"100111000",
79665=>"100100000",
79666=>"001111011",
79667=>"000000001",
79668=>"000000000",
79669=>"000000010",
79670=>"000000000",
79671=>"101000000",
79672=>"111010010",
79673=>"000100110",
79674=>"100100000",
79675=>"101101101",
79676=>"100010110",
79677=>"111010111",
79678=>"000000111",
79679=>"011001001",
79680=>"100111111",
79681=>"010111100",
79682=>"110111010",
79683=>"000111100",
79684=>"010000000",
79685=>"110010000",
79686=>"101101111",
79687=>"000000001",
79688=>"011001000",
79689=>"000111010",
79690=>"110010001",
79691=>"000100111",
79692=>"101101111",
79693=>"010111010",
79694=>"001001001",
79695=>"111111111",
79696=>"000000101",
79697=>"010111111",
79698=>"000011100",
79699=>"000111011",
79700=>"000111111",
79701=>"000000010",
79702=>"011111000",
79703=>"000000101",
79704=>"111000000",
79705=>"100100100",
79706=>"100100000",
79707=>"010100100",
79708=>"010000000",
79709=>"001001000",
79710=>"111111000",
79711=>"010001011",
79712=>"111000000",
79713=>"100001000",
79714=>"110000111",
79715=>"001001011",
79716=>"000000110",
79717=>"101111000",
79718=>"101001100",
79719=>"101000100",
79720=>"000000000",
79721=>"001100000",
79722=>"111010111",
79723=>"110110100",
79724=>"110111010",
79725=>"001111111",
79726=>"011001111",
79727=>"000111111",
79728=>"011011110",
79729=>"000000000",
79730=>"000000100",
79731=>"111101111",
79732=>"101010101",
79733=>"011000000",
79734=>"010111100",
79735=>"010111111",
79736=>"110001001",
79737=>"111111000",
79738=>"000100111",
79739=>"111111011",
79740=>"101000101",
79741=>"100100100",
79742=>"000000011",
79743=>"110110001",
79744=>"000100111",
79745=>"101111111",
79746=>"000111100",
79747=>"010000110",
79748=>"000110111",
79749=>"110111011",
79750=>"000100000",
79751=>"011001000",
79752=>"100100001",
79753=>"000000110",
79754=>"110010000",
79755=>"111010011",
79756=>"001001101",
79757=>"101101111",
79758=>"111110010",
79759=>"100110111",
79760=>"100110000",
79761=>"100000000",
79762=>"101111111",
79763=>"101000110",
79764=>"101010111",
79765=>"000000000",
79766=>"111011010",
79767=>"011111111",
79768=>"111111011",
79769=>"100010000",
79770=>"110111111",
79771=>"101111010",
79772=>"110111000",
79773=>"010010000",
79774=>"111111010",
79775=>"001001000",
79776=>"110110000",
79777=>"000111101",
79778=>"111111010",
79779=>"111000000",
79780=>"001110111",
79781=>"110001001",
79782=>"110010001",
79783=>"000010010",
79784=>"000110111",
79785=>"111111110",
79786=>"101101000",
79787=>"000000100",
79788=>"111111000",
79789=>"001111111",
79790=>"000001001",
79791=>"011011010",
79792=>"001000000",
79793=>"111011001",
79794=>"111111000",
79795=>"100000000",
79796=>"101011000",
79797=>"100000111",
79798=>"100100000",
79799=>"111010110",
79800=>"001100000",
79801=>"101100111",
79802=>"101110110",
79803=>"010010000",
79804=>"101111111",
79805=>"110110000",
79806=>"111011000",
79807=>"000000000",
79808=>"000000101",
79809=>"111101111",
79810=>"101111001",
79811=>"110111000",
79812=>"000010010",
79813=>"001101110",
79814=>"010010000",
79815=>"100100101",
79816=>"111010010",
79817=>"111011011",
79818=>"101000000",
79819=>"001001011",
79820=>"111101101",
79821=>"001101101",
79822=>"101101101",
79823=>"010000000",
79824=>"010001111",
79825=>"110110110",
79826=>"100111111",
79827=>"110000110",
79828=>"000000111",
79829=>"110110000",
79830=>"111111000",
79831=>"111000000",
79832=>"000000111",
79833=>"001000000",
79834=>"111111000",
79835=>"001111111",
79836=>"001001100",
79837=>"111111000",
79838=>"000101101",
79839=>"100001001",
79840=>"110010000",
79841=>"010111101",
79842=>"000000101",
79843=>"111011000",
79844=>"111100001",
79845=>"000000000",
79846=>"000000010",
79847=>"000000000",
79848=>"111101111",
79849=>"000000000",
79850=>"000001011",
79851=>"100000001",
79852=>"010111000",
79853=>"000000000",
79854=>"010010000",
79855=>"000101111",
79856=>"101000000",
79857=>"100001001",
79858=>"101101110",
79859=>"111101000",
79860=>"010011001",
79861=>"000000101",
79862=>"000000100",
79863=>"100101001",
79864=>"000000000",
79865=>"001011110",
79866=>"000111111",
79867=>"100101101",
79868=>"110110000",
79869=>"000000001",
79870=>"011111001",
79871=>"110110111",
79872=>"101111110",
79873=>"111111010",
79874=>"111111100",
79875=>"111101000",
79876=>"111110100",
79877=>"111111000",
79878=>"100000000",
79879=>"000000000",
79880=>"001001001",
79881=>"111111100",
79882=>"000001011",
79883=>"111000001",
79884=>"000000001",
79885=>"111010010",
79886=>"100100000",
79887=>"010010001",
79888=>"001010001",
79889=>"100000100",
79890=>"001000000",
79891=>"000111111",
79892=>"000100110",
79893=>"000000000",
79894=>"111111011",
79895=>"010111111",
79896=>"101101111",
79897=>"000000000",
79898=>"111100111",
79899=>"000000000",
79900=>"000101000",
79901=>"101101010",
79902=>"000001000",
79903=>"100000110",
79904=>"111111011",
79905=>"111111111",
79906=>"110000000",
79907=>"101100000",
79908=>"010110110",
79909=>"001000001",
79910=>"000000111",
79911=>"000100101",
79912=>"111111111",
79913=>"001001010",
79914=>"000010011",
79915=>"101111111",
79916=>"000000011",
79917=>"000000110",
79918=>"011111110",
79919=>"111111111",
79920=>"111111010",
79921=>"001000011",
79922=>"010110000",
79923=>"000001001",
79924=>"111001000",
79925=>"000000001",
79926=>"001011011",
79927=>"000001000",
79928=>"000000000",
79929=>"000001000",
79930=>"111111110",
79931=>"011101100",
79932=>"011011011",
79933=>"010111111",
79934=>"000111111",
79935=>"101111101",
79936=>"000111000",
79937=>"101111101",
79938=>"111101111",
79939=>"111000110",
79940=>"000000111",
79941=>"001101101",
79942=>"000001000",
79943=>"011101110",
79944=>"100000011",
79945=>"111000000",
79946=>"111111111",
79947=>"000110000",
79948=>"000000000",
79949=>"110100110",
79950=>"010011011",
79951=>"001000000",
79952=>"111101100",
79953=>"111111100",
79954=>"101111110",
79955=>"110011111",
79956=>"111001111",
79957=>"001000011",
79958=>"100111111",
79959=>"000000111",
79960=>"111111001",
79961=>"000100010",
79962=>"111110011",
79963=>"000110111",
79964=>"111101011",
79965=>"110110110",
79966=>"000111000",
79967=>"110000001",
79968=>"001001111",
79969=>"010000010",
79970=>"111101101",
79971=>"111111011",
79972=>"011111011",
79973=>"000000000",
79974=>"010010000",
79975=>"000101111",
79976=>"101110111",
79977=>"000000011",
79978=>"111111010",
79979=>"011111111",
79980=>"000011011",
79981=>"000111000",
79982=>"100100000",
79983=>"000001000",
79984=>"110110110",
79985=>"000010000",
79986=>"001111011",
79987=>"000001111",
79988=>"111111111",
79989=>"111110110",
79990=>"111101000",
79991=>"001001110",
79992=>"111101000",
79993=>"111101100",
79994=>"000010010",
79995=>"111110010",
79996=>"011001001",
79997=>"011111111",
79998=>"000101111",
79999=>"000001111",
80000=>"111111111",
80001=>"011111110",
80002=>"001010010",
80003=>"001101111",
80004=>"111000000",
80005=>"100111100",
80006=>"100100110",
80007=>"000011100",
80008=>"000010111",
80009=>"001001001",
80010=>"000101111",
80011=>"000100110",
80012=>"011111001",
80013=>"001000100",
80014=>"111111011",
80015=>"111110000",
80016=>"100100110",
80017=>"111000000",
80018=>"110111001",
80019=>"110000000",
80020=>"000000000",
80021=>"111111111",
80022=>"000010000",
80023=>"101111100",
80024=>"000000000",
80025=>"000011101",
80026=>"111111110",
80027=>"111111111",
80028=>"000000000",
80029=>"101011101",
80030=>"100111111",
80031=>"000000110",
80032=>"100111110",
80033=>"111011101",
80034=>"001101011",
80035=>"000000000",
80036=>"111111110",
80037=>"000110111",
80038=>"000000110",
80039=>"100111111",
80040=>"010101000",
80041=>"000001001",
80042=>"111111000",
80043=>"001000001",
80044=>"111101111",
80045=>"000000000",
80046=>"001011011",
80047=>"100101000",
80048=>"111111000",
80049=>"110110010",
80050=>"111111111",
80051=>"111000000",
80052=>"000001111",
80053=>"000010011",
80054=>"000001110",
80055=>"010111000",
80056=>"110100010",
80057=>"000001001",
80058=>"111111111",
80059=>"111110000",
80060=>"000000010",
80061=>"111111111",
80062=>"100100101",
80063=>"010011000",
80064=>"000111010",
80065=>"001001111",
80066=>"000000001",
80067=>"001001001",
80068=>"000000001",
80069=>"111000110",
80070=>"000001110",
80071=>"111110000",
80072=>"000000111",
80073=>"000001011",
80074=>"000111011",
80075=>"000101111",
80076=>"101000100",
80077=>"111000000",
80078=>"011101101",
80079=>"111010101",
80080=>"111011011",
80081=>"111110010",
80082=>"000000000",
80083=>"000101111",
80084=>"010000000",
80085=>"011111011",
80086=>"110110000",
80087=>"000001110",
80088=>"000000111",
80089=>"000000000",
80090=>"010111111",
80091=>"111111101",
80092=>"000111100",
80093=>"111101111",
80094=>"011010000",
80095=>"000000010",
80096=>"000000000",
80097=>"111000000",
80098=>"111000001",
80099=>"001011011",
80100=>"001101111",
80101=>"111000000",
80102=>"111111110",
80103=>"100101010",
80104=>"111100110",
80105=>"011000000",
80106=>"000000100",
80107=>"110011011",
80108=>"000000000",
80109=>"001111111",
80110=>"111111000",
80111=>"111111010",
80112=>"000000011",
80113=>"010110110",
80114=>"111111111",
80115=>"000001111",
80116=>"001111011",
80117=>"111111000",
80118=>"010010010",
80119=>"111000100",
80120=>"000110110",
80121=>"100001101",
80122=>"011110000",
80123=>"000100000",
80124=>"000000010",
80125=>"101000000",
80126=>"101011010",
80127=>"000000000",
80128=>"000000011",
80129=>"111111001",
80130=>"000111010",
80131=>"000000000",
80132=>"000000000",
80133=>"000010010",
80134=>"101111000",
80135=>"000000000",
80136=>"000001001",
80137=>"000011001",
80138=>"000000001",
80139=>"000000110",
80140=>"110000000",
80141=>"100111111",
80142=>"100100000",
80143=>"000011111",
80144=>"000000111",
80145=>"111100000",
80146=>"001000010",
80147=>"101111101",
80148=>"000000000",
80149=>"110111100",
80150=>"000111111",
80151=>"111000111",
80152=>"010000000",
80153=>"000000000",
80154=>"111100000",
80155=>"111111111",
80156=>"101000100",
80157=>"001000000",
80158=>"000000110",
80159=>"101101001",
80160=>"000010110",
80161=>"111110011",
80162=>"010101100",
80163=>"010111011",
80164=>"111011011",
80165=>"100001000",
80166=>"110100000",
80167=>"000000000",
80168=>"111111101",
80169=>"000101111",
80170=>"000000001",
80171=>"000000110",
80172=>"000010111",
80173=>"000000000",
80174=>"000000000",
80175=>"000000000",
80176=>"101111010",
80177=>"111011110",
80178=>"010001101",
80179=>"111001100",
80180=>"000000000",
80181=>"000000010",
80182=>"000000000",
80183=>"001000001",
80184=>"111000000",
80185=>"111101000",
80186=>"000000011",
80187=>"110110000",
80188=>"111111110",
80189=>"111111111",
80190=>"111100010",
80191=>"101111111",
80192=>"100010010",
80193=>"000001010",
80194=>"110111000",
80195=>"111011111",
80196=>"000000010",
80197=>"101001111",
80198=>"100110011",
80199=>"001001110",
80200=>"110111000",
80201=>"110000000",
80202=>"111101111",
80203=>"010001000",
80204=>"111100000",
80205=>"101110100",
80206=>"011110011",
80207=>"000000000",
80208=>"101101101",
80209=>"111101111",
80210=>"111111100",
80211=>"100000000",
80212=>"111111110",
80213=>"100011001",
80214=>"001000001",
80215=>"000000000",
80216=>"001111111",
80217=>"011001000",
80218=>"010111110",
80219=>"100111111",
80220=>"000001011",
80221=>"000110100",
80222=>"011110000",
80223=>"110100000",
80224=>"000000000",
80225=>"000101101",
80226=>"111010010",
80227=>"001001001",
80228=>"100000010",
80229=>"101111111",
80230=>"000000000",
80231=>"000000001",
80232=>"111010010",
80233=>"000000110",
80234=>"010110110",
80235=>"001111111",
80236=>"000000111",
80237=>"000001101",
80238=>"001000000",
80239=>"000000000",
80240=>"110111101",
80241=>"010111111",
80242=>"000000000",
80243=>"000000101",
80244=>"000111101",
80245=>"000010000",
80246=>"100000111",
80247=>"011101101",
80248=>"111111111",
80249=>"111110101",
80250=>"010000111",
80251=>"111111000",
80252=>"000001100",
80253=>"000011010",
80254=>"010111100",
80255=>"011111010",
80256=>"000101101",
80257=>"101000000",
80258=>"000001011",
80259=>"001001001",
80260=>"111000000",
80261=>"000111000",
80262=>"111110100",
80263=>"011100000",
80264=>"001011000",
80265=>"111111000",
80266=>"001000111",
80267=>"000000110",
80268=>"001000000",
80269=>"111010000",
80270=>"100000010",
80271=>"000000000",
80272=>"010100000",
80273=>"111111111",
80274=>"000000101",
80275=>"000000000",
80276=>"111111100",
80277=>"001000010",
80278=>"011011000",
80279=>"110100110",
80280=>"000010111",
80281=>"000000101",
80282=>"100111111",
80283=>"000011000",
80284=>"010010000",
80285=>"110111011",
80286=>"010111111",
80287=>"000000000",
80288=>"000111000",
80289=>"111000011",
80290=>"000000000",
80291=>"001000000",
80292=>"100000000",
80293=>"000101111",
80294=>"011001011",
80295=>"000000111",
80296=>"111111001",
80297=>"000000101",
80298=>"111110110",
80299=>"010010000",
80300=>"001101111",
80301=>"100100111",
80302=>"010110000",
80303=>"000011011",
80304=>"100111110",
80305=>"111101000",
80306=>"111101000",
80307=>"000000001",
80308=>"000001100",
80309=>"000000011",
80310=>"000000000",
80311=>"000111111",
80312=>"111111001",
80313=>"100101100",
80314=>"111111111",
80315=>"100111111",
80316=>"000000001",
80317=>"111111000",
80318=>"100100000",
80319=>"000011111",
80320=>"101101010",
80321=>"001000000",
80322=>"111101001",
80323=>"000001001",
80324=>"000000000",
80325=>"001010000",
80326=>"000000001",
80327=>"111101001",
80328=>"001000001",
80329=>"111001000",
80330=>"000000101",
80331=>"010111110",
80332=>"010011111",
80333=>"010000001",
80334=>"000000101",
80335=>"111111110",
80336=>"000111000",
80337=>"000100110",
80338=>"011101000",
80339=>"000000101",
80340=>"111110000",
80341=>"100100000",
80342=>"001000000",
80343=>"000111111",
80344=>"000000000",
80345=>"000000000",
80346=>"011010001",
80347=>"000110111",
80348=>"000110111",
80349=>"000111111",
80350=>"000000000",
80351=>"111111101",
80352=>"110111110",
80353=>"111011010",
80354=>"111111101",
80355=>"000001101",
80356=>"000000100",
80357=>"100110111",
80358=>"111111010",
80359=>"000100111",
80360=>"111111111",
80361=>"000001101",
80362=>"000000110",
80363=>"000000000",
80364=>"001000000",
80365=>"001000101",
80366=>"000111000",
80367=>"010111101",
80368=>"000000101",
80369=>"000000000",
80370=>"000101111",
80371=>"010110101",
80372=>"000001000",
80373=>"000110101",
80374=>"111111000",
80375=>"000010000",
80376=>"000000101",
80377=>"000000000",
80378=>"000000100",
80379=>"000000011",
80380=>"111011000",
80381=>"111111111",
80382=>"000110011",
80383=>"100100010",
80384=>"001000001",
80385=>"000000000",
80386=>"010111010",
80387=>"101000000",
80388=>"000000100",
80389=>"000000001",
80390=>"101111101",
80391=>"110000000",
80392=>"000000000",
80393=>"110001000",
80394=>"000100100",
80395=>"110111111",
80396=>"001011011",
80397=>"111001001",
80398=>"000111011",
80399=>"000000000",
80400=>"111000100",
80401=>"001110000",
80402=>"000000000",
80403=>"110000111",
80404=>"000000000",
80405=>"010111111",
80406=>"001111100",
80407=>"010010110",
80408=>"000000000",
80409=>"011000100",
80410=>"000000101",
80411=>"111111001",
80412=>"101010110",
80413=>"001111000",
80414=>"101000000",
80415=>"111111001",
80416=>"111111111",
80417=>"111000111",
80418=>"110111000",
80419=>"111111111",
80420=>"111001001",
80421=>"001011101",
80422=>"000111000",
80423=>"110001101",
80424=>"111001111",
80425=>"010000000",
80426=>"111111111",
80427=>"000111000",
80428=>"111110110",
80429=>"101000001",
80430=>"101111111",
80431=>"111000100",
80432=>"000000010",
80433=>"000000000",
80434=>"000000000",
80435=>"110110000",
80436=>"000001001",
80437=>"000000000",
80438=>"110111111",
80439=>"111001000",
80440=>"001000000",
80441=>"100000101",
80442=>"000000000",
80443=>"000000010",
80444=>"110011100",
80445=>"111111111",
80446=>"000000101",
80447=>"000000000",
80448=>"111000110",
80449=>"111111111",
80450=>"110100000",
80451=>"001101001",
80452=>"000000100",
80453=>"000000000",
80454=>"111101110",
80455=>"000111111",
80456=>"111111111",
80457=>"000000101",
80458=>"101000101",
80459=>"111111110",
80460=>"000100110",
80461=>"011000000",
80462=>"011001000",
80463=>"100011111",
80464=>"100101111",
80465=>"111111010",
80466=>"001000000",
80467=>"001010100",
80468=>"000000000",
80469=>"000111100",
80470=>"111001001",
80471=>"010000010",
80472=>"010010010",
80473=>"110110111",
80474=>"010111101",
80475=>"001000100",
80476=>"101101101",
80477=>"000000001",
80478=>"010111111",
80479=>"100100111",
80480=>"111101111",
80481=>"101111111",
80482=>"000000010",
80483=>"000111110",
80484=>"000001100",
80485=>"101000011",
80486=>"100110111",
80487=>"111000000",
80488=>"000000000",
80489=>"000000000",
80490=>"101000001",
80491=>"100110111",
80492=>"111101000",
80493=>"101000000",
80494=>"111000000",
80495=>"111000000",
80496=>"101001000",
80497=>"000000000",
80498=>"111111111",
80499=>"111100101",
80500=>"010100000",
80501=>"101000000",
80502=>"010000000",
80503=>"110101000",
80504=>"010111011",
80505=>"111111111",
80506=>"000011111",
80507=>"011001000",
80508=>"000100100",
80509=>"100000000",
80510=>"111111111",
80511=>"000111111",
80512=>"101101000",
80513=>"000111011",
80514=>"000000000",
80515=>"111000111",
80516=>"101000000",
80517=>"100000000",
80518=>"011111011",
80519=>"100110111",
80520=>"000000001",
80521=>"111111111",
80522=>"111101100",
80523=>"111101010",
80524=>"010010000",
80525=>"101111100",
80526=>"110111111",
80527=>"001001000",
80528=>"000000000",
80529=>"111111101",
80530=>"111101101",
80531=>"111010000",
80532=>"001011111",
80533=>"111000000",
80534=>"011111111",
80535=>"000000011",
80536=>"001000000",
80537=>"000000000",
80538=>"111111111",
80539=>"110010001",
80540=>"000000000",
80541=>"000000000",
80542=>"000000101",
80543=>"000000111",
80544=>"110111110",
80545=>"111011111",
80546=>"111111111",
80547=>"110000000",
80548=>"110101000",
80549=>"010001001",
80550=>"100100100",
80551=>"000000010",
80552=>"111111000",
80553=>"110101100",
80554=>"111010000",
80555=>"000000111",
80556=>"101100111",
80557=>"111000000",
80558=>"000000100",
80559=>"100111111",
80560=>"000100000",
80561=>"111111111",
80562=>"000001011",
80563=>"000010100",
80564=>"100100000",
80565=>"110111010",
80566=>"000000000",
80567=>"000000010",
80568=>"011010001",
80569=>"001000101",
80570=>"111111001",
80571=>"111001000",
80572=>"000100000",
80573=>"000011010",
80574=>"000000000",
80575=>"011000000",
80576=>"111101000",
80577=>"000110000",
80578=>"111101000",
80579=>"001001001",
80580=>"100000000",
80581=>"100110001",
80582=>"111100000",
80583=>"000000110",
80584=>"001000010",
80585=>"111111111",
80586=>"000000000",
80587=>"111101111",
80588=>"011000100",
80589=>"000001010",
80590=>"101000011",
80591=>"000000000",
80592=>"111111111",
80593=>"111011011",
80594=>"100011000",
80595=>"001000000",
80596=>"001001111",
80597=>"100101100",
80598=>"000000000",
80599=>"000000000",
80600=>"111000011",
80601=>"010010111",
80602=>"011001001",
80603=>"000010000",
80604=>"001111011",
80605=>"000000000",
80606=>"010110110",
80607=>"111001100",
80608=>"011100001",
80609=>"000011101",
80610=>"001000101",
80611=>"000011000",
80612=>"101001101",
80613=>"011111100",
80614=>"000001111",
80615=>"001101001",
80616=>"000000000",
80617=>"100000100",
80618=>"000000001",
80619=>"010011000",
80620=>"000001000",
80621=>"100000100",
80622=>"000010000",
80623=>"111100000",
80624=>"111000000",
80625=>"011111110",
80626=>"111111000",
80627=>"011001011",
80628=>"110110100",
80629=>"000111111",
80630=>"000000000",
80631=>"000010000",
80632=>"011010011",
80633=>"001000001",
80634=>"101100100",
80635=>"101010010",
80636=>"011111011",
80637=>"110111111",
80638=>"100000000",
80639=>"001000000",
80640=>"011101100",
80641=>"111000000",
80642=>"000000000",
80643=>"111010110",
80644=>"110110000",
80645=>"101110110",
80646=>"010111000",
80647=>"000000001",
80648=>"111011110",
80649=>"000001110",
80650=>"000011011",
80651=>"000010000",
80652=>"000000111",
80653=>"110000000",
80654=>"110100010",
80655=>"111101100",
80656=>"110010011",
80657=>"111011000",
80658=>"010000000",
80659=>"000000000",
80660=>"111000000",
80661=>"111111111",
80662=>"001111111",
80663=>"111111000",
80664=>"000000011",
80665=>"111111111",
80666=>"000000000",
80667=>"000111000",
80668=>"110100000",
80669=>"000100001",
80670=>"000110100",
80671=>"000000111",
80672=>"101001000",
80673=>"111001001",
80674=>"111101101",
80675=>"100111110",
80676=>"110111100",
80677=>"100001011",
80678=>"000000010",
80679=>"010100010",
80680=>"000000001",
80681=>"011001111",
80682=>"100110110",
80683=>"110100110",
80684=>"000000011",
80685=>"000000111",
80686=>"111101110",
80687=>"111011111",
80688=>"010010000",
80689=>"000110100",
80690=>"110001000",
80691=>"111000000",
80692=>"111111101",
80693=>"000000000",
80694=>"000000101",
80695=>"011111011",
80696=>"001000000",
80697=>"111000000",
80698=>"111000000",
80699=>"011111100",
80700=>"111101000",
80701=>"000111111",
80702=>"000000000",
80703=>"010001111",
80704=>"111110111",
80705=>"000101111",
80706=>"101111111",
80707=>"000111111",
80708=>"000110110",
80709=>"001010000",
80710=>"000111011",
80711=>"111111111",
80712=>"110001111",
80713=>"000101111",
80714=>"101000000",
80715=>"111111011",
80716=>"000011110",
80717=>"011111111",
80718=>"000111011",
80719=>"010000001",
80720=>"000001000",
80721=>"101010111",
80722=>"110101100",
80723=>"101000000",
80724=>"000100111",
80725=>"011001001",
80726=>"010011101",
80727=>"100111000",
80728=>"000000111",
80729=>"000110100",
80730=>"111000100",
80731=>"011100010",
80732=>"000111111",
80733=>"111101100",
80734=>"111001000",
80735=>"000011111",
80736=>"000110111",
80737=>"000111111",
80738=>"000000111",
80739=>"111000010",
80740=>"111001100",
80741=>"010011001",
80742=>"000110110",
80743=>"101011111",
80744=>"110111111",
80745=>"000010111",
80746=>"000010111",
80747=>"111001111",
80748=>"111111011",
80749=>"111111000",
80750=>"011000001",
80751=>"111111011",
80752=>"001011011",
80753=>"000010000",
80754=>"000000110",
80755=>"001001000",
80756=>"000000110",
80757=>"100111111",
80758=>"111111011",
80759=>"000001100",
80760=>"000001010",
80761=>"110111101",
80762=>"010111101",
80763=>"110111101",
80764=>"001001000",
80765=>"111000011",
80766=>"001101110",
80767=>"000000111",
80768=>"110111110",
80769=>"111011000",
80770=>"000111111",
80771=>"111111111",
80772=>"010000111",
80773=>"000000100",
80774=>"001000110",
80775=>"000110100",
80776=>"010110110",
80777=>"100111111",
80778=>"010110100",
80779=>"101111000",
80780=>"111000001",
80781=>"101111111",
80782=>"111000000",
80783=>"000101000",
80784=>"110100100",
80785=>"001101111",
80786=>"111001101",
80787=>"000000100",
80788=>"111110000",
80789=>"111000000",
80790=>"111111111",
80791=>"010010011",
80792=>"000111010",
80793=>"100101011",
80794=>"000001111",
80795=>"010011101",
80796=>"100001111",
80797=>"000110111",
80798=>"001010100",
80799=>"000111111",
80800=>"011110000",
80801=>"111111000",
80802=>"000000101",
80803=>"100001100",
80804=>"111101010",
80805=>"000010010",
80806=>"111101100",
80807=>"000001000",
80808=>"111110000",
80809=>"100101111",
80810=>"111000000",
80811=>"011010000",
80812=>"111101111",
80813=>"000000111",
80814=>"100000001",
80815=>"110011011",
80816=>"000110010",
80817=>"001000100",
80818=>"101111011",
80819=>"000011011",
80820=>"010100110",
80821=>"111101000",
80822=>"010000011",
80823=>"111000000",
80824=>"111001100",
80825=>"000000001",
80826=>"111000000",
80827=>"111001110",
80828=>"101100111",
80829=>"000000111",
80830=>"100110111",
80831=>"000000100",
80832=>"101000111",
80833=>"111100000",
80834=>"111011000",
80835=>"110100110",
80836=>"000101010",
80837=>"111111001",
80838=>"110111111",
80839=>"111101111",
80840=>"101110101",
80841=>"000001111",
80842=>"000100110",
80843=>"000101111",
80844=>"000000111",
80845=>"101100100",
80846=>"000000000",
80847=>"110110111",
80848=>"000000100",
80849=>"001111100",
80850=>"111111001",
80851=>"011001000",
80852=>"000101111",
80853=>"001011000",
80854=>"111000111",
80855=>"111000000",
80856=>"000000100",
80857=>"000111000",
80858=>"111111011",
80859=>"000111010",
80860=>"011111111",
80861=>"111111111",
80862=>"010001100",
80863=>"000111010",
80864=>"000110111",
80865=>"111001101",
80866=>"111000000",
80867=>"011011011",
80868=>"000000000",
80869=>"011011111",
80870=>"111000001",
80871=>"000011000",
80872=>"010111110",
80873=>"000100101",
80874=>"000000110",
80875=>"000101010",
80876=>"000000000",
80877=>"000000111",
80878=>"000000010",
80879=>"101000000",
80880=>"111111111",
80881=>"111110100",
80882=>"101000110",
80883=>"000011000",
80884=>"001101011",
80885=>"000000000",
80886=>"100100110",
80887=>"111111000",
80888=>"111000000",
80889=>"001001000",
80890=>"111100100",
80891=>"111011100",
80892=>"101111010",
80893=>"000000000",
80894=>"000011000",
80895=>"111000111",
80896=>"111011001",
80897=>"011011000",
80898=>"000000000",
80899=>"011011011",
80900=>"100100000",
80901=>"100111111",
80902=>"001111000",
80903=>"000011111",
80904=>"100110110",
80905=>"000001011",
80906=>"001001000",
80907=>"101110110",
80908=>"111101111",
80909=>"000000000",
80910=>"111111110",
80911=>"110110101",
80912=>"100000001",
80913=>"110111011",
80914=>"000000000",
80915=>"011001001",
80916=>"111111001",
80917=>"000000000",
80918=>"111101001",
80919=>"111111111",
80920=>"000001101",
80921=>"100000001",
80922=>"110111001",
80923=>"000010001",
80924=>"000100000",
80925=>"111010011",
80926=>"111100000",
80927=>"000100100",
80928=>"101111001",
80929=>"111010011",
80930=>"110101010",
80931=>"101101001",
80932=>"101101001",
80933=>"000000000",
80934=>"000011011",
80935=>"101111111",
80936=>"101110100",
80937=>"010001001",
80938=>"000000000",
80939=>"110111101",
80940=>"100011000",
80941=>"110001011",
80942=>"111010011",
80943=>"101110000",
80944=>"011001111",
80945=>"111111100",
80946=>"110000101",
80947=>"110010000",
80948=>"111110011",
80949=>"111001010",
80950=>"111011111",
80951=>"101011111",
80952=>"100001111",
80953=>"000001111",
80954=>"001101111",
80955=>"111000010",
80956=>"000101100",
80957=>"110110110",
80958=>"000000000",
80959=>"101111000",
80960=>"000010111",
80961=>"000000010",
80962=>"111101000",
80963=>"001001001",
80964=>"001110110",
80965=>"111000101",
80966=>"001010000",
80967=>"110100110",
80968=>"011001101",
80969=>"100000011",
80970=>"001001111",
80971=>"110110010",
80972=>"100010000",
80973=>"111001001",
80974=>"111111100",
80975=>"011110111",
80976=>"010110110",
80977=>"100110111",
80978=>"111010001",
80979=>"011001100",
80980=>"000010010",
80981=>"101100000",
80982=>"011101101",
80983=>"000000001",
80984=>"000100010",
80985=>"001001000",
80986=>"001111111",
80987=>"011011010",
80988=>"000011111",
80989=>"000000101",
80990=>"111011111",
80991=>"111110011",
80992=>"000111110",
80993=>"000011000",
80994=>"001111011",
80995=>"001000000",
80996=>"000101101",
80997=>"011001000",
80998=>"111111111",
80999=>"000101110",
81000=>"111000011",
81001=>"111001011",
81002=>"110111111",
81003=>"111110111",
81004=>"000100101",
81005=>"100000100",
81006=>"001011011",
81007=>"111111110",
81008=>"001101101",
81009=>"111111111",
81010=>"011001000",
81011=>"111100000",
81012=>"100000000",
81013=>"111000001",
81014=>"110000010",
81015=>"111000000",
81016=>"000000000",
81017=>"000001010",
81018=>"110010000",
81019=>"000000000",
81020=>"110101101",
81021=>"100000001",
81022=>"101111111",
81023=>"000000000",
81024=>"110000000",
81025=>"010011000",
81026=>"110000001",
81027=>"111110110",
81028=>"101111111",
81029=>"101010110",
81030=>"011100101",
81031=>"000110000",
81032=>"001001001",
81033=>"000000000",
81034=>"000000001",
81035=>"111000111",
81036=>"000110100",
81037=>"101110010",
81038=>"101111111",
81039=>"100100110",
81040=>"000100100",
81041=>"101000110",
81042=>"000010001",
81043=>"001100111",
81044=>"011011010",
81045=>"100001011",
81046=>"010010010",
81047=>"011101110",
81048=>"110100010",
81049=>"000010100",
81050=>"000110000",
81051=>"000001111",
81052=>"111011000",
81053=>"000100010",
81054=>"110110011",
81055=>"000000000",
81056=>"000011111",
81057=>"010001000",
81058=>"110000001",
81059=>"110000110",
81060=>"111001110",
81061=>"000110111",
81062=>"110000001",
81063=>"000100000",
81064=>"100000000",
81065=>"010011111",
81066=>"001100100",
81067=>"010001111",
81068=>"111100000",
81069=>"111110111",
81070=>"000000000",
81071=>"001001111",
81072=>"100000001",
81073=>"011011110",
81074=>"010010100",
81075=>"101100110",
81076=>"101111111",
81077=>"011001110",
81078=>"111000001",
81079=>"100100100",
81080=>"110000000",
81081=>"000000000",
81082=>"000100000",
81083=>"111111100",
81084=>"101000001",
81085=>"111110100",
81086=>"110000011",
81087=>"000001000",
81088=>"111110000",
81089=>"000000100",
81090=>"111101101",
81091=>"011001100",
81092=>"001001001",
81093=>"100110000",
81094=>"000000111",
81095=>"011101101",
81096=>"100100000",
81097=>"000010010",
81098=>"111001111",
81099=>"000000010",
81100=>"010011000",
81101=>"000100111",
81102=>"011111111",
81103=>"001001111",
81104=>"010010110",
81105=>"101111111",
81106=>"000100110",
81107=>"010111101",
81108=>"100110100",
81109=>"000100101",
81110=>"100000001",
81111=>"110100011",
81112=>"011011000",
81113=>"000000111",
81114=>"011101001",
81115=>"000000000",
81116=>"111111111",
81117=>"000000000",
81118=>"110010111",
81119=>"000000110",
81120=>"000000111",
81121=>"111111101",
81122=>"111111000",
81123=>"001011110",
81124=>"000010000",
81125=>"100101011",
81126=>"110111111",
81127=>"111111111",
81128=>"011011011",
81129=>"010001101",
81130=>"111111111",
81131=>"110100001",
81132=>"011001111",
81133=>"111111001",
81134=>"100001000",
81135=>"100001001",
81136=>"000001000",
81137=>"110011100",
81138=>"001001000",
81139=>"001101001",
81140=>"000000000",
81141=>"001111101",
81142=>"000000001",
81143=>"001110110",
81144=>"001011001",
81145=>"111111111",
81146=>"111111111",
81147=>"111110111",
81148=>"010010000",
81149=>"010010000",
81150=>"010110100",
81151=>"010111000",
81152=>"000110011",
81153=>"000000010",
81154=>"111000000",
81155=>"011000101",
81156=>"100110110",
81157=>"111000000",
81158=>"000010010",
81159=>"101110111",
81160=>"000011111",
81161=>"000110011",
81162=>"110001001",
81163=>"111001111",
81164=>"101101101",
81165=>"000110111",
81166=>"101000000",
81167=>"100000101",
81168=>"111000010",
81169=>"101000010",
81170=>"000111101",
81171=>"100111011",
81172=>"101000000",
81173=>"111100100",
81174=>"011011011",
81175=>"000111011",
81176=>"111000001",
81177=>"111101101",
81178=>"010100100",
81179=>"010100111",
81180=>"000000100",
81181=>"111100111",
81182=>"111011111",
81183=>"101110100",
81184=>"100000000",
81185=>"000010111",
81186=>"010111000",
81187=>"100110010",
81188=>"000110100",
81189=>"011011001",
81190=>"000000110",
81191=>"000000100",
81192=>"111001111",
81193=>"110011010",
81194=>"110100111",
81195=>"011111001",
81196=>"000110010",
81197=>"101000100",
81198=>"010001100",
81199=>"111010101",
81200=>"101011000",
81201=>"110010011",
81202=>"110011111",
81203=>"100001100",
81204=>"011000100",
81205=>"101010111",
81206=>"000011011",
81207=>"000011111",
81208=>"111011100",
81209=>"000101111",
81210=>"100000100",
81211=>"100011101",
81212=>"001111001",
81213=>"111111011",
81214=>"010000100",
81215=>"000001111",
81216=>"111111100",
81217=>"010111010",
81218=>"000000000",
81219=>"111101100",
81220=>"100010011",
81221=>"000000100",
81222=>"000001111",
81223=>"111101000",
81224=>"000100001",
81225=>"101101101",
81226=>"010000000",
81227=>"111101101",
81228=>"110100110",
81229=>"011111100",
81230=>"010000100",
81231=>"100101011",
81232=>"100101100",
81233=>"111111111",
81234=>"111011010",
81235=>"110011001",
81236=>"111100000",
81237=>"000000101",
81238=>"000111110",
81239=>"000000000",
81240=>"111101111",
81241=>"000011011",
81242=>"110110010",
81243=>"000001000",
81244=>"100111111",
81245=>"010000000",
81246=>"010111010",
81247=>"111100000",
81248=>"000001111",
81249=>"001101101",
81250=>"011000100",
81251=>"100001001",
81252=>"000000000",
81253=>"000111011",
81254=>"101000101",
81255=>"110100000",
81256=>"000011011",
81257=>"011111100",
81258=>"000001010",
81259=>"111101010",
81260=>"100111011",
81261=>"111100000",
81262=>"000000100",
81263=>"000000000",
81264=>"001010100",
81265=>"100000010",
81266=>"000011010",
81267=>"111101101",
81268=>"011111100",
81269=>"110000100",
81270=>"000001110",
81271=>"111111111",
81272=>"000100000",
81273=>"000110111",
81274=>"111101000",
81275=>"101101111",
81276=>"001110100",
81277=>"000110100",
81278=>"110011000",
81279=>"111000000",
81280=>"000011011",
81281=>"111111000",
81282=>"100100011",
81283=>"111000111",
81284=>"101111000",
81285=>"001010000",
81286=>"100110010",
81287=>"000000000",
81288=>"101011000",
81289=>"111000000",
81290=>"011000001",
81291=>"100100100",
81292=>"000000101",
81293=>"111000111",
81294=>"000000111",
81295=>"011000001",
81296=>"111011101",
81297=>"000011111",
81298=>"100000011",
81299=>"000000000",
81300=>"000000000",
81301=>"001101111",
81302=>"101110000",
81303=>"000110011",
81304=>"100110111",
81305=>"011000010",
81306=>"111000100",
81307=>"111101100",
81308=>"000000011",
81309=>"011000101",
81310=>"111011100",
81311=>"111101101",
81312=>"000011111",
81313=>"111010010",
81314=>"101111010",
81315=>"011000111",
81316=>"011111010",
81317=>"000100111",
81318=>"011001101",
81319=>"000001010",
81320=>"000101111",
81321=>"010101101",
81322=>"101110100",
81323=>"010100100",
81324=>"001100001",
81325=>"000000000",
81326=>"000011111",
81327=>"111001100",
81328=>"101101001",
81329=>"111110100",
81330=>"111000011",
81331=>"000101000",
81332=>"110101111",
81333=>"100011001",
81334=>"000101100",
81335=>"111111000",
81336=>"000101100",
81337=>"011101000",
81338=>"000010000",
81339=>"000111000",
81340=>"110000000",
81341=>"111000000",
81342=>"000110111",
81343=>"111000010",
81344=>"111100000",
81345=>"000100100",
81346=>"111111100",
81347=>"110011001",
81348=>"000000101",
81349=>"111100000",
81350=>"001010010",
81351=>"000000000",
81352=>"000010111",
81353=>"011000000",
81354=>"101011111",
81355=>"000110011",
81356=>"000011011",
81357=>"110011001",
81358=>"010000010",
81359=>"000000100",
81360=>"111011110",
81361=>"000111111",
81362=>"111000100",
81363=>"000111111",
81364=>"110000111",
81365=>"011101000",
81366=>"110100000",
81367=>"111110110",
81368=>"000011000",
81369=>"110000111",
81370=>"000010111",
81371=>"111000100",
81372=>"110000101",
81373=>"111101101",
81374=>"111110101",
81375=>"101011000",
81376=>"111000000",
81377=>"111100000",
81378=>"111110100",
81379=>"111010000",
81380=>"111101000",
81381=>"011011011",
81382=>"000001101",
81383=>"000110110",
81384=>"011001111",
81385=>"101101000",
81386=>"001100100",
81387=>"111101100",
81388=>"111100110",
81389=>"110111000",
81390=>"000000001",
81391=>"100000001",
81392=>"000010111",
81393=>"011001000",
81394=>"000100000",
81395=>"000010111",
81396=>"000011010",
81397=>"111001000",
81398=>"110100010",
81399=>"111000000",
81400=>"000010011",
81401=>"000000000",
81402=>"111100111",
81403=>"000000000",
81404=>"100111010",
81405=>"111000111",
81406=>"000011001",
81407=>"110000001",
81408=>"010111001",
81409=>"100000010",
81410=>"000110010",
81411=>"100000010",
81412=>"011111110",
81413=>"100000110",
81414=>"001101111",
81415=>"100101011",
81416=>"000111111",
81417=>"000000000",
81418=>"011001110",
81419=>"111111111",
81420=>"111010000",
81421=>"100010111",
81422=>"111100001",
81423=>"100000000",
81424=>"000111111",
81425=>"000000011",
81426=>"000000000",
81427=>"000000111",
81428=>"101011111",
81429=>"110111101",
81430=>"000100011",
81431=>"000010111",
81432=>"000000000",
81433=>"111110000",
81434=>"111111111",
81435=>"000111111",
81436=>"111000111",
81437=>"101010010",
81438=>"111111110",
81439=>"011101000",
81440=>"000000000",
81441=>"111111011",
81442=>"111010111",
81443=>"010000010",
81444=>"011101111",
81445=>"000001101",
81446=>"000000000",
81447=>"100111110",
81448=>"111101111",
81449=>"000111000",
81450=>"000111111",
81451=>"001101000",
81452=>"111110001",
81453=>"111010000",
81454=>"101000001",
81455=>"001000001",
81456=>"000000000",
81457=>"001000000",
81458=>"010111101",
81459=>"111010010",
81460=>"000000100",
81461=>"011000000",
81462=>"110000011",
81463=>"000000010",
81464=>"001001001",
81465=>"001111101",
81466=>"100000000",
81467=>"010000000",
81468=>"011011001",
81469=>"111101101",
81470=>"000000110",
81471=>"000101101",
81472=>"111000110",
81473=>"111111101",
81474=>"000101101",
81475=>"001001110",
81476=>"000111010",
81477=>"000000100",
81478=>"000001101",
81479=>"111000111",
81480=>"111100110",
81481=>"111011100",
81482=>"101101111",
81483=>"101010111",
81484=>"000000111",
81485=>"001011111",
81486=>"110111000",
81487=>"101010111",
81488=>"101000000",
81489=>"000111111",
81490=>"010000110",
81491=>"001000011",
81492=>"110111111",
81493=>"000100111",
81494=>"111001001",
81495=>"011010000",
81496=>"010001010",
81497=>"011110001",
81498=>"110100100",
81499=>"001001010",
81500=>"110011000",
81501=>"000000001",
81502=>"010011111",
81503=>"100010111",
81504=>"000011010",
81505=>"101111110",
81506=>"000000000",
81507=>"111101011",
81508=>"110101100",
81509=>"111011000",
81510=>"110000000",
81511=>"000000000",
81512=>"111111000",
81513=>"000111111",
81514=>"000000111",
81515=>"111001111",
81516=>"111001111",
81517=>"010010001",
81518=>"111000010",
81519=>"000000010",
81520=>"110110100",
81521=>"001101101",
81522=>"001000100",
81523=>"111100000",
81524=>"000000111",
81525=>"001000001",
81526=>"111111000",
81527=>"010000101",
81528=>"001111111",
81529=>"010000000",
81530=>"110111111",
81531=>"000001110",
81532=>"001001100",
81533=>"100100100",
81534=>"000111011",
81535=>"111000000",
81536=>"000000111",
81537=>"000000000",
81538=>"000010111",
81539=>"000000111",
81540=>"010000000",
81541=>"100111110",
81542=>"001101101",
81543=>"010011001",
81544=>"011011001",
81545=>"000000001",
81546=>"111000100",
81547=>"001010111",
81548=>"000111111",
81549=>"000000010",
81550=>"000111111",
81551=>"101000110",
81552=>"110100100",
81553=>"111101111",
81554=>"000010111",
81555=>"100000010",
81556=>"111000101",
81557=>"000010111",
81558=>"001111011",
81559=>"000001001",
81560=>"111111111",
81561=>"000000110",
81562=>"000000100",
81563=>"000000100",
81564=>"000001001",
81565=>"010010111",
81566=>"000100001",
81567=>"101000000",
81568=>"101111111",
81569=>"100100000",
81570=>"001111111",
81571=>"000011111",
81572=>"010000100",
81573=>"100000000",
81574=>"111000110",
81575=>"010111111",
81576=>"100010111",
81577=>"000000000",
81578=>"100110110",
81579=>"000000000",
81580=>"110000100",
81581=>"111111000",
81582=>"111101000",
81583=>"111000000",
81584=>"111011010",
81585=>"011111011",
81586=>"000010101",
81587=>"000001110",
81588=>"111101101",
81589=>"100100101",
81590=>"000000000",
81591=>"010110101",
81592=>"100110100",
81593=>"111001000",
81594=>"011000111",
81595=>"101000000",
81596=>"101111101",
81597=>"000111101",
81598=>"110011100",
81599=>"000000001",
81600=>"111000000",
81601=>"001001000",
81602=>"111000010",
81603=>"011000001",
81604=>"010010000",
81605=>"110000101",
81606=>"100000001",
81607=>"011000111",
81608=>"000111111",
81609=>"000000101",
81610=>"000001101",
81611=>"000010000",
81612=>"000000001",
81613=>"100101001",
81614=>"000000010",
81615=>"010010000",
81616=>"000111011",
81617=>"111101110",
81618=>"000000010",
81619=>"011011001",
81620=>"111000010",
81621=>"001111100",
81622=>"000111000",
81623=>"000100000",
81624=>"100000000",
81625=>"110010000",
81626=>"100101101",
81627=>"000000110",
81628=>"001011111",
81629=>"000011000",
81630=>"111011000",
81631=>"000000000",
81632=>"000011001",
81633=>"111010100",
81634=>"000011010",
81635=>"111111000",
81636=>"111000000",
81637=>"101101100",
81638=>"100110000",
81639=>"111011011",
81640=>"111010101",
81641=>"000100111",
81642=>"100100010",
81643=>"001010000",
81644=>"000001000",
81645=>"000111111",
81646=>"001000000",
81647=>"101000101",
81648=>"000000010",
81649=>"011000101",
81650=>"111000000",
81651=>"011011001",
81652=>"110110110",
81653=>"100001101",
81654=>"000000000",
81655=>"111111111",
81656=>"000111011",
81657=>"000000000",
81658=>"000101101",
81659=>"111001001",
81660=>"000111111",
81661=>"000000110",
81662=>"100101111",
81663=>"101001100",
81664=>"011010100",
81665=>"110010110",
81666=>"101000001",
81667=>"111000000",
81668=>"100000000",
81669=>"110111001",
81670=>"100010111",
81671=>"010111111",
81672=>"000000000",
81673=>"001000110",
81674=>"001110110",
81675=>"111111000",
81676=>"010100000",
81677=>"111110110",
81678=>"111111100",
81679=>"111110111",
81680=>"001000000",
81681=>"000000100",
81682=>"111101111",
81683=>"011010100",
81684=>"101111000",
81685=>"111111000",
81686=>"001000000",
81687=>"000000101",
81688=>"000000101",
81689=>"111111001",
81690=>"111101000",
81691=>"011000000",
81692=>"110000000",
81693=>"101110111",
81694=>"010000111",
81695=>"000110000",
81696=>"111101000",
81697=>"001011000",
81698=>"000000111",
81699=>"010010010",
81700=>"100101000",
81701=>"110000010",
81702=>"111001110",
81703=>"000000111",
81704=>"011110010",
81705=>"001011011",
81706=>"111001001",
81707=>"111100010",
81708=>"111111011",
81709=>"111110000",
81710=>"110011101",
81711=>"000000011",
81712=>"110001000",
81713=>"001001101",
81714=>"000000000",
81715=>"010000010",
81716=>"000111111",
81717=>"010110110",
81718=>"100100111",
81719=>"111100000",
81720=>"001000001",
81721=>"111101001",
81722=>"100101000",
81723=>"000000000",
81724=>"101000000",
81725=>"010101111",
81726=>"100000000",
81727=>"111100100",
81728=>"001000000",
81729=>"111000000",
81730=>"111111000",
81731=>"001111010",
81732=>"110100000",
81733=>"000000101",
81734=>"110010111",
81735=>"000111111",
81736=>"001011111",
81737=>"000111111",
81738=>"101101000",
81739=>"111101111",
81740=>"111000111",
81741=>"011101001",
81742=>"100100101",
81743=>"000000101",
81744=>"000111110",
81745=>"110111111",
81746=>"111111010",
81747=>"011100010",
81748=>"110110000",
81749=>"001000000",
81750=>"101000110",
81751=>"000000000",
81752=>"111111110",
81753=>"000101111",
81754=>"101100111",
81755=>"000111111",
81756=>"110000100",
81757=>"001101000",
81758=>"111100000",
81759=>"101101111",
81760=>"111010000",
81761=>"000100010",
81762=>"100000000",
81763=>"001101110",
81764=>"111011000",
81765=>"111111110",
81766=>"111000001",
81767=>"101011111",
81768=>"000000000",
81769=>"001000000",
81770=>"010000000",
81771=>"111111111",
81772=>"001111111",
81773=>"110110000",
81774=>"010110100",
81775=>"011001111",
81776=>"001000001",
81777=>"000000001",
81778=>"001001011",
81779=>"000010000",
81780=>"111011011",
81781=>"000000101",
81782=>"101000000",
81783=>"010010010",
81784=>"111000101",
81785=>"110000000",
81786=>"111101000",
81787=>"000000110",
81788=>"100010110",
81789=>"000001001",
81790=>"000101111",
81791=>"100101011",
81792=>"000000000",
81793=>"100111101",
81794=>"110010000",
81795=>"101110111",
81796=>"000110111",
81797=>"101111111",
81798=>"011011111",
81799=>"101100000",
81800=>"100100000",
81801=>"000011111",
81802=>"111010010",
81803=>"101111000",
81804=>"110000000",
81805=>"000100110",
81806=>"111111101",
81807=>"100000000",
81808=>"100101101",
81809=>"111001010",
81810=>"010000000",
81811=>"011000000",
81812=>"100000000",
81813=>"110000000",
81814=>"010111000",
81815=>"110100100",
81816=>"010000110",
81817=>"100111010",
81818=>"001001100",
81819=>"000000000",
81820=>"111110100",
81821=>"000000100",
81822=>"010001101",
81823=>"101101000",
81824=>"001100100",
81825=>"000000010",
81826=>"000101101",
81827=>"000000000",
81828=>"110111011",
81829=>"110111001",
81830=>"001110001",
81831=>"111011111",
81832=>"011010000",
81833=>"111000000",
81834=>"111000000",
81835=>"000001111",
81836=>"000100000",
81837=>"100100000",
81838=>"100111110",
81839=>"000110101",
81840=>"101101101",
81841=>"101011001",
81842=>"000000100",
81843=>"000010011",
81844=>"000001100",
81845=>"000100100",
81846=>"111011011",
81847=>"010000101",
81848=>"101000000",
81849=>"110000000",
81850=>"010111001",
81851=>"011100010",
81852=>"010000010",
81853=>"111111111",
81854=>"011010000",
81855=>"000000011",
81856=>"000111100",
81857=>"011001001",
81858=>"110111010",
81859=>"011001000",
81860=>"111000100",
81861=>"110110101",
81862=>"110010111",
81863=>"000000000",
81864=>"111011101",
81865=>"111010000",
81866=>"111111111",
81867=>"111101100",
81868=>"010100110",
81869=>"001011011",
81870=>"000000111",
81871=>"000111010",
81872=>"110110111",
81873=>"110001001",
81874=>"111000001",
81875=>"110111011",
81876=>"111101001",
81877=>"101100010",
81878=>"111111000",
81879=>"100000010",
81880=>"010000000",
81881=>"111111010",
81882=>"100000111",
81883=>"000000111",
81884=>"000001000",
81885=>"111111000",
81886=>"011111101",
81887=>"000000000",
81888=>"101000101",
81889=>"001001111",
81890=>"010000011",
81891=>"111001101",
81892=>"111000000",
81893=>"001111010",
81894=>"111011010",
81895=>"111101100",
81896=>"111011010",
81897=>"000000110",
81898=>"000011011",
81899=>"111001000",
81900=>"000000010",
81901=>"000010110",
81902=>"111000010",
81903=>"000111111",
81904=>"010111010",
81905=>"001001001",
81906=>"111000010",
81907=>"000110111",
81908=>"110110001",
81909=>"000101111",
81910=>"000111110",
81911=>"000100111",
81912=>"010000100",
81913=>"000010111",
81914=>"111111111",
81915=>"111101000",
81916=>"000101111",
81917=>"111010000",
81918=>"001011000",
81919=>"000111111",
81920=>"001001111",
81921=>"000001000",
81922=>"011000100",
81923=>"000111000",
81924=>"111011111",
81925=>"001001000",
81926=>"000000011",
81927=>"111110111",
81928=>"101000111",
81929=>"000000001",
81930=>"110011011",
81931=>"000111101",
81932=>"111001000",
81933=>"111101100",
81934=>"110000100",
81935=>"000010010",
81936=>"111100011",
81937=>"111000011",
81938=>"110111100",
81939=>"001000001",
81940=>"000001101",
81941=>"011001000",
81942=>"000000100",
81943=>"001111110",
81944=>"100000110",
81945=>"000000000",
81946=>"000111111",
81947=>"000000100",
81948=>"000111010",
81949=>"000111100",
81950=>"101111101",
81951=>"000000000",
81952=>"000000000",
81953=>"100111111",
81954=>"010110001",
81955=>"000000000",
81956=>"110111100",
81957=>"000011010",
81958=>"000111110",
81959=>"110000111",
81960=>"000001000",
81961=>"001111111",
81962=>"000000010",
81963=>"000000100",
81964=>"100000111",
81965=>"111111111",
81966=>"000000111",
81967=>"110111110",
81968=>"101111110",
81969=>"111111100",
81970=>"011100010",
81971=>"000101101",
81972=>"111111000",
81973=>"001101111",
81974=>"000000101",
81975=>"111111110",
81976=>"000001100",
81977=>"000000111",
81978=>"001000000",
81979=>"000001000",
81980=>"001100011",
81981=>"111111011",
81982=>"101001001",
81983=>"111111100",
81984=>"001010011",
81985=>"111111100",
81986=>"110111001",
81987=>"101101111",
81988=>"000000111",
81989=>"101101101",
81990=>"000000011",
81991=>"110011011",
81992=>"100111111",
81993=>"100111111",
81994=>"000000000",
81995=>"000000000",
81996=>"111111111",
81997=>"111000010",
81998=>"111111001",
81999=>"111000000",
82000=>"111000000",
82001=>"111111000",
82002=>"101111000",
82003=>"000100101",
82004=>"000000111",
82005=>"010110110",
82006=>"110010000",
82007=>"000000110",
82008=>"000001100",
82009=>"111111110",
82010=>"110000101",
82011=>"111111011",
82012=>"110010111",
82013=>"000000001",
82014=>"100110000",
82015=>"001000110",
82016=>"000111011",
82017=>"000000001",
82018=>"011011001",
82019=>"111011000",
82020=>"000000001",
82021=>"010111101",
82022=>"000111111",
82023=>"000101000",
82024=>"000111111",
82025=>"111111111",
82026=>"000010111",
82027=>"101000101",
82028=>"111110111",
82029=>"111110010",
82030=>"101000001",
82031=>"000111111",
82032=>"111111111",
82033=>"110000110",
82034=>"000001100",
82035=>"111111011",
82036=>"111111000",
82037=>"001011001",
82038=>"110010001",
82039=>"000001000",
82040=>"000000111",
82041=>"000000111",
82042=>"111111011",
82043=>"101111100",
82044=>"011001001",
82045=>"000001011",
82046=>"000001000",
82047=>"001001001",
82048=>"000000100",
82049=>"000000011",
82050=>"100111111",
82051=>"111000000",
82052=>"111111000",
82053=>"100100110",
82054=>"000100110",
82055=>"111000000",
82056=>"110110000",
82057=>"000101111",
82058=>"000111000",
82059=>"111011000",
82060=>"000000110",
82061=>"001001001",
82062=>"000000000",
82063=>"000000000",
82064=>"111111000",
82065=>"100100000",
82066=>"000001010",
82067=>"000000010",
82068=>"111000000",
82069=>"000000111",
82070=>"111110000",
82071=>"100101100",
82072=>"111001000",
82073=>"001000000",
82074=>"000010010",
82075=>"010010000",
82076=>"010001101",
82077=>"000000000",
82078=>"000001101",
82079=>"000000111",
82080=>"111011100",
82081=>"111110000",
82082=>"000000111",
82083=>"111000000",
82084=>"100100000",
82085=>"111000000",
82086=>"000000011",
82087=>"000000111",
82088=>"001000011",
82089=>"110010000",
82090=>"111111011",
82091=>"001000000",
82092=>"111001110",
82093=>"111111100",
82094=>"010011011",
82095=>"111000001",
82096=>"100000000",
82097=>"111000110",
82098=>"000000001",
82099=>"111001001",
82100=>"111100100",
82101=>"000111110",
82102=>"011011010",
82103=>"100000010",
82104=>"000001110",
82105=>"110000010",
82106=>"000000000",
82107=>"000101111",
82108=>"101000000",
82109=>"010010100",
82110=>"111111011",
82111=>"111110101",
82112=>"000100111",
82113=>"100000110",
82114=>"101000010",
82115=>"101101000",
82116=>"000111111",
82117=>"011111111",
82118=>"100000000",
82119=>"000000111",
82120=>"111101110",
82121=>"001000000",
82122=>"101110000",
82123=>"110101100",
82124=>"011110110",
82125=>"100000100",
82126=>"110000000",
82127=>"000011000",
82128=>"010110110",
82129=>"111111001",
82130=>"000000101",
82131=>"110010011",
82132=>"111000001",
82133=>"111000011",
82134=>"000011111",
82135=>"000110111",
82136=>"000110111",
82137=>"000000001",
82138=>"111100011",
82139=>"111000000",
82140=>"000000100",
82141=>"111010000",
82142=>"000000000",
82143=>"101001000",
82144=>"111000100",
82145=>"111100001",
82146=>"101110010",
82147=>"011110110",
82148=>"111100000",
82149=>"111110101",
82150=>"000001110",
82151=>"000000100",
82152=>"101001000",
82153=>"000000100",
82154=>"101100110",
82155=>"000000001",
82156=>"000000100",
82157=>"111111001",
82158=>"111000000",
82159=>"000000000",
82160=>"000001111",
82161=>"100111111",
82162=>"101111101",
82163=>"111011011",
82164=>"000000001",
82165=>"111000000",
82166=>"111000000",
82167=>"111111001",
82168=>"000000111",
82169=>"111111111",
82170=>"000000000",
82171=>"000000000",
82172=>"111111000",
82173=>"000111111",
82174=>"111000001",
82175=>"111111110",
82176=>"110100000",
82177=>"000101101",
82178=>"111101100",
82179=>"010110000",
82180=>"111000110",
82181=>"110000000",
82182=>"010110010",
82183=>"011001110",
82184=>"010000100",
82185=>"111101100",
82186=>"010000000",
82187=>"000010011",
82188=>"111100000",
82189=>"000000011",
82190=>"110100100",
82191=>"110111100",
82192=>"000011011",
82193=>"010000000",
82194=>"011111000",
82195=>"010000000",
82196=>"110111101",
82197=>"111001100",
82198=>"001101111",
82199=>"010111101",
82200=>"010010000",
82201=>"000100111",
82202=>"000000000",
82203=>"000001111",
82204=>"001000000",
82205=>"010011010",
82206=>"001100010",
82207=>"111010001",
82208=>"101000010",
82209=>"000010011",
82210=>"111000100",
82211=>"000101000",
82212=>"000100111",
82213=>"011011111",
82214=>"111100100",
82215=>"000100110",
82216=>"010011011",
82217=>"011101100",
82218=>"000010100",
82219=>"000000000",
82220=>"100001011",
82221=>"110011110",
82222=>"000011101",
82223=>"101011100",
82224=>"111100000",
82225=>"011001011",
82226=>"000000000",
82227=>"111100000",
82228=>"010001101",
82229=>"111111111",
82230=>"001111111",
82231=>"111010100",
82232=>"010111000",
82233=>"011001100",
82234=>"011000100",
82235=>"001101100",
82236=>"010001011",
82237=>"010111100",
82238=>"000000000",
82239=>"001011111",
82240=>"001101011",
82241=>"000101111",
82242=>"111110111",
82243=>"100000000",
82244=>"111000000",
82245=>"111100000",
82246=>"010000111",
82247=>"010010000",
82248=>"000001110",
82249=>"000011011",
82250=>"000100000",
82251=>"111111011",
82252=>"111101101",
82253=>"110001101",
82254=>"100100111",
82255=>"001111100",
82256=>"100100111",
82257=>"010010111",
82258=>"101111111",
82259=>"000011000",
82260=>"111101101",
82261=>"111011011",
82262=>"000000000",
82263=>"000100000",
82264=>"000010110",
82265=>"001001101",
82266=>"110001001",
82267=>"100100110",
82268=>"010000111",
82269=>"010000001",
82270=>"111100000",
82271=>"100100100",
82272=>"000000010",
82273=>"000010011",
82274=>"001000100",
82275=>"001001101",
82276=>"011000000",
82277=>"010100011",
82278=>"000010011",
82279=>"111100100",
82280=>"001011011",
82281=>"111110111",
82282=>"001001010",
82283=>"111111111",
82284=>"110110000",
82285=>"111111101",
82286=>"000000000",
82287=>"010001001",
82288=>"000110110",
82289=>"000100010",
82290=>"011111110",
82291=>"000001000",
82292=>"010101110",
82293=>"111100100",
82294=>"011111010",
82295=>"000011010",
82296=>"110000100",
82297=>"111000100",
82298=>"011111010",
82299=>"011100100",
82300=>"011111100",
82301=>"011110000",
82302=>"000100000",
82303=>"001001000",
82304=>"111111000",
82305=>"000010000",
82306=>"010001000",
82307=>"111011111",
82308=>"101101110",
82309=>"111000000",
82310=>"100110100",
82311=>"000100111",
82312=>"000001001",
82313=>"001000000",
82314=>"000001011",
82315=>"100100000",
82316=>"110010000",
82317=>"111101100",
82318=>"001000000",
82319=>"000100000",
82320=>"111100111",
82321=>"011111111",
82322=>"011101100",
82323=>"000111111",
82324=>"000111111",
82325=>"111000000",
82326=>"101011110",
82327=>"010010100",
82328=>"000001011",
82329=>"111000001",
82330=>"000000111",
82331=>"000000000",
82332=>"110100100",
82333=>"000011011",
82334=>"111111000",
82335=>"100100000",
82336=>"001000100",
82337=>"010000000",
82338=>"101010100",
82339=>"011000000",
82340=>"111101101",
82341=>"010000001",
82342=>"011011001",
82343=>"000011111",
82344=>"010001101",
82345=>"000000000",
82346=>"111000100",
82347=>"000111010",
82348=>"111111011",
82349=>"010000000",
82350=>"110011111",
82351=>"011011011",
82352=>"000100001",
82353=>"000011000",
82354=>"011111111",
82355=>"000101000",
82356=>"000000110",
82357=>"111110111",
82358=>"011111011",
82359=>"111100000",
82360=>"001100011",
82361=>"001111111",
82362=>"000010011",
82363=>"000110010",
82364=>"111110000",
82365=>"010111111",
82366=>"010000000",
82367=>"011111001",
82368=>"000001000",
82369=>"010110100",
82370=>"000000100",
82371=>"011001000",
82372=>"000010010",
82373=>"110111011",
82374=>"111010100",
82375=>"001101101",
82376=>"000100010",
82377=>"010010010",
82378=>"101000101",
82379=>"000100111",
82380=>"000011011",
82381=>"100001011",
82382=>"111110110",
82383=>"110100000",
82384=>"000010010",
82385=>"110100101",
82386=>"000000010",
82387=>"011111111",
82388=>"000000011",
82389=>"011100100",
82390=>"011101000",
82391=>"100111000",
82392=>"000100100",
82393=>"001011111",
82394=>"010110100",
82395=>"110000000",
82396=>"110111101",
82397=>"110010001",
82398=>"011010101",
82399=>"000010010",
82400=>"111101001",
82401=>"111111101",
82402=>"111101101",
82403=>"000001001",
82404=>"100100000",
82405=>"011001100",
82406=>"100110100",
82407=>"010000000",
82408=>"000000111",
82409=>"110111010",
82410=>"000000000",
82411=>"111100000",
82412=>"010010011",
82413=>"111100000",
82414=>"000000000",
82415=>"111110000",
82416=>"001100100",
82417=>"001111100",
82418=>"010111100",
82419=>"000000100",
82420=>"010110101",
82421=>"101100100",
82422=>"100000000",
82423=>"110000100",
82424=>"000111111",
82425=>"101001100",
82426=>"111101111",
82427=>"100000101",
82428=>"101011001",
82429=>"000000010",
82430=>"011011101",
82431=>"000100000",
82432=>"000011011",
82433=>"011011111",
82434=>"101100000",
82435=>"000100010",
82436=>"000000100",
82437=>"111111100",
82438=>"100000110",
82439=>"001000011",
82440=>"000000011",
82441=>"000111111",
82442=>"101100000",
82443=>"010011001",
82444=>"000000110",
82445=>"000000000",
82446=>"101101001",
82447=>"000000011",
82448=>"011111111",
82449=>"010010011",
82450=>"110100000",
82451=>"011100000",
82452=>"101111110",
82453=>"000011010",
82454=>"100100100",
82455=>"111111110",
82456=>"000000011",
82457=>"010111101",
82458=>"010111100",
82459=>"010010110",
82460=>"111100100",
82461=>"000100100",
82462=>"111010000",
82463=>"000111111",
82464=>"000110000",
82465=>"011111011",
82466=>"100010011",
82467=>"000101111",
82468=>"010011001",
82469=>"001101100",
82470=>"000000000",
82471=>"100001000",
82472=>"001111101",
82473=>"001111011",
82474=>"100000000",
82475=>"000000000",
82476=>"000001001",
82477=>"011000011",
82478=>"110000100",
82479=>"001110100",
82480=>"100101111",
82481=>"001011111",
82482=>"111011011",
82483=>"100100100",
82484=>"111000000",
82485=>"101000001",
82486=>"110100001",
82487=>"000000010",
82488=>"111000110",
82489=>"111101000",
82490=>"111100100",
82491=>"111101101",
82492=>"011010001",
82493=>"111111110",
82494=>"000000110",
82495=>"001111111",
82496=>"000111010",
82497=>"011111100",
82498=>"000000110",
82499=>"111011001",
82500=>"111100010",
82501=>"001010011",
82502=>"101000000",
82503=>"111111000",
82504=>"010110111",
82505=>"001011011",
82506=>"101000000",
82507=>"011100001",
82508=>"111111000",
82509=>"001110100",
82510=>"000110111",
82511=>"111101111",
82512=>"101111000",
82513=>"110111101",
82514=>"000100010",
82515=>"011001000",
82516=>"111000000",
82517=>"110110111",
82518=>"011011001",
82519=>"010001111",
82520=>"111101001",
82521=>"001110001",
82522=>"000111111",
82523=>"010111111",
82524=>"000000000",
82525=>"110001001",
82526=>"111111100",
82527=>"111100000",
82528=>"000011111",
82529=>"111111101",
82530=>"111100111",
82531=>"100000000",
82532=>"111111111",
82533=>"111110110",
82534=>"111110111",
82535=>"000000111",
82536=>"101000010",
82537=>"011010000",
82538=>"010000111",
82539=>"111111000",
82540=>"111111111",
82541=>"000000010",
82542=>"000111010",
82543=>"011010111",
82544=>"101111001",
82545=>"000100110",
82546=>"111001000",
82547=>"000011001",
82548=>"000001001",
82549=>"110000000",
82550=>"000000000",
82551=>"000001000",
82552=>"000000000",
82553=>"111011100",
82554=>"110111111",
82555=>"000000100",
82556=>"000110111",
82557=>"011110000",
82558=>"000000000",
82559=>"111000101",
82560=>"000010100",
82561=>"111100000",
82562=>"001111111",
82563=>"000000011",
82564=>"011011011",
82565=>"111111100",
82566=>"100011001",
82567=>"000000001",
82568=>"101100100",
82569=>"001000000",
82570=>"000000001",
82571=>"011011000",
82572=>"000100111",
82573=>"000000000",
82574=>"100000000",
82575=>"100000101",
82576=>"111111001",
82577=>"100111101",
82578=>"101000001",
82579=>"110000000",
82580=>"001010011",
82581=>"111000010",
82582=>"111111111",
82583=>"000011011",
82584=>"011011111",
82585=>"000000111",
82586=>"111000100",
82587=>"000100110",
82588=>"111100100",
82589=>"010111011",
82590=>"100000100",
82591=>"111000000",
82592=>"001000001",
82593=>"110000010",
82594=>"100010110",
82595=>"000000111",
82596=>"011011001",
82597=>"100011111",
82598=>"001110111",
82599=>"010111111",
82600=>"111011111",
82601=>"000010011",
82602=>"101110110",
82603=>"111100100",
82604=>"010000000",
82605=>"001001001",
82606=>"001100100",
82607=>"000000011",
82608=>"100011111",
82609=>"000011001",
82610=>"111111111",
82611=>"000010010",
82612=>"010111011",
82613=>"000000011",
82614=>"000111011",
82615=>"001000000",
82616=>"110101011",
82617=>"100000110",
82618=>"111111001",
82619=>"101111010",
82620=>"010110010",
82621=>"111111111",
82622=>"000110011",
82623=>"101001111",
82624=>"111100100",
82625=>"111101110",
82626=>"111101111",
82627=>"000110010",
82628=>"101101000",
82629=>"011000101",
82630=>"110100000",
82631=>"000100000",
82632=>"000010010",
82633=>"000100001",
82634=>"000011111",
82635=>"000011011",
82636=>"100101111",
82637=>"100001011",
82638=>"100100110",
82639=>"010111000",
82640=>"000100000",
82641=>"000110000",
82642=>"000011011",
82643=>"001011001",
82644=>"011100100",
82645=>"010110110",
82646=>"100000010",
82647=>"000011011",
82648=>"001011000",
82649=>"111000101",
82650=>"100100100",
82651=>"100000000",
82652=>"001111011",
82653=>"010011111",
82654=>"101111111",
82655=>"111010000",
82656=>"101000100",
82657=>"101100100",
82658=>"000000000",
82659=>"000000110",
82660=>"101000000",
82661=>"000000000",
82662=>"000001000",
82663=>"000001001",
82664=>"000000010",
82665=>"000001010",
82666=>"111001000",
82667=>"000000001",
82668=>"000000111",
82669=>"000000001",
82670=>"000100000",
82671=>"000101010",
82672=>"111111000",
82673=>"010100101",
82674=>"010010011",
82675=>"000111011",
82676=>"100110100",
82677=>"000000101",
82678=>"010000010",
82679=>"000111011",
82680=>"111010010",
82681=>"100111111",
82682=>"000000000",
82683=>"011101101",
82684=>"101000010",
82685=>"100111011",
82686=>"000000001",
82687=>"101000000",
82688=>"011001000",
82689=>"010000111",
82690=>"010011010",
82691=>"101000000",
82692=>"111110111",
82693=>"000001000",
82694=>"110100010",
82695=>"000000111",
82696=>"111111111",
82697=>"001000000",
82698=>"110110110",
82699=>"001101001",
82700=>"101101101",
82701=>"000001000",
82702=>"001011011",
82703=>"111110010",
82704=>"111111001",
82705=>"110000000",
82706=>"110000000",
82707=>"000000111",
82708=>"110000100",
82709=>"111100100",
82710=>"011011101",
82711=>"110111111",
82712=>"100100110",
82713=>"001001101",
82714=>"101101101",
82715=>"111010010",
82716=>"000000000",
82717=>"000000010",
82718=>"000000000",
82719=>"101001101",
82720=>"100101111",
82721=>"111111011",
82722=>"010110110",
82723=>"110000110",
82724=>"110110100",
82725=>"011011111",
82726=>"010000000",
82727=>"111111111",
82728=>"111111011",
82729=>"011011001",
82730=>"000000111",
82731=>"101000100",
82732=>"010111011",
82733=>"000000000",
82734=>"000000000",
82735=>"000100000",
82736=>"000000100",
82737=>"111111011",
82738=>"000000100",
82739=>"000000000",
82740=>"011110110",
82741=>"101011110",
82742=>"111111111",
82743=>"000100011",
82744=>"000000000",
82745=>"000000111",
82746=>"000010100",
82747=>"111000000",
82748=>"000000001",
82749=>"011101001",
82750=>"100100100",
82751=>"111111111",
82752=>"000000000",
82753=>"101111111",
82754=>"000100000",
82755=>"010001001",
82756=>"000000110",
82757=>"001101101",
82758=>"100101100",
82759=>"001001001",
82760=>"000000000",
82761=>"101101101",
82762=>"101101100",
82763=>"101011101",
82764=>"000000000",
82765=>"111111111",
82766=>"111111011",
82767=>"111101110",
82768=>"001101000",
82769=>"111001000",
82770=>"000000100",
82771=>"011000010",
82772=>"010111111",
82773=>"100100100",
82774=>"111111001",
82775=>"000100100",
82776=>"101111111",
82777=>"001011111",
82778=>"111111110",
82779=>"001000101",
82780=>"101000111",
82781=>"011011011",
82782=>"010111011",
82783=>"000100100",
82784=>"111111111",
82785=>"101000101",
82786=>"100000000",
82787=>"111111011",
82788=>"101111110",
82789=>"111111111",
82790=>"111111100",
82791=>"011000111",
82792=>"000000000",
82793=>"000000011",
82794=>"000000001",
82795=>"010011001",
82796=>"010101001",
82797=>"111011011",
82798=>"111000000",
82799=>"000000000",
82800=>"100100100",
82801=>"000000010",
82802=>"111011111",
82803=>"011111010",
82804=>"000000000",
82805=>"000101101",
82806=>"000000000",
82807=>"011111000",
82808=>"000010011",
82809=>"000000000",
82810=>"000011010",
82811=>"111111111",
82812=>"001000110",
82813=>"110110110",
82814=>"111000000",
82815=>"010111010",
82816=>"000000000",
82817=>"000000100",
82818=>"000000000",
82819=>"000000000",
82820=>"000000000",
82821=>"000000100",
82822=>"110110110",
82823=>"011011011",
82824=>"011011001",
82825=>"010011010",
82826=>"011011010",
82827=>"110100100",
82828=>"101111011",
82829=>"111101110",
82830=>"101001110",
82831=>"101101100",
82832=>"111110110",
82833=>"111111110",
82834=>"001010000",
82835=>"000000000",
82836=>"101110110",
82837=>"110100101",
82838=>"110111011",
82839=>"001101111",
82840=>"000100111",
82841=>"000000111",
82842=>"000010011",
82843=>"000000000",
82844=>"000000000",
82845=>"000000010",
82846=>"000000000",
82847=>"110011000",
82848=>"011111011",
82849=>"000000000",
82850=>"111011000",
82851=>"000000000",
82852=>"000000000",
82853=>"110101110",
82854=>"101011111",
82855=>"111111111",
82856=>"000000001",
82857=>"000001010",
82858=>"000001111",
82859=>"000000000",
82860=>"111111111",
82861=>"000000000",
82862=>"110101010",
82863=>"101101100",
82864=>"000000100",
82865=>"000001111",
82866=>"111010111",
82867=>"100000100",
82868=>"111111111",
82869=>"011010000",
82870=>"000100100",
82871=>"011000000",
82872=>"000000100",
82873=>"001111010",
82874=>"000000000",
82875=>"000000000",
82876=>"111101010",
82877=>"000110111",
82878=>"110100110",
82879=>"000000000",
82880=>"111100110",
82881=>"000000101",
82882=>"000100001",
82883=>"001001011",
82884=>"000000000",
82885=>"100000001",
82886=>"000000101",
82887=>"000000111",
82888=>"111111111",
82889=>"010010000",
82890=>"101101110",
82891=>"111111110",
82892=>"001000000",
82893=>"110100111",
82894=>"111111001",
82895=>"000000000",
82896=>"010010000",
82897=>"111111111",
82898=>"010010010",
82899=>"111110100",
82900=>"001000101",
82901=>"111111111",
82902=>"010111010",
82903=>"000000000",
82904=>"111111111",
82905=>"111011011",
82906=>"110111111",
82907=>"010011000",
82908=>"000000000",
82909=>"000001000",
82910=>"011100101",
82911=>"000000000",
82912=>"010010000",
82913=>"000000000",
82914=>"100011011",
82915=>"111100001",
82916=>"001000101",
82917=>"001100111",
82918=>"000010000",
82919=>"010001111",
82920=>"001000000",
82921=>"111111111",
82922=>"011111101",
82923=>"111111100",
82924=>"100111000",
82925=>"000000000",
82926=>"100000000",
82927=>"100101111",
82928=>"010010010",
82929=>"101000001",
82930=>"000110000",
82931=>"111111111",
82932=>"110000001",
82933=>"111111111",
82934=>"001001000",
82935=>"000000000",
82936=>"111111111",
82937=>"000000000",
82938=>"111000101",
82939=>"111111010",
82940=>"111001011",
82941=>"111010111",
82942=>"111101110",
82943=>"011110000",
82944=>"011111001",
82945=>"001000000",
82946=>"111101100",
82947=>"010000000",
82948=>"000111011",
82949=>"000000000",
82950=>"111000101",
82951=>"101101110",
82952=>"010010011",
82953=>"000000000",
82954=>"111001111",
82955=>"000011111",
82956=>"000101010",
82957=>"010001000",
82958=>"000111111",
82959=>"111111000",
82960=>"010100000",
82961=>"000100101",
82962=>"000000100",
82963=>"000010010",
82964=>"101000000",
82965=>"101100000",
82966=>"111111000",
82967=>"111110111",
82968=>"000000000",
82969=>"101001111",
82970=>"111110011",
82971=>"110000000",
82972=>"011000000",
82973=>"001101001",
82974=>"011010000",
82975=>"000000111",
82976=>"110101001",
82977=>"100101010",
82978=>"000000110",
82979=>"000111111",
82980=>"111101101",
82981=>"011111110",
82982=>"100000010",
82983=>"101000000",
82984=>"111000111",
82985=>"101010000",
82986=>"001010000",
82987=>"101100000",
82988=>"001011001",
82989=>"110000011",
82990=>"001011000",
82991=>"010111101",
82992=>"001111100",
82993=>"000111011",
82994=>"011000111",
82995=>"000000000",
82996=>"000110000",
82997=>"100111111",
82998=>"011110000",
82999=>"010111111",
83000=>"111101111",
83001=>"111101001",
83002=>"100101110",
83003=>"001010010",
83004=>"000011111",
83005=>"100011111",
83006=>"011101000",
83007=>"110011011",
83008=>"100111111",
83009=>"001111111",
83010=>"000000101",
83011=>"110000110",
83012=>"010010000",
83013=>"101101010",
83014=>"100100000",
83015=>"010001111",
83016=>"110110110",
83017=>"000111111",
83018=>"101100100",
83019=>"111100100",
83020=>"000110000",
83021=>"111101100",
83022=>"000010110",
83023=>"011111101",
83024=>"111100000",
83025=>"010010000",
83026=>"000010011",
83027=>"000011011",
83028=>"000000111",
83029=>"010010000",
83030=>"010011011",
83031=>"100001101",
83032=>"000001111",
83033=>"100100011",
83034=>"111110100",
83035=>"000011111",
83036=>"010001000",
83037=>"111001001",
83038=>"111111000",
83039=>"001010110",
83040=>"000000011",
83041=>"000000011",
83042=>"010000000",
83043=>"011000000",
83044=>"000111010",
83045=>"000000100",
83046=>"000000000",
83047=>"100111011",
83048=>"100001010",
83049=>"000001111",
83050=>"111000111",
83051=>"000101111",
83052=>"010010010",
83053=>"111101101",
83054=>"000000000",
83055=>"110101001",
83056=>"011011111",
83057=>"111001111",
83058=>"110001000",
83059=>"000001011",
83060=>"011111000",
83061=>"000100001",
83062=>"000111010",
83063=>"000000011",
83064=>"010000000",
83065=>"110101110",
83066=>"111001100",
83067=>"000100011",
83068=>"011100100",
83069=>"000110000",
83070=>"111000000",
83071=>"000000111",
83072=>"010010011",
83073=>"100110101",
83074=>"000000011",
83075=>"000111111",
83076=>"101100000",
83077=>"000111111",
83078=>"100110011",
83079=>"110000011",
83080=>"011111111",
83081=>"111111001",
83082=>"100111000",
83083=>"000010110",
83084=>"111000100",
83085=>"000101101",
83086=>"110111100",
83087=>"001101100",
83088=>"000111111",
83089=>"111100101",
83090=>"110100101",
83091=>"010010111",
83092=>"100000111",
83093=>"111000000",
83094=>"111000101",
83095=>"100101110",
83096=>"000000001",
83097=>"010110111",
83098=>"111000100",
83099=>"000100110",
83100=>"011011110",
83101=>"000000011",
83102=>"011111001",
83103=>"000111111",
83104=>"111011000",
83105=>"111000000",
83106=>"000111111",
83107=>"111010000",
83108=>"100111111",
83109=>"000110110",
83110=>"000110110",
83111=>"011111100",
83112=>"100000000",
83113=>"000000001",
83114=>"111000000",
83115=>"111000000",
83116=>"100101111",
83117=>"011000111",
83118=>"111101001",
83119=>"111001000",
83120=>"100101101",
83121=>"011100111",
83122=>"000000000",
83123=>"011001100",
83124=>"111111111",
83125=>"100000010",
83126=>"000100101",
83127=>"010010011",
83128=>"000100011",
83129=>"010000111",
83130=>"000010010",
83131=>"011111101",
83132=>"000011111",
83133=>"111111111",
83134=>"000011110",
83135=>"001000100",
83136=>"111001000",
83137=>"001011011",
83138=>"111111000",
83139=>"011111110",
83140=>"000111110",
83141=>"000100100",
83142=>"000011111",
83143=>"111101100",
83144=>"001000101",
83145=>"101000000",
83146=>"000001000",
83147=>"000010111",
83148=>"011010000",
83149=>"111111000",
83150=>"011101011",
83151=>"111000000",
83152=>"110111111",
83153=>"000111010",
83154=>"111101110",
83155=>"101111100",
83156=>"000000010",
83157=>"101001010",
83158=>"010000000",
83159=>"111001101",
83160=>"000011011",
83161=>"100000111",
83162=>"111111000",
83163=>"000000000",
83164=>"111111000",
83165=>"111000110",
83166=>"101111111",
83167=>"010001000",
83168=>"111000000",
83169=>"111101100",
83170=>"100000110",
83171=>"100110100",
83172=>"001000100",
83173=>"000111111",
83174=>"000111111",
83175=>"111111001",
83176=>"000111111",
83177=>"011110110",
83178=>"110110111",
83179=>"001000000",
83180=>"100000111",
83181=>"000001000",
83182=>"000001011",
83183=>"010010111",
83184=>"000011111",
83185=>"010001011",
83186=>"000000010",
83187=>"000010110",
83188=>"010110000",
83189=>"100100000",
83190=>"000000010",
83191=>"000000111",
83192=>"111010000",
83193=>"001010000",
83194=>"011111000",
83195=>"000101101",
83196=>"111111000",
83197=>"000011111",
83198=>"000111001",
83199=>"001111000",
83200=>"010101111",
83201=>"000010010",
83202=>"111110000",
83203=>"000011011",
83204=>"010000111",
83205=>"001111111",
83206=>"100000101",
83207=>"100000000",
83208=>"000011111",
83209=>"110000000",
83210=>"111100010",
83211=>"000100100",
83212=>"000000111",
83213=>"000111111",
83214=>"000100011",
83215=>"111100100",
83216=>"111000000",
83217=>"010000000",
83218=>"111010011",
83219=>"000000000",
83220=>"101111001",
83221=>"110000010",
83222=>"101111111",
83223=>"111111010",
83224=>"000000000",
83225=>"111001001",
83226=>"000000000",
83227=>"000000111",
83228=>"011000000",
83229=>"101111110",
83230=>"010000101",
83231=>"101001111",
83232=>"111111001",
83233=>"101111111",
83234=>"101101110",
83235=>"110111111",
83236=>"110111101",
83237=>"111001011",
83238=>"000000000",
83239=>"011001000",
83240=>"111000000",
83241=>"110110000",
83242=>"000110111",
83243=>"001000110",
83244=>"000111111",
83245=>"000010000",
83246=>"101111111",
83247=>"010001100",
83248=>"000000000",
83249=>"001110100",
83250=>"111000111",
83251=>"000100001",
83252=>"011000111",
83253=>"000001110",
83254=>"110110111",
83255=>"011111111",
83256=>"000000110",
83257=>"110110101",
83258=>"111010101",
83259=>"111000111",
83260=>"000100111",
83261=>"111001001",
83262=>"000000100",
83263=>"001000001",
83264=>"001000000",
83265=>"101111011",
83266=>"001110111",
83267=>"100110110",
83268=>"111110100",
83269=>"001001100",
83270=>"100100100",
83271=>"000010110",
83272=>"111111111",
83273=>"111000000",
83274=>"111111001",
83275=>"000000000",
83276=>"111000000",
83277=>"010000111",
83278=>"001001000",
83279=>"000000110",
83280=>"101101100",
83281=>"111000000",
83282=>"000000011",
83283=>"110000001",
83284=>"000000111",
83285=>"111010100",
83286=>"111100101",
83287=>"111000000",
83288=>"000001000",
83289=>"000000011",
83290=>"000000010",
83291=>"111000000",
83292=>"101010000",
83293=>"110110001",
83294=>"111000000",
83295=>"011011011",
83296=>"000000111",
83297=>"000101111",
83298=>"000000001",
83299=>"001000100",
83300=>"000000100",
83301=>"111011111",
83302=>"111110000",
83303=>"110110010",
83304=>"000000000",
83305=>"111000101",
83306=>"000000111",
83307=>"111101110",
83308=>"000011111",
83309=>"111000010",
83310=>"000000010",
83311=>"000000001",
83312=>"100011011",
83313=>"011110111",
83314=>"011011100",
83315=>"001101110",
83316=>"110000000",
83317=>"100000000",
83318=>"000000000",
83319=>"000010111",
83320=>"001110111",
83321=>"111101011",
83322=>"000000000",
83323=>"011111011",
83324=>"011011101",
83325=>"100000100",
83326=>"101010001",
83327=>"111111000",
83328=>"101000001",
83329=>"111000111",
83330=>"111010010",
83331=>"000000110",
83332=>"000000000",
83333=>"001111110",
83334=>"111101111",
83335=>"111111110",
83336=>"101100100",
83337=>"001101000",
83338=>"000100010",
83339=>"111111001",
83340=>"000000000",
83341=>"111110001",
83342=>"000000111",
83343=>"000001001",
83344=>"000000011",
83345=>"000000111",
83346=>"111000000",
83347=>"000111101",
83348=>"000110100",
83349=>"000010111",
83350=>"111111111",
83351=>"000000011",
83352=>"101100111",
83353=>"111001110",
83354=>"111011000",
83355=>"100110000",
83356=>"000001101",
83357=>"111011000",
83358=>"000000111",
83359=>"000000111",
83360=>"111010011",
83361=>"011111010",
83362=>"111111011",
83363=>"111100111",
83364=>"011010111",
83365=>"100110110",
83366=>"001001000",
83367=>"000010110",
83368=>"111010000",
83369=>"000000111",
83370=>"010111111",
83371=>"100000101",
83372=>"000001000",
83373=>"000000111",
83374=>"111110110",
83375=>"000100111",
83376=>"000000111",
83377=>"110111111",
83378=>"111000100",
83379=>"010001110",
83380=>"000011011",
83381=>"001011010",
83382=>"001000100",
83383=>"000000111",
83384=>"000010011",
83385=>"001111111",
83386=>"000000110",
83387=>"111111000",
83388=>"000100010",
83389=>"110000101",
83390=>"000000100",
83391=>"000010101",
83392=>"111111010",
83393=>"111111000",
83394=>"111001010",
83395=>"101100111",
83396=>"000000000",
83397=>"111111011",
83398=>"000001111",
83399=>"111111110",
83400=>"001010110",
83401=>"000111100",
83402=>"111111110",
83403=>"111000101",
83404=>"111000000",
83405=>"000100110",
83406=>"111111000",
83407=>"110111001",
83408=>"000000111",
83409=>"011110111",
83410=>"110110100",
83411=>"000000111",
83412=>"000000111",
83413=>"111110100",
83414=>"111111111",
83415=>"101001100",
83416=>"000000000",
83417=>"010001000",
83418=>"001100110",
83419=>"110101000",
83420=>"111101100",
83421=>"000001111",
83422=>"000001111",
83423=>"000000011",
83424=>"111000000",
83425=>"000000110",
83426=>"001000010",
83427=>"010011001",
83428=>"010000000",
83429=>"000000000",
83430=>"000111111",
83431=>"111001111",
83432=>"000110111",
83433=>"101101111",
83434=>"111011110",
83435=>"000010000",
83436=>"101000000",
83437=>"100001111",
83438=>"111000000",
83439=>"000000110",
83440=>"010000001",
83441=>"111111111",
83442=>"000111110",
83443=>"010011100",
83444=>"100100101",
83445=>"000001000",
83446=>"101000000",
83447=>"000001010",
83448=>"111110000",
83449=>"001000010",
83450=>"110101111",
83451=>"000011011",
83452=>"011000010",
83453=>"000110111",
83454=>"001001111",
83455=>"100101000",
83456=>"011001000",
83457=>"000000101",
83458=>"000000000",
83459=>"111101111",
83460=>"100000000",
83461=>"001100100",
83462=>"111111000",
83463=>"111111111",
83464=>"111001000",
83465=>"110111011",
83466=>"100100110",
83467=>"001101111",
83468=>"000000001",
83469=>"111001000",
83470=>"101011011",
83471=>"101111101",
83472=>"011101011",
83473=>"000111000",
83474=>"000010010",
83475=>"101111111",
83476=>"111010000",
83477=>"000000111",
83478=>"011001111",
83479=>"010111111",
83480=>"101000000",
83481=>"011000111",
83482=>"111101111",
83483=>"111011110",
83484=>"110010111",
83485=>"000100000",
83486=>"111000010",
83487=>"000111011",
83488=>"101000100",
83489=>"101001001",
83490=>"101000010",
83491=>"111111011",
83492=>"111110100",
83493=>"010111000",
83494=>"101000111",
83495=>"000110111",
83496=>"101001111",
83497=>"111111111",
83498=>"000000111",
83499=>"111000010",
83500=>"111111010",
83501=>"011000111",
83502=>"011000000",
83503=>"111111000",
83504=>"111000101",
83505=>"111101100",
83506=>"111101010",
83507=>"111000001",
83508=>"101111100",
83509=>"011101100",
83510=>"110111111",
83511=>"110000111",
83512=>"000000001",
83513=>"111010110",
83514=>"000000111",
83515=>"111000110",
83516=>"111110011",
83517=>"010111010",
83518=>"000000000",
83519=>"011001001",
83520=>"001000000",
83521=>"111111000",
83522=>"000001111",
83523=>"100110100",
83524=>"100000000",
83525=>"010000001",
83526=>"010010000",
83527=>"110100000",
83528=>"000010000",
83529=>"111111000",
83530=>"000000111",
83531=>"010110000",
83532=>"000000000",
83533=>"111101000",
83534=>"101101000",
83535=>"111100111",
83536=>"111101101",
83537=>"010111000",
83538=>"111010000",
83539=>"011011000",
83540=>"000000010",
83541=>"001100110",
83542=>"111111110",
83543=>"010110000",
83544=>"001000100",
83545=>"101001001",
83546=>"111110100",
83547=>"000001000",
83548=>"010111111",
83549=>"001000001",
83550=>"101000011",
83551=>"101111000",
83552=>"101001111",
83553=>"000010111",
83554=>"000111000",
83555=>"010001001",
83556=>"111001000",
83557=>"111011010",
83558=>"001000010",
83559=>"010111001",
83560=>"000100101",
83561=>"000000000",
83562=>"101001000",
83563=>"000010111",
83564=>"000000110",
83565=>"110000000",
83566=>"000000111",
83567=>"000000111",
83568=>"001001100",
83569=>"111000011",
83570=>"011011110",
83571=>"001000100",
83572=>"101110000",
83573=>"000000110",
83574=>"000111111",
83575=>"000000001",
83576=>"010000011",
83577=>"110010111",
83578=>"101000000",
83579=>"001000000",
83580=>"110110110",
83581=>"100100010",
83582=>"010001101",
83583=>"010110100",
83584=>"000000101",
83585=>"010000110",
83586=>"111010000",
83587=>"111111111",
83588=>"111101111",
83589=>"010110111",
83590=>"011110000",
83591=>"011010000",
83592=>"000100000",
83593=>"011111111",
83594=>"111111111",
83595=>"000000010",
83596=>"000000001",
83597=>"000000100",
83598=>"001000000",
83599=>"000001101",
83600=>"100100100",
83601=>"000111000",
83602=>"000111111",
83603=>"011000000",
83604=>"000000111",
83605=>"111111001",
83606=>"101001010",
83607=>"110100100",
83608=>"010101000",
83609=>"100010111",
83610=>"001000111",
83611=>"000000010",
83612=>"001011111",
83613=>"000000000",
83614=>"111001000",
83615=>"011111010",
83616=>"000001000",
83617=>"101010011",
83618=>"000000001",
83619=>"111110111",
83620=>"000111111",
83621=>"000100110",
83622=>"001101001",
83623=>"001001000",
83624=>"111111011",
83625=>"000000000",
83626=>"100000000",
83627=>"000111011",
83628=>"011001000",
83629=>"000000110",
83630=>"110110010",
83631=>"111001010",
83632=>"000000111",
83633=>"111000011",
83634=>"000000000",
83635=>"000100110",
83636=>"111110111",
83637=>"101110111",
83638=>"111100011",
83639=>"111111111",
83640=>"111011011",
83641=>"010011111",
83642=>"000000010",
83643=>"111010000",
83644=>"000000101",
83645=>"000000000",
83646=>"100111001",
83647=>"000000101",
83648=>"011010010",
83649=>"111110111",
83650=>"000110111",
83651=>"010101001",
83652=>"000000101",
83653=>"001101000",
83654=>"000000111",
83655=>"110111000",
83656=>"101110111",
83657=>"111000000",
83658=>"100000000",
83659=>"111111000",
83660=>"000000001",
83661=>"110111011",
83662=>"010010000",
83663=>"110111101",
83664=>"011000000",
83665=>"011011000",
83666=>"111110011",
83667=>"110101111",
83668=>"110000000",
83669=>"100000000",
83670=>"111111111",
83671=>"111111001",
83672=>"010110101",
83673=>"000000111",
83674=>"001110000",
83675=>"001001000",
83676=>"100000111",
83677=>"000000100",
83678=>"011100111",
83679=>"111001011",
83680=>"010000000",
83681=>"101000000",
83682=>"110111000",
83683=>"101101110",
83684=>"000110000",
83685=>"110101101",
83686=>"000000000",
83687=>"011111101",
83688=>"000000001",
83689=>"111010000",
83690=>"001001011",
83691=>"111101110",
83692=>"000000011",
83693=>"101101001",
83694=>"000000000",
83695=>"000100001",
83696=>"111111101",
83697=>"010111010",
83698=>"101101111",
83699=>"111101111",
83700=>"111001011",
83701=>"111111101",
83702=>"000000000",
83703=>"101000111",
83704=>"111010010",
83705=>"000000010",
83706=>"111110010",
83707=>"111111111",
83708=>"011001111",
83709=>"011010111",
83710=>"001001001",
83711=>"000010111",
83712=>"011011001",
83713=>"000101111",
83714=>"001100100",
83715=>"000000101",
83716=>"110111111",
83717=>"010010000",
83718=>"101000001",
83719=>"000000111",
83720=>"011111010",
83721=>"111111011",
83722=>"100100000",
83723=>"010010101",
83724=>"100000111",
83725=>"010011111",
83726=>"010100001",
83727=>"001000100",
83728=>"000000000",
83729=>"100100100",
83730=>"000111001",
83731=>"010000000",
83732=>"100000011",
83733=>"000010000",
83734=>"000101100",
83735=>"111010101",
83736=>"111100111",
83737=>"111111110",
83738=>"011011001",
83739=>"100111010",
83740=>"000101111",
83741=>"000100100",
83742=>"111111000",
83743=>"100000000",
83744=>"011000111",
83745=>"000011011",
83746=>"100100000",
83747=>"000010000",
83748=>"111011011",
83749=>"011111111",
83750=>"010000010",
83751=>"100101101",
83752=>"011011011",
83753=>"100111001",
83754=>"001011000",
83755=>"000111111",
83756=>"000100100",
83757=>"010100100",
83758=>"010111111",
83759=>"000110110",
83760=>"000100100",
83761=>"001111011",
83762=>"000011011",
83763=>"101101100",
83764=>"101110010",
83765=>"100000010",
83766=>"011010111",
83767=>"011011111",
83768=>"011111001",
83769=>"100100000",
83770=>"111000011",
83771=>"100010100",
83772=>"110011111",
83773=>"110111111",
83774=>"000000100",
83775=>"100111101",
83776=>"100100000",
83777=>"010100111",
83778=>"001011111",
83779=>"000001000",
83780=>"001001111",
83781=>"100101111",
83782=>"000000111",
83783=>"111011000",
83784=>"000110111",
83785=>"000000100",
83786=>"101100000",
83787=>"111001010",
83788=>"011111111",
83789=>"011111110",
83790=>"111111111",
83791=>"101100100",
83792=>"101100100",
83793=>"011111111",
83794=>"010100101",
83795=>"011101100",
83796=>"100100110",
83797=>"101001011",
83798=>"001001001",
83799=>"000000000",
83800=>"111110101",
83801=>"001100110",
83802=>"101111011",
83803=>"110110110",
83804=>"000000000",
83805=>"000000001",
83806=>"001011011",
83807=>"010000000",
83808=>"000010000",
83809=>"000000000",
83810=>"001000000",
83811=>"111111001",
83812=>"110010110",
83813=>"000100100",
83814=>"000000000",
83815=>"011011011",
83816=>"111011111",
83817=>"011011000",
83818=>"000011001",
83819=>"010010000",
83820=>"010110111",
83821=>"100000000",
83822=>"111110111",
83823=>"101100111",
83824=>"111111011",
83825=>"000000000",
83826=>"110010001",
83827=>"100100000",
83828=>"111011010",
83829=>"100000000",
83830=>"111111011",
83831=>"000100011",
83832=>"111100101",
83833=>"100000000",
83834=>"101000010",
83835=>"101111101",
83836=>"110110111",
83837=>"010010100",
83838=>"100101101",
83839=>"010010010",
83840=>"000000000",
83841=>"111100000",
83842=>"011011010",
83843=>"000000111",
83844=>"011101000",
83845=>"000000001",
83846=>"010111111",
83847=>"000100110",
83848=>"100000001",
83849=>"000000110",
83850=>"111100100",
83851=>"111010000",
83852=>"111111011",
83853=>"111001101",
83854=>"100011111",
83855=>"101000000",
83856=>"111011011",
83857=>"010111111",
83858=>"000000000",
83859=>"111101100",
83860=>"101111011",
83861=>"011011000",
83862=>"111011010",
83863=>"001001111",
83864=>"111011111",
83865=>"101101011",
83866=>"010010000",
83867=>"000010000",
83868=>"011011011",
83869=>"000011010",
83870=>"011001010",
83871=>"100100100",
83872=>"101111111",
83873=>"100100001",
83874=>"000000000",
83875=>"101000001",
83876=>"111111111",
83877=>"001011001",
83878=>"111111000",
83879=>"010111111",
83880=>"100111111",
83881=>"000111101",
83882=>"010010010",
83883=>"000100000",
83884=>"111111111",
83885=>"111000100",
83886=>"110010001",
83887=>"000000011",
83888=>"001111110",
83889=>"001001011",
83890=>"111000011",
83891=>"000100010",
83892=>"100100000",
83893=>"000000110",
83894=>"110100100",
83895=>"010000010",
83896=>"011111111",
83897=>"101011011",
83898=>"011000111",
83899=>"011000000",
83900=>"111110111",
83901=>"111111011",
83902=>"111011001",
83903=>"011011110",
83904=>"100000100",
83905=>"000000000",
83906=>"111000010",
83907=>"100111110",
83908=>"101000000",
83909=>"111011110",
83910=>"101111111",
83911=>"010111011",
83912=>"010010000",
83913=>"100101000",
83914=>"000000101",
83915=>"011110111",
83916=>"011011011",
83917=>"001011111",
83918=>"010000010",
83919=>"111111011",
83920=>"010000000",
83921=>"110110110",
83922=>"000110111",
83923=>"100100000",
83924=>"000000111",
83925=>"000010111",
83926=>"000000000",
83927=>"000000001",
83928=>"100000100",
83929=>"010000000",
83930=>"101101101",
83931=>"101100100",
83932=>"100110110",
83933=>"111111111",
83934=>"100101101",
83935=>"010000000",
83936=>"111100110",
83937=>"101000100",
83938=>"101001111",
83939=>"000000101",
83940=>"000000000",
83941=>"011111111",
83942=>"010011010",
83943=>"000100110",
83944=>"011111011",
83945=>"010000111",
83946=>"100000000",
83947=>"000000000",
83948=>"000000000",
83949=>"000000011",
83950=>"111111000",
83951=>"000111111",
83952=>"010011000",
83953=>"111011000",
83954=>"010000100",
83955=>"001000001",
83956=>"110000110",
83957=>"000100000",
83958=>"000000100",
83959=>"010111111",
83960=>"000000010",
83961=>"100101000",
83962=>"100100100",
83963=>"111110101",
83964=>"010011010",
83965=>"111011111",
83966=>"110111010",
83967=>"000100100",
83968=>"011011110",
83969=>"110111110",
83970=>"000000010",
83971=>"000110110",
83972=>"000000100",
83973=>"000111111",
83974=>"111001101",
83975=>"000000111",
83976=>"000000000",
83977=>"000000000",
83978=>"111111011",
83979=>"111111111",
83980=>"000110100",
83981=>"101000101",
83982=>"101011001",
83983=>"111010001",
83984=>"110000000",
83985=>"111110111",
83986=>"111010000",
83987=>"110111111",
83988=>"111011010",
83989=>"111110110",
83990=>"110110110",
83991=>"111000000",
83992=>"000000000",
83993=>"111101111",
83994=>"111111111",
83995=>"111110110",
83996=>"111111111",
83997=>"101100111",
83998=>"010000001",
83999=>"000000001",
84000=>"111110111",
84001=>"111111111",
84002=>"001000000",
84003=>"000101000",
84004=>"110111011",
84005=>"111110101",
84006=>"010000010",
84007=>"000011000",
84008=>"010010110",
84009=>"000110110",
84010=>"111111100",
84011=>"111111010",
84012=>"111011111",
84013=>"000110110",
84014=>"111111111",
84015=>"000001000",
84016=>"000000000",
84017=>"110110110",
84018=>"011100000",
84019=>"111111001",
84020=>"111001101",
84021=>"111111101",
84022=>"111111110",
84023=>"000000000",
84024=>"110111110",
84025=>"110111010",
84026=>"000000000",
84027=>"010011111",
84028=>"101010010",
84029=>"111011011",
84030=>"000101101",
84031=>"000000000",
84032=>"010110110",
84033=>"111110110",
84034=>"010000000",
84035=>"000010110",
84036=>"100000001",
84037=>"001001000",
84038=>"111001111",
84039=>"011001111",
84040=>"111111010",
84041=>"111110101",
84042=>"000110010",
84043=>"001000000",
84044=>"000111101",
84045=>"111011100",
84046=>"000111100",
84047=>"000111110",
84048=>"111110111",
84049=>"000010010",
84050=>"000000000",
84051=>"001000100",
84052=>"010000010",
84053=>"110010110",
84054=>"111000000",
84055=>"101111111",
84056=>"100110110",
84057=>"110100001",
84058=>"111111111",
84059=>"111000011",
84060=>"000000000",
84061=>"001001001",
84062=>"010010000",
84063=>"110110111",
84064=>"000000101",
84065=>"101111111",
84066=>"000110110",
84067=>"110000000",
84068=>"101111101",
84069=>"000000000",
84070=>"111111101",
84071=>"000000000",
84072=>"000000000",
84073=>"111100100",
84074=>"010011101",
84075=>"111110110",
84076=>"000000000",
84077=>"111111010",
84078=>"100000000",
84079=>"111111101",
84080=>"101101101",
84081=>"111110100",
84082=>"110111111",
84083=>"001101000",
84084=>"100000011",
84085=>"110000001",
84086=>"111111111",
84087=>"000000110",
84088=>"000111011",
84089=>"111111101",
84090=>"000000011",
84091=>"000000011",
84092=>"100110100",
84093=>"000000001",
84094=>"000000001",
84095=>"101000111",
84096=>"111111000",
84097=>"111111000",
84098=>"000000000",
84099=>"010111111",
84100=>"000000000",
84101=>"010001111",
84102=>"110011011",
84103=>"101110110",
84104=>"011001111",
84105=>"111100001",
84106=>"000000000",
84107=>"001000000",
84108=>"000000100",
84109=>"011101101",
84110=>"000000011",
84111=>"001001000",
84112=>"011011001",
84113=>"110110101",
84114=>"111011111",
84115=>"111101000",
84116=>"111101101",
84117=>"111111111",
84118=>"110110000",
84119=>"000001111",
84120=>"011111101",
84121=>"010101111",
84122=>"111011111",
84123=>"000000010",
84124=>"101001001",
84125=>"000000001",
84126=>"100110111",
84127=>"111110110",
84128=>"011110000",
84129=>"110111111",
84130=>"110100010",
84131=>"110111011",
84132=>"111000001",
84133=>"110011110",
84134=>"011010000",
84135=>"111111111",
84136=>"111111110",
84137=>"000000010",
84138=>"000000110",
84139=>"111111000",
84140=>"000101011",
84141=>"111011111",
84142=>"111111111",
84143=>"000111111",
84144=>"000000100",
84145=>"111111110",
84146=>"000101001",
84147=>"001001000",
84148=>"111100001",
84149=>"000000000",
84150=>"110000111",
84151=>"111111111",
84152=>"011000111",
84153=>"100100111",
84154=>"010010111",
84155=>"100110111",
84156=>"101101010",
84157=>"111001001",
84158=>"000000000",
84159=>"110000111",
84160=>"100010000",
84161=>"011000001",
84162=>"111111110",
84163=>"000010110",
84164=>"000000000",
84165=>"110100010",
84166=>"100000000",
84167=>"011111101",
84168=>"010011011",
84169=>"110110010",
84170=>"001111111",
84171=>"000010110",
84172=>"110110111",
84173=>"001011001",
84174=>"110110100",
84175=>"000000000",
84176=>"111111111",
84177=>"110001001",
84178=>"101111100",
84179=>"111010000",
84180=>"000000000",
84181=>"110110000",
84182=>"011110101",
84183=>"010000000",
84184=>"000000000",
84185=>"111101001",
84186=>"111011111",
84187=>"101011000",
84188=>"110110011",
84189=>"000001001",
84190=>"110100100",
84191=>"011000000",
84192=>"000000000",
84193=>"000010010",
84194=>"000000000",
84195=>"110111000",
84196=>"000000000",
84197=>"000110111",
84198=>"000000101",
84199=>"101111110",
84200=>"000101111",
84201=>"000000000",
84202=>"111101111",
84203=>"001111101",
84204=>"000100000",
84205=>"000000000",
84206=>"001110000",
84207=>"001001111",
84208=>"111000110",
84209=>"111110001",
84210=>"010000000",
84211=>"011111100",
84212=>"100100111",
84213=>"101111000",
84214=>"000000000",
84215=>"001000001",
84216=>"111110000",
84217=>"000001000",
84218=>"111111110",
84219=>"001011111",
84220=>"010110000",
84221=>"100100111",
84222=>"110110111",
84223=>"110111010",
84224=>"111100010",
84225=>"101000000",
84226=>"000000111",
84227=>"111111000",
84228=>"001011000",
84229=>"001000001",
84230=>"000111100",
84231=>"111111111",
84232=>"111101000",
84233=>"110110111",
84234=>"000000101",
84235=>"111110100",
84236=>"010110000",
84237=>"001101000",
84238=>"011000000",
84239=>"111001101",
84240=>"111001111",
84241=>"010000000",
84242=>"001110101",
84243=>"111111000",
84244=>"010111101",
84245=>"111000000",
84246=>"111011001",
84247=>"001010000",
84248=>"101111000",
84249=>"110111000",
84250=>"111011000",
84251=>"000010000",
84252=>"111001000",
84253=>"110110110",
84254=>"000110111",
84255=>"010000000",
84256=>"111001011",
84257=>"010000001",
84258=>"001000000",
84259=>"111101000",
84260=>"101000000",
84261=>"111011000",
84262=>"111110000",
84263=>"111101001",
84264=>"000000101",
84265=>"111111001",
84266=>"011011000",
84267=>"001000101",
84268=>"111000000",
84269=>"001111000",
84270=>"000000011",
84271=>"011011001",
84272=>"000110000",
84273=>"111000000",
84274=>"111111000",
84275=>"101111001",
84276=>"111000111",
84277=>"000000000",
84278=>"111010001",
84279=>"110111000",
84280=>"000000111",
84281=>"000011000",
84282=>"001111000",
84283=>"100011000",
84284=>"111011010",
84285=>"111000111",
84286=>"011000000",
84287=>"111000000",
84288=>"000101000",
84289=>"000001110",
84290=>"111111000",
84291=>"100100111",
84292=>"000000100",
84293=>"000010111",
84294=>"110111010",
84295=>"000010111",
84296=>"011111000",
84297=>"001000000",
84298=>"111001011",
84299=>"110000001",
84300=>"000110111",
84301=>"101000000",
84302=>"101000000",
84303=>"111101000",
84304=>"101000101",
84305=>"000111111",
84306=>"111011000",
84307=>"110000000",
84308=>"011110000",
84309=>"100111011",
84310=>"111000010",
84311=>"010111000",
84312=>"111110000",
84313=>"111010000",
84314=>"111001000",
84315=>"100111001",
84316=>"111101001",
84317=>"011000000",
84318=>"011101111",
84319=>"011001001",
84320=>"111000000",
84321=>"111101001",
84322=>"000111111",
84323=>"111000000",
84324=>"111000000",
84325=>"101000101",
84326=>"010011000",
84327=>"111000000",
84328=>"111111000",
84329=>"101000111",
84330=>"111111111",
84331=>"111111110",
84332=>"111101010",
84333=>"010110000",
84334=>"000101111",
84335=>"111111100",
84336=>"111000000",
84337=>"101111101",
84338=>"111010000",
84339=>"010010000",
84340=>"111101000",
84341=>"010011110",
84342=>"111111000",
84343=>"010000001",
84344=>"011111111",
84345=>"000100100",
84346=>"101101011",
84347=>"001000001",
84348=>"011011000",
84349=>"000000000",
84350=>"011000111",
84351=>"111000010",
84352=>"010011001",
84353=>"000000100",
84354=>"010001000",
84355=>"000111111",
84356=>"010111100",
84357=>"111010010",
84358=>"100100000",
84359=>"001100000",
84360=>"110000000",
84361=>"101000111",
84362=>"111011000",
84363=>"000111111",
84364=>"000000110",
84365=>"100000111",
84366=>"001111111",
84367=>"000000011",
84368=>"100000000",
84369=>"111101000",
84370=>"110111110",
84371=>"001101001",
84372=>"111101000",
84373=>"000111101",
84374=>"011010100",
84375=>"111000000",
84376=>"101111000",
84377=>"000110110",
84378=>"100111100",
84379=>"111111000",
84380=>"000111111",
84381=>"101100000",
84382=>"111110011",
84383=>"000010000",
84384=>"000111000",
84385=>"100111110",
84386=>"000000000",
84387=>"001101000",
84388=>"111111000",
84389=>"001001000",
84390=>"110001111",
84391=>"111000000",
84392=>"111111101",
84393=>"110001000",
84394=>"000001001",
84395=>"111000101",
84396=>"000111111",
84397=>"001010000",
84398=>"110001000",
84399=>"001000001",
84400=>"011000111",
84401=>"111001000",
84402=>"000110111",
84403=>"100000000",
84404=>"111000000",
84405=>"101101000",
84406=>"011011100",
84407=>"111111000",
84408=>"111111010",
84409=>"101001001",
84410=>"000101111",
84411=>"000001110",
84412=>"111110101",
84413=>"000110111",
84414=>"001000000",
84415=>"000000000",
84416=>"001101000",
84417=>"111011001",
84418=>"010010000",
84419=>"111100000",
84420=>"000000000",
84421=>"000000111",
84422=>"111111001",
84423=>"111111111",
84424=>"000111111",
84425=>"010110101",
84426=>"000001000",
84427=>"000110010",
84428=>"011010000",
84429=>"110111000",
84430=>"110000110",
84431=>"000111000",
84432=>"110111000",
84433=>"110000000",
84434=>"000111100",
84435=>"000111000",
84436=>"111010111",
84437=>"101000000",
84438=>"101111000",
84439=>"111111000",
84440=>"000000000",
84441=>"110111001",
84442=>"000000000",
84443=>"000101111",
84444=>"101111100",
84445=>"011111011",
84446=>"101110110",
84447=>"110111111",
84448=>"000001000",
84449=>"000000111",
84450=>"100000000",
84451=>"111001000",
84452=>"111000000",
84453=>"110100000",
84454=>"111111000",
84455=>"011010000",
84456=>"111111000",
84457=>"111111000",
84458=>"010000000",
84459=>"001000011",
84460=>"110000000",
84461=>"111111110",
84462=>"000000111",
84463=>"001011000",
84464=>"000000000",
84465=>"000000011",
84466=>"111111010",
84467=>"111000000",
84468=>"111001001",
84469=>"101000111",
84470=>"111111111",
84471=>"010000100",
84472=>"000111101",
84473=>"010001000",
84474=>"000111111",
84475=>"110000000",
84476=>"101000100",
84477=>"111000000",
84478=>"011001001",
84479=>"110110000",
84480=>"101101100",
84481=>"011011000",
84482=>"100000111",
84483=>"101000000",
84484=>"111000000",
84485=>"111111010",
84486=>"111110111",
84487=>"011010000",
84488=>"000011000",
84489=>"000000110",
84490=>"001000001",
84491=>"011111000",
84492=>"001101011",
84493=>"000000000",
84494=>"111101000",
84495=>"001000010",
84496=>"111000000",
84497=>"000011011",
84498=>"100101111",
84499=>"010000000",
84500=>"100111111",
84501=>"000000000",
84502=>"111010100",
84503=>"010111010",
84504=>"000100111",
84505=>"110101011",
84506=>"100100000",
84507=>"101100111",
84508=>"000000000",
84509=>"101110100",
84510=>"111100000",
84511=>"010111000",
84512=>"111000000",
84513=>"000000001",
84514=>"101111111",
84515=>"110111111",
84516=>"010110000",
84517=>"111110000",
84518=>"010000000",
84519=>"000110110",
84520=>"100101111",
84521=>"010010000",
84522=>"101101000",
84523=>"000000111",
84524=>"010011001",
84525=>"100101111",
84526=>"010010110",
84527=>"001111110",
84528=>"111010000",
84529=>"011001000",
84530=>"000010111",
84531=>"000100111",
84532=>"101100111",
84533=>"111111111",
84534=>"011001001",
84535=>"100000000",
84536=>"000000111",
84537=>"000100011",
84538=>"100111010",
84539=>"000011010",
84540=>"111011001",
84541=>"111000111",
84542=>"000000101",
84543=>"001001000",
84544=>"000111111",
84545=>"111010100",
84546=>"111010111",
84547=>"101001100",
84548=>"000010110",
84549=>"000000100",
84550=>"101111111",
84551=>"000010111",
84552=>"101111111",
84553=>"000101111",
84554=>"101011111",
84555=>"000000000",
84556=>"110000000",
84557=>"000001110",
84558=>"010110100",
84559=>"101000000",
84560=>"011001100",
84561=>"000111011",
84562=>"110010010",
84563=>"001100000",
84564=>"000010001",
84565=>"111110010",
84566=>"111001000",
84567=>"111010111",
84568=>"101111010",
84569=>"000011001",
84570=>"001011000",
84571=>"011110000",
84572=>"000000010",
84573=>"001111000",
84574=>"111000111",
84575=>"100100001",
84576=>"111010000",
84577=>"111110000",
84578=>"000000111",
84579=>"100100001",
84580=>"100001101",
84581=>"100011011",
84582=>"111001000",
84583=>"101101100",
84584=>"101000000",
84585=>"101110111",
84586=>"101101111",
84587=>"010010000",
84588=>"011000000",
84589=>"000111011",
84590=>"111000000",
84591=>"100111111",
84592=>"001001000",
84593=>"000010010",
84594=>"010110100",
84595=>"011010000",
84596=>"000101101",
84597=>"000111110",
84598=>"010000001",
84599=>"011000100",
84600=>"000000101",
84601=>"101000011",
84602=>"101101111",
84603=>"000111010",
84604=>"111100100",
84605=>"110100000",
84606=>"000000111",
84607=>"010000001",
84608=>"001101000",
84609=>"010010001",
84610=>"010001000",
84611=>"000011110",
84612=>"111111110",
84613=>"111111111",
84614=>"010111000",
84615=>"110000001",
84616=>"110100000",
84617=>"111111000",
84618=>"111000000",
84619=>"011110110",
84620=>"111100101",
84621=>"101001101",
84622=>"111111100",
84623=>"010100111",
84624=>"010000110",
84625=>"100000111",
84626=>"000000000",
84627=>"101000000",
84628=>"111011011",
84629=>"101000111",
84630=>"111111111",
84631=>"011101000",
84632=>"101100000",
84633=>"000010000",
84634=>"000011010",
84635=>"101000111",
84636=>"000011000",
84637=>"101100000",
84638=>"010000000",
84639=>"110100111",
84640=>"100111011",
84641=>"110010010",
84642=>"011000000",
84643=>"111111111",
84644=>"101111111",
84645=>"000101000",
84646=>"110011000",
84647=>"101101000",
84648=>"000000011",
84649=>"111010000",
84650=>"101101011",
84651=>"111000001",
84652=>"001101111",
84653=>"000000111",
84654=>"011111001",
84655=>"000010001",
84656=>"001000111",
84657=>"001011100",
84658=>"010001000",
84659=>"111100100",
84660=>"010111000",
84661=>"111111000",
84662=>"000111111",
84663=>"000100000",
84664=>"111110100",
84665=>"000011110",
84666=>"010010000",
84667=>"110010100",
84668=>"111110110",
84669=>"100000000",
84670=>"010110000",
84671=>"000110111",
84672=>"000000111",
84673=>"100000000",
84674=>"101111000",
84675=>"110101100",
84676=>"000111010",
84677=>"100100111",
84678=>"001000000",
84679=>"111111010",
84680=>"000100101",
84681=>"000000000",
84682=>"000111101",
84683=>"000100111",
84684=>"011000100",
84685=>"011000001",
84686=>"000000000",
84687=>"000000111",
84688=>"110010000",
84689=>"110110000",
84690=>"000000101",
84691=>"110000100",
84692=>"111001111",
84693=>"110000000",
84694=>"111001111",
84695=>"001001001",
84696=>"000000000",
84697=>"000010110",
84698=>"100110111",
84699=>"001101111",
84700=>"001000001",
84701=>"010011000",
84702=>"011110101",
84703=>"100001111",
84704=>"000000000",
84705=>"111001111",
84706=>"000010100",
84707=>"111011000",
84708=>"111000111",
84709=>"000000101",
84710=>"011111000",
84711=>"101111000",
84712=>"101001000",
84713=>"001000101",
84714=>"100000100",
84715=>"010000101",
84716=>"010000010",
84717=>"010000011",
84718=>"000000000",
84719=>"001000000",
84720=>"111101000",
84721=>"000001111",
84722=>"010011000",
84723=>"001100000",
84724=>"100010000",
84725=>"100000101",
84726=>"000000001",
84727=>"001100000",
84728=>"101011010",
84729=>"101111000",
84730=>"011111110",
84731=>"111100101",
84732=>"001111000",
84733=>"111100101",
84734=>"001000000",
84735=>"001100101",
84736=>"010000000",
84737=>"100000110",
84738=>"010100001",
84739=>"100000011",
84740=>"000111111",
84741=>"000100100",
84742=>"100110101",
84743=>"000010110",
84744=>"100001000",
84745=>"010110100",
84746=>"111111011",
84747=>"110100100",
84748=>"110100000",
84749=>"010111101",
84750=>"011011111",
84751=>"011101001",
84752=>"110110110",
84753=>"010010100",
84754=>"010000000",
84755=>"000010110",
84756=>"100000100",
84757=>"110110111",
84758=>"111000001",
84759=>"000110110",
84760=>"100000000",
84761=>"110100001",
84762=>"100000110",
84763=>"110000001",
84764=>"110110110",
84765=>"011000100",
84766=>"100101000",
84767=>"011010000",
84768=>"110000100",
84769=>"001101101",
84770=>"101100100",
84771=>"111111100",
84772=>"011011010",
84773=>"100000000",
84774=>"010110100",
84775=>"001000000",
84776=>"011111110",
84777=>"010000000",
84778=>"001100100",
84779=>"010000010",
84780=>"111011111",
84781=>"100100000",
84782=>"111011001",
84783=>"000000100",
84784=>"111110000",
84785=>"000000011",
84786=>"000100000",
84787=>"101001110",
84788=>"110000001",
84789=>"110001010",
84790=>"111110010",
84791=>"111001000",
84792=>"001001001",
84793=>"100001010",
84794=>"000001001",
84795=>"111111011",
84796=>"000000000",
84797=>"111011010",
84798=>"000100000",
84799=>"111111000",
84800=>"100100001",
84801=>"000000000",
84802=>"001011110",
84803=>"000010000",
84804=>"001001001",
84805=>"000001101",
84806=>"111110010",
84807=>"111111111",
84808=>"011101001",
84809=>"110100000",
84810=>"110100100",
84811=>"010111111",
84812=>"000001001",
84813=>"101011111",
84814=>"111011000",
84815=>"110001111",
84816=>"000100000",
84817=>"011011111",
84818=>"100110111",
84819=>"011101000",
84820=>"100111010",
84821=>"000000011",
84822=>"101000001",
84823=>"110110101",
84824=>"100110111",
84825=>"011011011",
84826=>"101101001",
84827=>"111111111",
84828=>"110100000",
84829=>"001001001",
84830=>"010110110",
84831=>"010000000",
84832=>"001001100",
84833=>"100110100",
84834=>"010110111",
84835=>"001011010",
84836=>"000000001",
84837=>"011111100",
84838=>"011111000",
84839=>"011010010",
84840=>"000010101",
84841=>"101001111",
84842=>"011111110",
84843=>"011110110",
84844=>"111000011",
84845=>"111111100",
84846=>"010100100",
84847=>"001001011",
84848=>"011011111",
84849=>"010001101",
84850=>"111101001",
84851=>"111000000",
84852=>"111101110",
84853=>"000101100",
84854=>"000001100",
84855=>"001001011",
84856=>"110100100",
84857=>"010001011",
84858=>"001111110",
84859=>"110100111",
84860=>"111101101",
84861=>"000000000",
84862=>"011010110",
84863=>"000100110",
84864=>"100100101",
84865=>"001001111",
84866=>"100000000",
84867=>"001100000",
84868=>"000110100",
84869=>"111100010",
84870=>"000101111",
84871=>"111000001",
84872=>"001011011",
84873=>"000100000",
84874=>"111110010",
84875=>"111000000",
84876=>"000000110",
84877=>"000111110",
84878=>"111101000",
84879=>"110001001",
84880=>"111001011",
84881=>"000010110",
84882=>"000011010",
84883=>"001000000",
84884=>"111010110",
84885=>"010100100",
84886=>"000010011",
84887=>"000001001",
84888=>"110100110",
84889=>"011111101",
84890=>"010000010",
84891=>"011010000",
84892=>"000100111",
84893=>"000000111",
84894=>"010000010",
84895=>"001001101",
84896=>"101111001",
84897=>"000101100",
84898=>"010001001",
84899=>"011110001",
84900=>"001111111",
84901=>"010010001",
84902=>"101001001",
84903=>"111001110",
84904=>"100100111",
84905=>"100001001",
84906=>"101001001",
84907=>"000000100",
84908=>"100000001",
84909=>"100010010",
84910=>"010111111",
84911=>"111110000",
84912=>"000000100",
84913=>"011101100",
84914=>"000001001",
84915=>"001001001",
84916=>"010111111",
84917=>"101010000",
84918=>"000000101",
84919=>"011000000",
84920=>"000100111",
84921=>"010010100",
84922=>"010010100",
84923=>"110011110",
84924=>"101000000",
84925=>"001011101",
84926=>"100000101",
84927=>"010110000",
84928=>"100110101",
84929=>"000110010",
84930=>"110001011",
84931=>"011011011",
84932=>"001000001",
84933=>"000000001",
84934=>"000011011",
84935=>"010000100",
84936=>"000001001",
84937=>"001000001",
84938=>"011111011",
84939=>"110000101",
84940=>"010010011",
84941=>"001001111",
84942=>"110100000",
84943=>"110111010",
84944=>"001011011",
84945=>"101001010",
84946=>"111000000",
84947=>"011111000",
84948=>"000001001",
84949=>"100100000",
84950=>"110100001",
84951=>"000010000",
84952=>"100101000",
84953=>"111000110",
84954=>"000101011",
84955=>"110100100",
84956=>"000000011",
84957=>"001011111",
84958=>"001001111",
84959=>"101000001",
84960=>"110110100",
84961=>"111001000",
84962=>"101111100",
84963=>"110110001",
84964=>"000000000",
84965=>"000011011",
84966=>"101000111",
84967=>"110000001",
84968=>"011101011",
84969=>"110101100",
84970=>"110110000",
84971=>"001011001",
84972=>"110110000",
84973=>"101001011",
84974=>"010000000",
84975=>"100001011",
84976=>"000100110",
84977=>"111011001",
84978=>"110100101",
84979=>"010000000",
84980=>"000000011",
84981=>"001011010",
84982=>"001100000",
84983=>"011011110",
84984=>"100100101",
84985=>"100000000",
84986=>"110110110",
84987=>"001011011",
84988=>"111011011",
84989=>"011010000",
84990=>"111111110",
84991=>"011111111",
84992=>"000000000",
84993=>"000100111",
84994=>"010000000",
84995=>"000101101",
84996=>"001001001",
84997=>"000000000",
84998=>"000000000",
84999=>"000111110",
85000=>"010000101",
85001=>"001000001",
85002=>"111000000",
85003=>"111100001",
85004=>"000111000",
85005=>"000000000",
85006=>"001011000",
85007=>"010000110",
85008=>"001000000",
85009=>"111111000",
85010=>"000000000",
85011=>"101101100",
85012=>"111101000",
85013=>"101001111",
85014=>"101101001",
85015=>"110110110",
85016=>"000000001",
85017=>"111000001",
85018=>"101111111",
85019=>"110010000",
85020=>"011100001",
85021=>"010000100",
85022=>"000000000",
85023=>"111000101",
85024=>"111000111",
85025=>"000000000",
85026=>"110110001",
85027=>"111111000",
85028=>"110101001",
85029=>"000100100",
85030=>"111011000",
85031=>"000100000",
85032=>"000111111",
85033=>"111110000",
85034=>"101011111",
85035=>"000110111",
85036=>"000011111",
85037=>"111111111",
85038=>"000000000",
85039=>"001001110",
85040=>"000000011",
85041=>"101111001",
85042=>"111111111",
85043=>"111000101",
85044=>"000000000",
85045=>"001101111",
85046=>"110001000",
85047=>"110000000",
85048=>"000010101",
85049=>"111100000",
85050=>"000000111",
85051=>"111101110",
85052=>"110110100",
85053=>"000000010",
85054=>"110000000",
85055=>"001001000",
85056=>"010010001",
85057=>"110000000",
85058=>"111111110",
85059=>"000110000",
85060=>"111111111",
85061=>"110111111",
85062=>"010111001",
85063=>"110100111",
85064=>"001011111",
85065=>"111111000",
85066=>"001111011",
85067=>"000111010",
85068=>"000010000",
85069=>"101101101",
85070=>"011111100",
85071=>"111100001",
85072=>"110000000",
85073=>"011001111",
85074=>"100101000",
85075=>"000100110",
85076=>"000110000",
85077=>"110101001",
85078=>"001011100",
85079=>"101000000",
85080=>"010000111",
85081=>"001000110",
85082=>"110010011",
85083=>"011110000",
85084=>"111001000",
85085=>"001000111",
85086=>"001111011",
85087=>"000011000",
85088=>"101111010",
85089=>"000000111",
85090=>"111001000",
85091=>"100000011",
85092=>"000100000",
85093=>"111010010",
85094=>"110111000",
85095=>"111001000",
85096=>"001111110",
85097=>"111001000",
85098=>"111111111",
85099=>"111100111",
85100=>"101001000",
85101=>"010010110",
85102=>"100000000",
85103=>"111010011",
85104=>"000000000",
85105=>"010010111",
85106=>"011100000",
85107=>"111110000",
85108=>"111111010",
85109=>"000000000",
85110=>"000111111",
85111=>"001110000",
85112=>"010010111",
85113=>"100000000",
85114=>"000001000",
85115=>"000101111",
85116=>"100110110",
85117=>"100000000",
85118=>"110000000",
85119=>"000000000",
85120=>"110010000",
85121=>"000000000",
85122=>"000000111",
85123=>"101000111",
85124=>"111111011",
85125=>"100000000",
85126=>"000000101",
85127=>"001100000",
85128=>"000100010",
85129=>"000000000",
85130=>"111101001",
85131=>"111101100",
85132=>"000000101",
85133=>"111001001",
85134=>"000000010",
85135=>"010001000",
85136=>"100111011",
85137=>"111111000",
85138=>"100100110",
85139=>"000001000",
85140=>"000111001",
85141=>"000000001",
85142=>"001001001",
85143=>"000001011",
85144=>"111000000",
85145=>"000111111",
85146=>"001000111",
85147=>"111001001",
85148=>"000001000",
85149=>"000001001",
85150=>"010101111",
85151=>"000010011",
85152=>"111100101",
85153=>"111010111",
85154=>"101001000",
85155=>"111111111",
85156=>"010000000",
85157=>"011001001",
85158=>"100100101",
85159=>"001111011",
85160=>"111110111",
85161=>"000111111",
85162=>"000100100",
85163=>"000110000",
85164=>"110111111",
85165=>"111110010",
85166=>"000001100",
85167=>"111111000",
85168=>"010101010",
85169=>"111000000",
85170=>"000000100",
85171=>"110100100",
85172=>"110110111",
85173=>"111101101",
85174=>"110100100",
85175=>"101111111",
85176=>"011011001",
85177=>"000100101",
85178=>"111000100",
85179=>"000000000",
85180=>"111111111",
85181=>"111110010",
85182=>"000000000",
85183=>"111000110",
85184=>"111000101",
85185=>"111010000",
85186=>"000110110",
85187=>"000100110",
85188=>"010111111",
85189=>"011001001",
85190=>"010010111",
85191=>"110111111",
85192=>"011011000",
85193=>"000010000",
85194=>"100000000",
85195=>"111010000",
85196=>"110110000",
85197=>"001011111",
85198=>"000000000",
85199=>"000000011",
85200=>"000010110",
85201=>"000111110",
85202=>"111000000",
85203=>"010000010",
85204=>"000000000",
85205=>"100000111",
85206=>"101101001",
85207=>"000111111",
85208=>"101101111",
85209=>"011011011",
85210=>"100011001",
85211=>"000000000",
85212=>"111001100",
85213=>"000111110",
85214=>"111101000",
85215=>"010000000",
85216=>"111110000",
85217=>"001101001",
85218=>"111101111",
85219=>"000110010",
85220=>"111010000",
85221=>"000101101",
85222=>"011011001",
85223=>"010000100",
85224=>"010111111",
85225=>"111001011",
85226=>"011000000",
85227=>"100101101",
85228=>"000111010",
85229=>"010100001",
85230=>"000000000",
85231=>"111000100",
85232=>"010000010",
85233=>"110101000",
85234=>"101000101",
85235=>"000001111",
85236=>"100010001",
85237=>"101000000",
85238=>"000000000",
85239=>"101111111",
85240=>"000001111",
85241=>"000111111",
85242=>"111000100",
85243=>"111101100",
85244=>"111010000",
85245=>"010011001",
85246=>"101101100",
85247=>"000111010",
85248=>"000011011",
85249=>"000001101",
85250=>"111101000",
85251=>"000000001",
85252=>"011000111",
85253=>"101100000",
85254=>"111101000",
85255=>"000000111",
85256=>"111111000",
85257=>"111101000",
85258=>"001111111",
85259=>"001011011",
85260=>"000000010",
85261=>"010111110",
85262=>"000101111",
85263=>"000001000",
85264=>"111101010",
85265=>"111101111",
85266=>"010010100",
85267=>"000000110",
85268=>"000010001",
85269=>"000010010",
85270=>"110101101",
85271=>"000111111",
85272=>"001000000",
85273=>"000110110",
85274=>"101000000",
85275=>"000000000",
85276=>"000010111",
85277=>"000000000",
85278=>"111010000",
85279=>"000000001",
85280=>"011010001",
85281=>"000010011",
85282=>"000000010",
85283=>"000100110",
85284=>"001011110",
85285=>"001110101",
85286=>"000010010",
85287=>"011100001",
85288=>"010110111",
85289=>"000010110",
85290=>"111101001",
85291=>"000000101",
85292=>"000100111",
85293=>"000111111",
85294=>"001000111",
85295=>"000000001",
85296=>"110111001",
85297=>"000100111",
85298=>"001000001",
85299=>"001111110",
85300=>"000100111",
85301=>"111010110",
85302=>"110001111",
85303=>"001001001",
85304=>"111111001",
85305=>"000000001",
85306=>"111001110",
85307=>"000101101",
85308=>"001111111",
85309=>"111000010",
85310=>"000000001",
85311=>"000011001",
85312=>"001100000",
85313=>"000010000",
85314=>"011101001",
85315=>"111001000",
85316=>"101001000",
85317=>"000000001",
85318=>"101000001",
85319=>"000000010",
85320=>"000111111",
85321=>"000110111",
85322=>"100000000",
85323=>"010011111",
85324=>"010010000",
85325=>"000110111",
85326=>"001001111",
85327=>"001100000",
85328=>"000010110",
85329=>"011010000",
85330=>"100110111",
85331=>"000001000",
85332=>"100111010",
85333=>"101110111",
85334=>"011011011",
85335=>"111000000",
85336=>"001110111",
85337=>"000100101",
85338=>"011001000",
85339=>"010100111",
85340=>"111001101",
85341=>"000001011",
85342=>"111111110",
85343=>"111001000",
85344=>"111111000",
85345=>"111111111",
85346=>"110000000",
85347=>"011000000",
85348=>"001111110",
85349=>"111111010",
85350=>"110110010",
85351=>"111000000",
85352=>"111100000",
85353=>"000000101",
85354=>"000100111",
85355=>"100011011",
85356=>"000000111",
85357=>"011001000",
85358=>"110110100",
85359=>"000000000",
85360=>"100111111",
85361=>"000000101",
85362=>"100100101",
85363=>"111000000",
85364=>"000000100",
85365=>"010001001",
85366=>"000000111",
85367=>"111111110",
85368=>"111000000",
85369=>"001000000",
85370=>"111111101",
85371=>"011101101",
85372=>"001000111",
85373=>"000100100",
85374=>"111101000",
85375=>"111111000",
85376=>"000111011",
85377=>"000000100",
85378=>"000000001",
85379=>"000000000",
85380=>"001010000",
85381=>"000000000",
85382=>"000100111",
85383=>"000000011",
85384=>"001111111",
85385=>"000100111",
85386=>"111111000",
85387=>"000011001",
85388=>"110100000",
85389=>"011111101",
85390=>"111011001",
85391=>"111001100",
85392=>"001111111",
85393=>"011110011",
85394=>"000001000",
85395=>"111110101",
85396=>"000000000",
85397=>"111101001",
85398=>"000111111",
85399=>"000000011",
85400=>"001101111",
85401=>"111001010",
85402=>"111010111",
85403=>"111101000",
85404=>"111011111",
85405=>"010000000",
85406=>"000111110",
85407=>"000000011",
85408=>"000111111",
85409=>"111111100",
85410=>"000000001",
85411=>"111100010",
85412=>"111111111",
85413=>"001111111",
85414=>"110010110",
85415=>"000001001",
85416=>"000110011",
85417=>"000111111",
85418=>"111000000",
85419=>"110101101",
85420=>"010011111",
85421=>"110111000",
85422=>"011000100",
85423=>"111010110",
85424=>"110000000",
85425=>"101110111",
85426=>"111111000",
85427=>"100000000",
85428=>"000000011",
85429=>"101110011",
85430=>"000000111",
85431=>"000111111",
85432=>"000010111",
85433=>"000000110",
85434=>"001001011",
85435=>"111111011",
85436=>"000010110",
85437=>"111111110",
85438=>"111011000",
85439=>"000110111",
85440=>"100010110",
85441=>"000011101",
85442=>"001111111",
85443=>"000000100",
85444=>"011110111",
85445=>"001010011",
85446=>"111100101",
85447=>"111000011",
85448=>"100000111",
85449=>"101001100",
85450=>"000110111",
85451=>"110110010",
85452=>"011001101",
85453=>"000000100",
85454=>"111111110",
85455=>"111000000",
85456=>"111000000",
85457=>"000100111",
85458=>"101000110",
85459=>"000101001",
85460=>"111000111",
85461=>"000110110",
85462=>"000011111",
85463=>"101001001",
85464=>"000000110",
85465=>"011000000",
85466=>"000000100",
85467=>"111100000",
85468=>"001001101",
85469=>"111010111",
85470=>"000111111",
85471=>"101011000",
85472=>"111101000",
85473=>"111101100",
85474=>"111000000",
85475=>"100001111",
85476=>"111101000",
85477=>"101101111",
85478=>"000001111",
85479=>"100010110",
85480=>"111101001",
85481=>"111000000",
85482=>"100110111",
85483=>"111000000",
85484=>"111010000",
85485=>"000000000",
85486=>"010100000",
85487=>"001000111",
85488=>"000000000",
85489=>"000010001",
85490=>"111111111",
85491=>"001001110",
85492=>"000000110",
85493=>"111111000",
85494=>"001000010",
85495=>"111000000",
85496=>"000000111",
85497=>"000001101",
85498=>"000111111",
85499=>"001010110",
85500=>"000111111",
85501=>"101001000",
85502=>"000100111",
85503=>"111000111",
85504=>"011011000",
85505=>"111100000",
85506=>"100000000",
85507=>"000000110",
85508=>"100111110",
85509=>"111101101",
85510=>"100111111",
85511=>"000110010",
85512=>"000110110",
85513=>"000000100",
85514=>"110000101",
85515=>"010010111",
85516=>"000000101",
85517=>"011101101",
85518=>"100100010",
85519=>"001100100",
85520=>"111111000",
85521=>"000111001",
85522=>"100110000",
85523=>"010111000",
85524=>"001011011",
85525=>"101010111",
85526=>"011111111",
85527=>"010101011",
85528=>"000010000",
85529=>"000110110",
85530=>"011000100",
85531=>"000000000",
85532=>"111111111",
85533=>"000000110",
85534=>"101010010",
85535=>"000000100",
85536=>"111000011",
85537=>"111101101",
85538=>"100000000",
85539=>"111111000",
85540=>"000101001",
85541=>"110110100",
85542=>"000000001",
85543=>"000000000",
85544=>"111110110",
85545=>"000010010",
85546=>"000000111",
85547=>"011001111",
85548=>"110101001",
85549=>"001111101",
85550=>"111100100",
85551=>"011101111",
85552=>"110100000",
85553=>"000001000",
85554=>"111101101",
85555=>"000010010",
85556=>"101100000",
85557=>"000110101",
85558=>"100100000",
85559=>"000110111",
85560=>"111010010",
85561=>"000001001",
85562=>"000101111",
85563=>"000000001",
85564=>"000100100",
85565=>"111111000",
85566=>"000000000",
85567=>"100000111",
85568=>"111000111",
85569=>"101010010",
85570=>"111000000",
85571=>"001001100",
85572=>"111101010",
85573=>"000010100",
85574=>"000000101",
85575=>"111010111",
85576=>"010000100",
85577=>"101001110",
85578=>"000000111",
85579=>"000010000",
85580=>"000000010",
85581=>"011101100",
85582=>"000100000",
85583=>"111111111",
85584=>"010000000",
85585=>"110100000",
85586=>"001000110",
85587=>"011001000",
85588=>"100000000",
85589=>"001100000",
85590=>"011000000",
85591=>"011010010",
85592=>"001101001",
85593=>"001111101",
85594=>"101000111",
85595=>"000011011",
85596=>"000010010",
85597=>"000100000",
85598=>"111000010",
85599=>"100000000",
85600=>"000010010",
85601=>"110111001",
85602=>"000000000",
85603=>"000100111",
85604=>"000000101",
85605=>"000000001",
85606=>"010100000",
85607=>"000010111",
85608=>"000001111",
85609=>"101000110",
85610=>"101111111",
85611=>"110000000",
85612=>"000101110",
85613=>"000101111",
85614=>"000000111",
85615=>"110010101",
85616=>"011111100",
85617=>"001001011",
85618=>"001001001",
85619=>"000111010",
85620=>"111100000",
85621=>"111000001",
85622=>"101000001",
85623=>"011110110",
85624=>"001000011",
85625=>"000011000",
85626=>"101111000",
85627=>"101101101",
85628=>"001001101",
85629=>"100000000",
85630=>"010000011",
85631=>"100101101",
85632=>"010000010",
85633=>"111101000",
85634=>"111111010",
85635=>"000000011",
85636=>"001010111",
85637=>"000100101",
85638=>"101011000",
85639=>"000100000",
85640=>"100111101",
85641=>"001101100",
85642=>"000011111",
85643=>"000110010",
85644=>"001000100",
85645=>"010110111",
85646=>"111100000",
85647=>"000000000",
85648=>"100111101",
85649=>"111001001",
85650=>"100000101",
85651=>"111010010",
85652=>"001101000",
85653=>"111010010",
85654=>"111101111",
85655=>"100000000",
85656=>"010010111",
85657=>"001111111",
85658=>"100100000",
85659=>"100000000",
85660=>"010101111",
85661=>"111100000",
85662=>"010010100",
85663=>"000010000",
85664=>"000011001",
85665=>"111111010",
85666=>"101000100",
85667=>"101111101",
85668=>"111000000",
85669=>"010110110",
85670=>"110110000",
85671=>"110110000",
85672=>"100001000",
85673=>"000000101",
85674=>"100000000",
85675=>"110111101",
85676=>"100000000",
85677=>"001101111",
85678=>"110110100",
85679=>"000000110",
85680=>"010000010",
85681=>"000101100",
85682=>"010101101",
85683=>"001001000",
85684=>"000101111",
85685=>"110111010",
85686=>"011011011",
85687=>"000000000",
85688=>"000001001",
85689=>"000001101",
85690=>"011111101",
85691=>"111001000",
85692=>"010100010",
85693=>"101001011",
85694=>"011101001",
85695=>"000010110",
85696=>"001001000",
85697=>"000000000",
85698=>"001010000",
85699=>"000110110",
85700=>"000001101",
85701=>"111111100",
85702=>"000000011",
85703=>"111001001",
85704=>"000000111",
85705=>"000010000",
85706=>"100110110",
85707=>"000111010",
85708=>"000111101",
85709=>"100100000",
85710=>"000101000",
85711=>"010110110",
85712=>"011111110",
85713=>"100101011",
85714=>"000111111",
85715=>"000010110",
85716=>"010010000",
85717=>"000100100",
85718=>"111100000",
85719=>"111111011",
85720=>"000111111",
85721=>"010111000",
85722=>"010110110",
85723=>"000000111",
85724=>"110101000",
85725=>"000111111",
85726=>"111111101",
85727=>"111111111",
85728=>"000000010",
85729=>"111100011",
85730=>"000000101",
85731=>"001011000",
85732=>"001000000",
85733=>"000111110",
85734=>"010001111",
85735=>"011011101",
85736=>"111001000",
85737=>"111101111",
85738=>"111001001",
85739=>"111000111",
85740=>"110000000",
85741=>"010000100",
85742=>"001000000",
85743=>"100000000",
85744=>"110110010",
85745=>"111111000",
85746=>"100010010",
85747=>"100111000",
85748=>"110110011",
85749=>"000000111",
85750=>"100000111",
85751=>"101000010",
85752=>"111000000",
85753=>"000100011",
85754=>"000001001",
85755=>"111111101",
85756=>"111100000",
85757=>"000000000",
85758=>"001111001",
85759=>"001010111",
85760=>"111000000",
85761=>"110000101",
85762=>"100100100",
85763=>"000111001",
85764=>"011010110",
85765=>"000110110",
85766=>"110111111",
85767=>"100110100",
85768=>"010000010",
85769=>"100100110",
85770=>"000101001",
85771=>"011001011",
85772=>"110110000",
85773=>"011000011",
85774=>"001011001",
85775=>"110111111",
85776=>"110100110",
85777=>"110110110",
85778=>"100100110",
85779=>"110110001",
85780=>"110100111",
85781=>"111111111",
85782=>"101111110",
85783=>"110110111",
85784=>"000010010",
85785=>"111111111",
85786=>"000001111",
85787=>"110110110",
85788=>"000011110",
85789=>"001110000",
85790=>"110110100",
85791=>"001011001",
85792=>"001100101",
85793=>"101100001",
85794=>"000011011",
85795=>"111111101",
85796=>"011101111",
85797=>"000001011",
85798=>"001011011",
85799=>"110100100",
85800=>"011011101",
85801=>"001110111",
85802=>"110100100",
85803=>"001001001",
85804=>"000101111",
85805=>"110100000",
85806=>"010100100",
85807=>"000000000",
85808=>"000110110",
85809=>"001000000",
85810=>"100111101",
85811=>"010110111",
85812=>"111001100",
85813=>"000000110",
85814=>"100100100",
85815=>"110110010",
85816=>"100000111",
85817=>"000110000",
85818=>"001001111",
85819=>"011000110",
85820=>"011101111",
85821=>"011001011",
85822=>"000000100",
85823=>"000000111",
85824=>"100111111",
85825=>"000000011",
85826=>"110110010",
85827=>"110010100",
85828=>"011001001",
85829=>"000000010",
85830=>"000100110",
85831=>"000110111",
85832=>"001000011",
85833=>"011101101",
85834=>"110100110",
85835=>"111101001",
85836=>"110101111",
85837=>"001101000",
85838=>"111111111",
85839=>"001100011",
85840=>"001001001",
85841=>"001100111",
85842=>"101100111",
85843=>"100110010",
85844=>"001001001",
85845=>"110100110",
85846=>"011001100",
85847=>"110110110",
85848=>"111111111",
85849=>"000000000",
85850=>"001001001",
85851=>"111010000",
85852=>"110110110",
85853=>"001001000",
85854=>"110110110",
85855=>"000100110",
85856=>"011011011",
85857=>"110011111",
85858=>"000100110",
85859=>"011011001",
85860=>"010111110",
85861=>"111111111",
85862=>"000001001",
85863=>"001000001",
85864=>"111101111",
85865=>"000100111",
85866=>"001100110",
85867=>"011011101",
85868=>"111001101",
85869=>"001001101",
85870=>"110110010",
85871=>"100110100",
85872=>"000000000",
85873=>"110110110",
85874=>"110110000",
85875=>"001001001",
85876=>"100111111",
85877=>"000000010",
85878=>"110110110",
85879=>"000011111",
85880=>"110110100",
85881=>"110111110",
85882=>"111011011",
85883=>"011101111",
85884=>"001100110",
85885=>"000000000",
85886=>"010100000",
85887=>"111011011",
85888=>"000100110",
85889=>"110110110",
85890=>"011000111",
85891=>"001011000",
85892=>"111111001",
85893=>"000110110",
85894=>"000110001",
85895=>"001001001",
85896=>"001001101",
85897=>"001001001",
85898=>"111110111",
85899=>"110100100",
85900=>"110010001",
85901=>"110111110",
85902=>"110110110",
85903=>"010000000",
85904=>"000000000",
85905=>"111011010",
85906=>"101000000",
85907=>"011000010",
85908=>"001000000",
85909=>"110110110",
85910=>"011111101",
85911=>"000111101",
85912=>"011011011",
85913=>"100100101",
85914=>"001111111",
85915=>"100110000",
85916=>"111110110",
85917=>"111111111",
85918=>"110111111",
85919=>"001100111",
85920=>"001001101",
85921=>"110111110",
85922=>"111110011",
85923=>"100110001",
85924=>"011110110",
85925=>"010001010",
85926=>"111100000",
85927=>"010001001",
85928=>"110110110",
85929=>"111111111",
85930=>"001010010",
85931=>"110000100",
85932=>"000101000",
85933=>"001001000",
85934=>"100100010",
85935=>"011011011",
85936=>"110100100",
85937=>"001000000",
85938=>"111011000",
85939=>"000000100",
85940=>"000001000",
85941=>"010000001",
85942=>"000011001",
85943=>"001010000",
85944=>"100100100",
85945=>"011000000",
85946=>"111101111",
85947=>"110110000",
85948=>"011011001",
85949=>"111011011",
85950=>"111101001",
85951=>"000000011",
85952=>"011001001",
85953=>"111011010",
85954=>"110000111",
85955=>"111011000",
85956=>"000000011",
85957=>"000100001",
85958=>"110100110",
85959=>"110110100",
85960=>"001000000",
85961=>"101111111",
85962=>"000100001",
85963=>"000000000",
85964=>"011111001",
85965=>"000100000",
85966=>"001001001",
85967=>"000110000",
85968=>"001001111",
85969=>"001001000",
85970=>"111111011",
85971=>"001000001",
85972=>"101000110",
85973=>"001011111",
85974=>"101100110",
85975=>"110100100",
85976=>"000000000",
85977=>"110000101",
85978=>"010101001",
85979=>"001011001",
85980=>"100110100",
85981=>"001001001",
85982=>"011001010",
85983=>"110000000",
85984=>"111110100",
85985=>"000011111",
85986=>"001101011",
85987=>"001000000",
85988=>"100000000",
85989=>"100000011",
85990=>"011011011",
85991=>"110110110",
85992=>"110010111",
85993=>"110010010",
85994=>"011001000",
85995=>"110101100",
85996=>"100110010",
85997=>"001001011",
85998=>"110000010",
85999=>"110000110",
86000=>"000000000",
86001=>"111110010",
86002=>"111110110",
86003=>"110111000",
86004=>"100100110",
86005=>"001011001",
86006=>"000000000",
86007=>"000001110",
86008=>"110110110",
86009=>"100000000",
86010=>"011011111",
86011=>"110100000",
86012=>"111001000",
86013=>"000100010",
86014=>"010011101",
86015=>"011111011",
86016=>"011011001",
86017=>"000001110",
86018=>"000100000",
86019=>"001001111",
86020=>"010101100",
86021=>"110110010",
86022=>"100110111",
86023=>"110001010",
86024=>"000000001",
86025=>"110001100",
86026=>"010110010",
86027=>"100100111",
86028=>"001110111",
86029=>"000010010",
86030=>"010001011",
86031=>"101001101",
86032=>"011111001",
86033=>"100111111",
86034=>"001011110",
86035=>"000001011",
86036=>"111111000",
86037=>"100110110",
86038=>"011000001",
86039=>"110100101",
86040=>"010000001",
86041=>"100111111",
86042=>"111111010",
86043=>"110000000",
86044=>"100000100",
86045=>"000000011",
86046=>"111000000",
86047=>"001001011",
86048=>"000110010",
86049=>"000001011",
86050=>"110101001",
86051=>"110011011",
86052=>"011001011",
86053=>"001001010",
86054=>"011011001",
86055=>"000010011",
86056=>"010111111",
86057=>"100000101",
86058=>"110011000",
86059=>"111100100",
86060=>"111111111",
86061=>"100000111",
86062=>"111101000",
86063=>"011001101",
86064=>"011000010",
86065=>"001001001",
86066=>"000111110",
86067=>"111111100",
86068=>"100110111",
86069=>"001000000",
86070=>"000001011",
86071=>"111110000",
86072=>"011101110",
86073=>"000100000",
86074=>"100000001",
86075=>"110000000",
86076=>"000000011",
86077=>"010001001",
86078=>"000010001",
86079=>"111111110",
86080=>"111110111",
86081=>"001111101",
86082=>"000110011",
86083=>"000000011",
86084=>"110000000",
86085=>"000100101",
86086=>"000100001",
86087=>"001011111",
86088=>"011001001",
86089=>"011010001",
86090=>"001001001",
86091=>"101111111",
86092=>"100110100",
86093=>"111011001",
86094=>"011001001",
86095=>"000100011",
86096=>"001010010",
86097=>"111000100",
86098=>"111110001",
86099=>"011000000",
86100=>"111111101",
86101=>"011000000",
86102=>"001001001",
86103=>"110100100",
86104=>"110000110",
86105=>"000001001",
86106=>"001001001",
86107=>"101101100",
86108=>"110101110",
86109=>"100000101",
86110=>"110011110",
86111=>"000111100",
86112=>"110110110",
86113=>"000010110",
86114=>"100110110",
86115=>"001001011",
86116=>"000000000",
86117=>"010001001",
86118=>"100011011",
86119=>"000011011",
86120=>"010001111",
86121=>"110000000",
86122=>"111001011",
86123=>"010111111",
86124=>"111001111",
86125=>"100100100",
86126=>"000110010",
86127=>"111100000",
86128=>"001001001",
86129=>"010111001",
86130=>"011011000",
86131=>"001001111",
86132=>"001000110",
86133=>"000100100",
86134=>"000100100",
86135=>"110111000",
86136=>"110110000",
86137=>"110101100",
86138=>"010011011",
86139=>"110000000",
86140=>"110010000",
86141=>"000000011",
86142=>"110010110",
86143=>"000110011",
86144=>"101110010",
86145=>"011000010",
86146=>"110111000",
86147=>"000000000",
86148=>"001001000",
86149=>"110110101",
86150=>"111001110",
86151=>"110100100",
86152=>"011001001",
86153=>"000001001",
86154=>"001011111",
86155=>"100110111",
86156=>"100101000",
86157=>"100110100",
86158=>"000111101",
86159=>"000000001",
86160=>"101001001",
86161=>"001000000",
86162=>"111111011",
86163=>"001000000",
86164=>"100111001",
86165=>"000010110",
86166=>"001110010",
86167=>"101101111",
86168=>"000001100",
86169=>"011110111",
86170=>"111101111",
86171=>"100111011",
86172=>"100110111",
86173=>"100110110",
86174=>"010001111",
86175=>"101100101",
86176=>"001110100",
86177=>"110100100",
86178=>"001001111",
86179=>"011110111",
86180=>"111001111",
86181=>"100110010",
86182=>"000000111",
86183=>"111011001",
86184=>"110100000",
86185=>"100010111",
86186=>"011111111",
86187=>"000000000",
86188=>"010100110",
86189=>"111101100",
86190=>"000000010",
86191=>"100010011",
86192=>"000100010",
86193=>"110100101",
86194=>"001000000",
86195=>"010000010",
86196=>"100100000",
86197=>"000000111",
86198=>"011110111",
86199=>"001001101",
86200=>"111000000",
86201=>"000100000",
86202=>"011001100",
86203=>"111000011",
86204=>"000101111",
86205=>"110111111",
86206=>"111101000",
86207=>"010111011",
86208=>"100100110",
86209=>"111010110",
86210=>"000110011",
86211=>"011001000",
86212=>"100100000",
86213=>"000110101",
86214=>"110100000",
86215=>"110010100",
86216=>"100110001",
86217=>"010000000",
86218=>"011111000",
86219=>"010011011",
86220=>"111000001",
86221=>"100101101",
86222=>"111100100",
86223=>"100000111",
86224=>"110001111",
86225=>"011111111",
86226=>"100100110",
86227=>"000001001",
86228=>"000110111",
86229=>"000000000",
86230=>"001111111",
86231=>"111011111",
86232=>"011001011",
86233=>"000011011",
86234=>"000101110",
86235=>"100110110",
86236=>"011011011",
86237=>"100001011",
86238=>"000101111",
86239=>"100000000",
86240=>"000011011",
86241=>"010110110",
86242=>"110111110",
86243=>"100100001",
86244=>"010010010",
86245=>"001001001",
86246=>"100001001",
86247=>"111001001",
86248=>"110111011",
86249=>"100110111",
86250=>"110110110",
86251=>"110111101",
86252=>"010110010",
86253=>"000000011",
86254=>"000100000",
86255=>"111110001",
86256=>"011001111",
86257=>"101000100",
86258=>"111101100",
86259=>"011001011",
86260=>"000000010",
86261=>"110110111",
86262=>"100110100",
86263=>"010110101",
86264=>"110100100",
86265=>"010011010",
86266=>"100100100",
86267=>"010000000",
86268=>"111111011",
86269=>"011111111",
86270=>"000001101",
86271=>"110111001",
86272=>"011011011",
86273=>"000110110",
86274=>"101000000",
86275=>"010111111",
86276=>"011000000",
86277=>"110010000",
86278=>"100010101",
86279=>"000101111",
86280=>"010110100",
86281=>"100111101",
86282=>"000001001",
86283=>"000000010",
86284=>"111011000",
86285=>"011000111",
86286=>"110110110",
86287=>"000110101",
86288=>"110110000",
86289=>"001101111",
86290=>"101000010",
86291=>"000010110",
86292=>"111000010",
86293=>"111000000",
86294=>"000101101",
86295=>"010111011",
86296=>"000000000",
86297=>"010000010",
86298=>"000000010",
86299=>"000111101",
86300=>"000100010",
86301=>"010010000",
86302=>"000000000",
86303=>"101000101",
86304=>"011101111",
86305=>"110110111",
86306=>"001000101",
86307=>"000000000",
86308=>"001100101",
86309=>"000000000",
86310=>"110111111",
86311=>"111111011",
86312=>"011010011",
86313=>"110111111",
86314=>"110011110",
86315=>"000100110",
86316=>"011111011",
86317=>"000111011",
86318=>"010111101",
86319=>"011000000",
86320=>"110111001",
86321=>"101110100",
86322=>"101110000",
86323=>"110101010",
86324=>"000001001",
86325=>"010110110",
86326=>"000100100",
86327=>"000010111",
86328=>"011111000",
86329=>"111010000",
86330=>"101101100",
86331=>"110111111",
86332=>"100001001",
86333=>"001101000",
86334=>"001000000",
86335=>"000101001",
86336=>"001101110",
86337=>"111111011",
86338=>"100010110",
86339=>"001001101",
86340=>"111000000",
86341=>"011000000",
86342=>"000100100",
86343=>"111111010",
86344=>"010100000",
86345=>"011111111",
86346=>"000110100",
86347=>"000101111",
86348=>"101000111",
86349=>"100001001",
86350=>"101001000",
86351=>"100110000",
86352=>"001101111",
86353=>"011000000",
86354=>"111111010",
86355=>"011011000",
86356=>"111111110",
86357=>"000101100",
86358=>"100101100",
86359=>"000000000",
86360=>"011101010",
86361=>"101100101",
86362=>"001000011",
86363=>"000000111",
86364=>"010011001",
86365=>"000000000",
86366=>"111111111",
86367=>"100100100",
86368=>"111110111",
86369=>"111111011",
86370=>"101000011",
86371=>"000100110",
86372=>"100000000",
86373=>"000001000",
86374=>"010011010",
86375=>"000000000",
86376=>"011101101",
86377=>"111111101",
86378=>"001101000",
86379=>"111111100",
86380=>"111001000",
86381=>"111000110",
86382=>"000000010",
86383=>"110111111",
86384=>"001001100",
86385=>"000111101",
86386=>"000001011",
86387=>"101000111",
86388=>"111111111",
86389=>"111000100",
86390=>"000110111",
86391=>"111111111",
86392=>"110010110",
86393=>"000001000",
86394=>"101110010",
86395=>"111000000",
86396=>"000011001",
86397=>"110110000",
86398=>"110101111",
86399=>"111000001",
86400=>"010010000",
86401=>"010000010",
86402=>"110010100",
86403=>"011110001",
86404=>"011111000",
86405=>"000010111",
86406=>"010001000",
86407=>"001000000",
86408=>"100101001",
86409=>"001010010",
86410=>"001000111",
86411=>"111011111",
86412=>"110000000",
86413=>"010010110",
86414=>"000110111",
86415=>"000110000",
86416=>"101111001",
86417=>"110000100",
86418=>"011000001",
86419=>"010100101",
86420=>"000100011",
86421=>"101111111",
86422=>"000010110",
86423=>"000000110",
86424=>"111010000",
86425=>"111001011",
86426=>"111101000",
86427=>"000010000",
86428=>"011110000",
86429=>"000111010",
86430=>"011111000",
86431=>"000111000",
86432=>"000100000",
86433=>"000100111",
86434=>"101001000",
86435=>"000000110",
86436=>"110111010",
86437=>"100000010",
86438=>"000000100",
86439=>"101100000",
86440=>"010011111",
86441=>"000000010",
86442=>"111101000",
86443=>"000101110",
86444=>"010111010",
86445=>"000001101",
86446=>"000110110",
86447=>"100000011",
86448=>"111010010",
86449=>"101001100",
86450=>"111000000",
86451=>"001001001",
86452=>"001001101",
86453=>"010010111",
86454=>"111111010",
86455=>"000000010",
86456=>"001100010",
86457=>"011011110",
86458=>"000000110",
86459=>"000111000",
86460=>"111010111",
86461=>"111011111",
86462=>"000011000",
86463=>"101001100",
86464=>"000111010",
86465=>"000111101",
86466=>"010110111",
86467=>"000001001",
86468=>"111010000",
86469=>"011101110",
86470=>"010111110",
86471=>"111110110",
86472=>"111010111",
86473=>"000000111",
86474=>"111111011",
86475=>"100101101",
86476=>"000001010",
86477=>"000100110",
86478=>"000101111",
86479=>"110101101",
86480=>"010010011",
86481=>"010011011",
86482=>"100001111",
86483=>"010010101",
86484=>"111011111",
86485=>"000101011",
86486=>"100001010",
86487=>"000110000",
86488=>"000011100",
86489=>"011000000",
86490=>"000001000",
86491=>"111000000",
86492=>"100101001",
86493=>"000000111",
86494=>"010010001",
86495=>"010010010",
86496=>"101000000",
86497=>"111100010",
86498=>"110001000",
86499=>"001001010",
86500=>"000000010",
86501=>"101100000",
86502=>"010000011",
86503=>"000011110",
86504=>"111101111",
86505=>"100101101",
86506=>"000100100",
86507=>"111011101",
86508=>"010010000",
86509=>"000100100",
86510=>"111010010",
86511=>"000001001",
86512=>"000101111",
86513=>"000111011",
86514=>"010011011",
86515=>"001001100",
86516=>"000110110",
86517=>"111000111",
86518=>"000000010",
86519=>"010000000",
86520=>"010111011",
86521=>"111101111",
86522=>"011111110",
86523=>"111111110",
86524=>"000110101",
86525=>"000000101",
86526=>"101101000",
86527=>"000000110",
86528=>"011001110",
86529=>"000000000",
86530=>"111000100",
86531=>"000100010",
86532=>"000000000",
86533=>"001000100",
86534=>"000111110",
86535=>"000000111",
86536=>"101011000",
86537=>"000011111",
86538=>"000110001",
86539=>"000010011",
86540=>"001101101",
86541=>"000010111",
86542=>"000000011",
86543=>"110000000",
86544=>"111000100",
86545=>"111000000",
86546=>"111000000",
86547=>"000000010",
86548=>"110100000",
86549=>"111100000",
86550=>"101101111",
86551=>"100000111",
86552=>"000000000",
86553=>"011111101",
86554=>"001011111",
86555=>"011000100",
86556=>"010000001",
86557=>"110011000",
86558=>"010010000",
86559=>"000000011",
86560=>"001110111",
86561=>"110000000",
86562=>"010111000",
86563=>"000111000",
86564=>"100110110",
86565=>"001000000",
86566=>"000110111",
86567=>"000100010",
86568=>"011101101",
86569=>"100000001",
86570=>"000000011",
86571=>"000100000",
86572=>"111111111",
86573=>"010111100",
86574=>"111111111",
86575=>"111101101",
86576=>"000010000",
86577=>"010001011",
86578=>"000001001",
86579=>"000100000",
86580=>"000011010",
86581=>"100000110",
86582=>"011011110",
86583=>"101000000",
86584=>"000000000",
86585=>"110110111",
86586=>"000000101",
86587=>"000000010",
86588=>"000110111",
86589=>"111111010",
86590=>"000010000",
86591=>"011001001",
86592=>"100110111",
86593=>"101010000",
86594=>"000111000",
86595=>"000101110",
86596=>"111111001",
86597=>"000000000",
86598=>"101111111",
86599=>"111111000",
86600=>"000010110",
86601=>"111100000",
86602=>"000000000",
86603=>"110010111",
86604=>"111101000",
86605=>"100001001",
86606=>"000100110",
86607=>"111111001",
86608=>"101001000",
86609=>"111000000",
86610=>"110110111",
86611=>"001001000",
86612=>"010110000",
86613=>"111011001",
86614=>"010000011",
86615=>"001000100",
86616=>"000110110",
86617=>"000001001",
86618=>"111000000",
86619=>"000111110",
86620=>"111000000",
86621=>"000001001",
86622=>"111111000",
86623=>"110110110",
86624=>"000000111",
86625=>"111110101",
86626=>"111000000",
86627=>"110111110",
86628=>"000100110",
86629=>"010000000",
86630=>"010111110",
86631=>"101110010",
86632=>"010000001",
86633=>"011000111",
86634=>"111111011",
86635=>"000000000",
86636=>"111111000",
86637=>"111100111",
86638=>"011010000",
86639=>"000000000",
86640=>"000001111",
86641=>"000000010",
86642=>"000100111",
86643=>"000000010",
86644=>"100101000",
86645=>"000000000",
86646=>"111010001",
86647=>"111001100",
86648=>"000111000",
86649=>"000010011",
86650=>"100111110",
86651=>"000000000",
86652=>"110110101",
86653=>"100100000",
86654=>"000100000",
86655=>"111101000",
86656=>"000000000",
86657=>"000000110",
86658=>"010010000",
86659=>"000000000",
86660=>"110111111",
86661=>"011011000",
86662=>"110110100",
86663=>"011110110",
86664=>"110110110",
86665=>"100000010",
86666=>"000100111",
86667=>"011000000",
86668=>"111000000",
86669=>"000000010",
86670=>"000101100",
86671=>"001011100",
86672=>"000111010",
86673=>"000000111",
86674=>"000000001",
86675=>"111001000",
86676=>"100110111",
86677=>"000010000",
86678=>"111110010",
86679=>"000001100",
86680=>"010110000",
86681=>"111101001",
86682=>"110000110",
86683=>"111101010",
86684=>"111001110",
86685=>"000100100",
86686=>"111000000",
86687=>"100000000",
86688=>"001010010",
86689=>"010010000",
86690=>"101111111",
86691=>"100000000",
86692=>"111010100",
86693=>"000111111",
86694=>"100111110",
86695=>"011111000",
86696=>"001110111",
86697=>"100100000",
86698=>"111000000",
86699=>"111100000",
86700=>"101001000",
86701=>"101100100",
86702=>"100000000",
86703=>"111110111",
86704=>"000000000",
86705=>"001111101",
86706=>"001111111",
86707=>"000000100",
86708=>"000010110",
86709=>"011111000",
86710=>"011100100",
86711=>"000100101",
86712=>"100100011",
86713=>"101111011",
86714=>"000011000",
86715=>"111000010",
86716=>"110000000",
86717=>"111110000",
86718=>"100100100",
86719=>"000000011",
86720=>"101100001",
86721=>"010010000",
86722=>"000000101",
86723=>"000111111",
86724=>"011010000",
86725=>"111001011",
86726=>"000110111",
86727=>"110111111",
86728=>"101100010",
86729=>"001100000",
86730=>"011000000",
86731=>"111000000",
86732=>"011011001",
86733=>"111101000",
86734=>"100010000",
86735=>"110000101",
86736=>"000010111",
86737=>"010110111",
86738=>"111010100",
86739=>"111000000",
86740=>"000111000",
86741=>"100100000",
86742=>"000011010",
86743=>"111111111",
86744=>"011000001",
86745=>"100000110",
86746=>"101010011",
86747=>"111000000",
86748=>"110100111",
86749=>"000000000",
86750=>"010111111",
86751=>"011000000",
86752=>"111010000",
86753=>"101100110",
86754=>"010111110",
86755=>"011001111",
86756=>"101000000",
86757=>"001111111",
86758=>"000010111",
86759=>"010011111",
86760=>"000010111",
86761=>"101110111",
86762=>"000111100",
86763=>"111101100",
86764=>"000000000",
86765=>"000010111",
86766=>"011000010",
86767=>"000000000",
86768=>"011011010",
86769=>"011100110",
86770=>"001000010",
86771=>"000110101",
86772=>"100100111",
86773=>"111111111",
86774=>"000000010",
86775=>"000010001",
86776=>"111011000",
86777=>"001010011",
86778=>"000001101",
86779=>"100111111",
86780=>"111000000",
86781=>"111100000",
86782=>"111001000",
86783=>"111011001",
86784=>"011011000",
86785=>"111000001",
86786=>"101000001",
86787=>"110000111",
86788=>"100111111",
86789=>"000000110",
86790=>"000111110",
86791=>"001101101",
86792=>"000001000",
86793=>"111000100",
86794=>"000010000",
86795=>"111101101",
86796=>"101000000",
86797=>"000000001",
86798=>"000000011",
86799=>"000001101",
86800=>"011010111",
86801=>"111100000",
86802=>"010110111",
86803=>"000001010",
86804=>"110111111",
86805=>"111111111",
86806=>"110000101",
86807=>"000111111",
86808=>"000001100",
86809=>"111111111",
86810=>"000101000",
86811=>"101000001",
86812=>"110110101",
86813=>"000000111",
86814=>"000111011",
86815=>"000000111",
86816=>"111000000",
86817=>"110100110",
86818=>"000000000",
86819=>"111111000",
86820=>"010111100",
86821=>"100111111",
86822=>"101000000",
86823=>"010010000",
86824=>"110100101",
86825=>"000001111",
86826=>"001111000",
86827=>"101000000",
86828=>"111111111",
86829=>"101011000",
86830=>"111001001",
86831=>"010000100",
86832=>"010101000",
86833=>"100100110",
86834=>"111100110",
86835=>"111101111",
86836=>"000010111",
86837=>"111000000",
86838=>"111111011",
86839=>"101000011",
86840=>"001000000",
86841=>"100100010",
86842=>"000001111",
86843=>"111101101",
86844=>"010011011",
86845=>"111111001",
86846=>"100000000",
86847=>"001100110",
86848=>"111100101",
86849=>"000111111",
86850=>"111111000",
86851=>"000110011",
86852=>"111101111",
86853=>"111000010",
86854=>"010010111",
86855=>"010110110",
86856=>"111101100",
86857=>"001000001",
86858=>"110001001",
86859=>"000011111",
86860=>"000000000",
86861=>"101101101",
86862=>"010111011",
86863=>"000000000",
86864=>"000000111",
86865=>"111000000",
86866=>"011000111",
86867=>"000011100",
86868=>"101000000",
86869=>"111101100",
86870=>"100111111",
86871=>"101111111",
86872=>"111000001",
86873=>"100100111",
86874=>"100101101",
86875=>"010011111",
86876=>"111000000",
86877=>"001001001",
86878=>"111101111",
86879=>"101110110",
86880=>"000111110",
86881=>"000011011",
86882=>"101000101",
86883=>"100101001",
86884=>"100110000",
86885=>"011000001",
86886=>"111110010",
86887=>"000011100",
86888=>"000000010",
86889=>"010100001",
86890=>"111000010",
86891=>"010000001",
86892=>"101000001",
86893=>"010111111",
86894=>"000010111",
86895=>"001000001",
86896=>"100100111",
86897=>"111111001",
86898=>"111011110",
86899=>"000000000",
86900=>"111101101",
86901=>"101001111",
86902=>"000011010",
86903=>"001000000",
86904=>"111000000",
86905=>"110111111",
86906=>"000000111",
86907=>"001001111",
86908=>"100110010",
86909=>"000100000",
86910=>"000000000",
86911=>"001000001",
86912=>"111010000",
86913=>"100101000",
86914=>"010000000",
86915=>"000000000",
86916=>"001000000",
86917=>"000010000",
86918=>"001011111",
86919=>"001010001",
86920=>"011111011",
86921=>"111111010",
86922=>"000101000",
86923=>"110000111",
86924=>"000000000",
86925=>"111111111",
86926=>"011101000",
86927=>"000000101",
86928=>"100100100",
86929=>"101001101",
86930=>"011010000",
86931=>"101000111",
86932=>"111000000",
86933=>"000010011",
86934=>"110110000",
86935=>"110100100",
86936=>"101110010",
86937=>"111111110",
86938=>"111010110",
86939=>"000000000",
86940=>"011111011",
86941=>"111010000",
86942=>"111010010",
86943=>"000000000",
86944=>"010100001",
86945=>"101000000",
86946=>"111101000",
86947=>"110000001",
86948=>"000000111",
86949=>"110110010",
86950=>"111001101",
86951=>"011101000",
86952=>"111110111",
86953=>"111011000",
86954=>"010000101",
86955=>"000001101",
86956=>"010001111",
86957=>"000000000",
86958=>"111111111",
86959=>"110111111",
86960=>"000000101",
86961=>"001100110",
86962=>"000000000",
86963=>"000000010",
86964=>"000000101",
86965=>"000000000",
86966=>"110000100",
86967=>"001000010",
86968=>"011110010",
86969=>"110010000",
86970=>"011001101",
86971=>"000000011",
86972=>"110101100",
86973=>"110101111",
86974=>"100000000",
86975=>"111000000",
86976=>"011111010",
86977=>"000111010",
86978=>"000010111",
86979=>"001001001",
86980=>"011000000",
86981=>"100010001",
86982=>"011000000",
86983=>"111111110",
86984=>"011010000",
86985=>"101101111",
86986=>"111000010",
86987=>"100110000",
86988=>"000011111",
86989=>"000110010",
86990=>"000111111",
86991=>"000000000",
86992=>"000000000",
86993=>"001011011",
86994=>"010111111",
86995=>"000100001",
86996=>"000010110",
86997=>"110100101",
86998=>"110100000",
86999=>"000000000",
87000=>"111111000",
87001=>"000101101",
87002=>"111011000",
87003=>"000000100",
87004=>"001000001",
87005=>"100111100",
87006=>"111111111",
87007=>"010110111",
87008=>"100000000",
87009=>"010000000",
87010=>"000000100",
87011=>"001111111",
87012=>"000011111",
87013=>"010000111",
87014=>"111101111",
87015=>"011000101",
87016=>"101100111",
87017=>"111000010",
87018=>"000111011",
87019=>"111101000",
87020=>"000000000",
87021=>"101101000",
87022=>"000000000",
87023=>"111000000",
87024=>"111101101",
87025=>"000000100",
87026=>"000000010",
87027=>"000000111",
87028=>"111111001",
87029=>"100111011",
87030=>"110101100",
87031=>"000000000",
87032=>"000111000",
87033=>"101000010",
87034=>"010111000",
87035=>"111111101",
87036=>"111010001",
87037=>"000011011",
87038=>"010000000",
87039=>"000010000",
87040=>"100110010",
87041=>"000101000",
87042=>"011001000",
87043=>"101000001",
87044=>"111110001",
87045=>"111001001",
87046=>"101101111",
87047=>"111111000",
87048=>"010001001",
87049=>"110000000",
87050=>"011111110",
87051=>"111110110",
87052=>"000000010",
87053=>"000010010",
87054=>"001110110",
87055=>"000000010",
87056=>"111110110",
87057=>"000000110",
87058=>"000000000",
87059=>"110100110",
87060=>"000111111",
87061=>"111110000",
87062=>"111110111",
87063=>"111000101",
87064=>"111000000",
87065=>"111000001",
87066=>"010000010",
87067=>"000000000",
87068=>"001000110",
87069=>"100000010",
87070=>"000001000",
87071=>"101101111",
87072=>"111111111",
87073=>"111111111",
87074=>"000010000",
87075=>"001000011",
87076=>"100010000",
87077=>"100000110",
87078=>"010000000",
87079=>"001000000",
87080=>"000001000",
87081=>"111111111",
87082=>"101000111",
87083=>"000000000",
87084=>"000001001",
87085=>"000000000",
87086=>"110110111",
87087=>"111111010",
87088=>"111111111",
87089=>"111110011",
87090=>"001000000",
87091=>"000011010",
87092=>"111111111",
87093=>"001011010",
87094=>"100001010",
87095=>"100101101",
87096=>"010111000",
87097=>"000000111",
87098=>"111111010",
87099=>"101000001",
87100=>"000001100",
87101=>"101111111",
87102=>"100001111",
87103=>"100100001",
87104=>"001111110",
87105=>"110000000",
87106=>"111000001",
87107=>"011011001",
87108=>"001111111",
87109=>"111111010",
87110=>"000000000",
87111=>"010010111",
87112=>"000000000",
87113=>"000000111",
87114=>"000111110",
87115=>"110111111",
87116=>"111001000",
87117=>"011110001",
87118=>"110110001",
87119=>"011111111",
87120=>"101000001",
87121=>"111111111",
87122=>"011101111",
87123=>"111110001",
87124=>"101000101",
87125=>"100111001",
87126=>"011000100",
87127=>"111000000",
87128=>"111010111",
87129=>"000110111",
87130=>"101001101",
87131=>"111111111",
87132=>"000110010",
87133=>"000111000",
87134=>"000000000",
87135=>"110101001",
87136=>"000000000",
87137=>"111000000",
87138=>"000110011",
87139=>"101101001",
87140=>"100110111",
87141=>"000000101",
87142=>"101000101",
87143=>"110000000",
87144=>"110111001",
87145=>"000000000",
87146=>"000000100",
87147=>"110000101",
87148=>"111111010",
87149=>"000111110",
87150=>"101001000",
87151=>"000010000",
87152=>"011110110",
87153=>"000000001",
87154=>"110100100",
87155=>"000000000",
87156=>"000000000",
87157=>"110000000",
87158=>"000000000",
87159=>"110100000",
87160=>"001010000",
87161=>"110000000",
87162=>"000101110",
87163=>"000000010",
87164=>"000000100",
87165=>"101011110",
87166=>"111010000",
87167=>"001010100",
87168=>"111000001",
87169=>"101110111",
87170=>"000011111",
87171=>"000111100",
87172=>"000111111",
87173=>"000000000",
87174=>"011100111",
87175=>"001001111",
87176=>"011011011",
87177=>"010010110",
87178=>"011111011",
87179=>"111000111",
87180=>"111111000",
87181=>"000011000",
87182=>"000110110",
87183=>"101110110",
87184=>"001000100",
87185=>"111111111",
87186=>"111110000",
87187=>"000011111",
87188=>"000011111",
87189=>"111111111",
87190=>"000110110",
87191=>"110111110",
87192=>"110000101",
87193=>"111111101",
87194=>"101000100",
87195=>"000000001",
87196=>"010011010",
87197=>"000100000",
87198=>"000000000",
87199=>"001101111",
87200=>"100110000",
87201=>"000000000",
87202=>"111000000",
87203=>"010001101",
87204=>"000001111",
87205=>"100111111",
87206=>"011111001",
87207=>"001001111",
87208=>"111100111",
87209=>"000010000",
87210=>"000011011",
87211=>"001000111",
87212=>"111111101",
87213=>"000100111",
87214=>"000011011",
87215=>"110111000",
87216=>"001000000",
87217=>"100100100",
87218=>"111111111",
87219=>"100010000",
87220=>"001000000",
87221=>"000000011",
87222=>"110110000",
87223=>"100000000",
87224=>"000100001",
87225=>"000110101",
87226=>"010010110",
87227=>"000110111",
87228=>"110000000",
87229=>"111101100",
87230=>"011101110",
87231=>"110111000",
87232=>"000000101",
87233=>"101000000",
87234=>"000010101",
87235=>"110010011",
87236=>"000000000",
87237=>"100100000",
87238=>"000001111",
87239=>"111000010",
87240=>"000011100",
87241=>"111111101",
87242=>"111111111",
87243=>"100000000",
87244=>"101000000",
87245=>"000001001",
87246=>"100101101",
87247=>"111111110",
87248=>"011000001",
87249=>"111100000",
87250=>"110101111",
87251=>"001101101",
87252=>"111000001",
87253=>"010111011",
87254=>"010000000",
87255=>"110000000",
87256=>"001000000",
87257=>"001000101",
87258=>"000100111",
87259=>"000111111",
87260=>"011111000",
87261=>"010010111",
87262=>"111001000",
87263=>"010010111",
87264=>"111100110",
87265=>"000001111",
87266=>"010100010",
87267=>"111111110",
87268=>"110110000",
87269=>"111011000",
87270=>"000000000",
87271=>"100000000",
87272=>"001011010",
87273=>"000110110",
87274=>"111011101",
87275=>"001000101",
87276=>"111111111",
87277=>"101111010",
87278=>"010000011",
87279=>"010010000",
87280=>"011000100",
87281=>"011000010",
87282=>"000000000",
87283=>"000100000",
87284=>"000001011",
87285=>"101101101",
87286=>"000001101",
87287=>"010000000",
87288=>"111111000",
87289=>"100000000",
87290=>"011000001",
87291=>"110101101",
87292=>"000000101",
87293=>"111111111",
87294=>"000000001",
87295=>"001000111",
87296=>"111101101",
87297=>"110111111",
87298=>"001000001",
87299=>"100001001",
87300=>"000000000",
87301=>"100010010",
87302=>"100000000",
87303=>"000111101",
87304=>"000000000",
87305=>"110010110",
87306=>"101101000",
87307=>"000100110",
87308=>"001001001",
87309=>"100000100",
87310=>"111010111",
87311=>"110110101",
87312=>"101000000",
87313=>"110010110",
87314=>"000000100",
87315=>"000000110",
87316=>"001101001",
87317=>"111001111",
87318=>"111101111",
87319=>"000000000",
87320=>"110110000",
87321=>"101000111",
87322=>"000000000",
87323=>"100110101",
87324=>"000101111",
87325=>"100000011",
87326=>"000011111",
87327=>"110100001",
87328=>"101101100",
87329=>"000000000",
87330=>"110110010",
87331=>"000110000",
87332=>"111111111",
87333=>"000010000",
87334=>"100000001",
87335=>"100110100",
87336=>"111101111",
87337=>"001001010",
87338=>"000010110",
87339=>"011011001",
87340=>"110100001",
87341=>"110011011",
87342=>"000011011",
87343=>"011110111",
87344=>"000000110",
87345=>"100100001",
87346=>"010001100",
87347=>"001111110",
87348=>"001000100",
87349=>"000010011",
87350=>"000100111",
87351=>"110111100",
87352=>"001001100",
87353=>"100100110",
87354=>"000000000",
87355=>"100010001",
87356=>"001001001",
87357=>"000000000",
87358=>"011011011",
87359=>"100001000",
87360=>"111001011",
87361=>"000001101",
87362=>"011000000",
87363=>"011011001",
87364=>"000010110",
87365=>"000010010",
87366=>"000100100",
87367=>"000000011",
87368=>"100111101",
87369=>"000100000",
87370=>"111111111",
87371=>"100000001",
87372=>"001001011",
87373=>"111100111",
87374=>"111011111",
87375=>"001011001",
87376=>"011001001",
87377=>"000000000",
87378=>"111110001",
87379=>"101100100",
87380=>"001000000",
87381=>"011010011",
87382=>"111101100",
87383=>"010011110",
87384=>"111110110",
87385=>"000100100",
87386=>"010000100",
87387=>"001101000",
87388=>"110110100",
87389=>"000100100",
87390=>"101001011",
87391=>"001001101",
87392=>"100110110",
87393=>"101111101",
87394=>"101001011",
87395=>"110110110",
87396=>"000100100",
87397=>"111111111",
87398=>"000100000",
87399=>"000000000",
87400=>"101111101",
87401=>"000111111",
87402=>"101011000",
87403=>"011101011",
87404=>"000001001",
87405=>"101000101",
87406=>"001000100",
87407=>"100101110",
87408=>"011010011",
87409=>"000001000",
87410=>"111011011",
87411=>"011111001",
87412=>"011111101",
87413=>"011011010",
87414=>"100100000",
87415=>"000000011",
87416=>"001011001",
87417=>"100100100",
87418=>"111111111",
87419=>"011000011",
87420=>"000000000",
87421=>"000000000",
87422=>"000000001",
87423=>"111000001",
87424=>"101011011",
87425=>"101001101",
87426=>"100101000",
87427=>"000011001",
87428=>"011001100",
87429=>"101111111",
87430=>"001101111",
87431=>"110110001",
87432=>"111111111",
87433=>"100000000",
87434=>"111001001",
87435=>"001000001",
87436=>"101101011",
87437=>"001101001",
87438=>"000000000",
87439=>"000010000",
87440=>"111111111",
87441=>"111101101",
87442=>"100100100",
87443=>"011001000",
87444=>"100000000",
87445=>"101011011",
87446=>"001001101",
87447=>"100100100",
87448=>"001000000",
87449=>"000011000",
87450=>"001001001",
87451=>"111011011",
87452=>"000100000",
87453=>"100000111",
87454=>"101111001",
87455=>"011011011",
87456=>"111101101",
87457=>"111000111",
87458=>"000000001",
87459=>"011001101",
87460=>"101001101",
87461=>"000000100",
87462=>"100110000",
87463=>"100101100",
87464=>"000110011",
87465=>"110100001",
87466=>"011001011",
87467=>"101000001",
87468=>"000000011",
87469=>"001001001",
87470=>"001001001",
87471=>"000000000",
87472=>"010100011",
87473=>"111011110",
87474=>"000000001",
87475=>"000001000",
87476=>"111100110",
87477=>"011001100",
87478=>"100110111",
87479=>"000101011",
87480=>"110100100",
87481=>"110010000",
87482=>"100110100",
87483=>"001001001",
87484=>"001101101",
87485=>"001001001",
87486=>"111000111",
87487=>"000011100",
87488=>"000011011",
87489=>"100100100",
87490=>"001000011",
87491=>"111000001",
87492=>"000000000",
87493=>"000001011",
87494=>"101101100",
87495=>"100111111",
87496=>"000100100",
87497=>"101010011",
87498=>"011101001",
87499=>"100011111",
87500=>"111111000",
87501=>"111100100",
87502=>"110100100",
87503=>"111101000",
87504=>"101001101",
87505=>"001010001",
87506=>"100101001",
87507=>"000000000",
87508=>"001101111",
87509=>"000000011",
87510=>"001001001",
87511=>"101111101",
87512=>"110000100",
87513=>"100100100",
87514=>"001001000",
87515=>"001000000",
87516=>"101001001",
87517=>"111000000",
87518=>"100100000",
87519=>"001000000",
87520=>"011001000",
87521=>"011000000",
87522=>"101011001",
87523=>"111100000",
87524=>"001000000",
87525=>"101100001",
87526=>"100000110",
87527=>"100001111",
87528=>"110011111",
87529=>"000111110",
87530=>"100000011",
87531=>"000010011",
87532=>"100010011",
87533=>"100100110",
87534=>"000000000",
87535=>"000000000",
87536=>"010011101",
87537=>"110111011",
87538=>"100111111",
87539=>"000000000",
87540=>"010110110",
87541=>"001011011",
87542=>"011101100",
87543=>"110000000",
87544=>"000001011",
87545=>"100111100",
87546=>"000001001",
87547=>"101111101",
87548=>"001001101",
87549=>"000001001",
87550=>"001010110",
87551=>"101111001",
87552=>"110011100",
87553=>"010000010",
87554=>"101000111",
87555=>"000000111",
87556=>"000000100",
87557=>"010001111",
87558=>"000110011",
87559=>"010111110",
87560=>"111001000",
87561=>"101000101",
87562=>"110011000",
87563=>"000011111",
87564=>"000000001",
87565=>"000110010",
87566=>"000101000",
87567=>"111110010",
87568=>"010110000",
87569=>"010111011",
87570=>"110000001",
87571=>"000000101",
87572=>"100100101",
87573=>"000000111",
87574=>"111111100",
87575=>"010010111",
87576=>"101000000",
87577=>"001111001",
87578=>"000000000",
87579=>"111111000",
87580=>"011010110",
87581=>"111001000",
87582=>"111111000",
87583=>"101111110",
87584=>"101101101",
87585=>"000101111",
87586=>"100000110",
87587=>"000000111",
87588=>"110100100",
87589=>"011010101",
87590=>"100110010",
87591=>"000111010",
87592=>"000010011",
87593=>"000111110",
87594=>"000010000",
87595=>"100111110",
87596=>"000111111",
87597=>"111110111",
87598=>"010000011",
87599=>"001001000",
87600=>"110111111",
87601=>"110111100",
87602=>"111001101",
87603=>"001101000",
87604=>"111111000",
87605=>"111100000",
87606=>"011010010",
87607=>"101000000",
87608=>"000000011",
87609=>"111000000",
87610=>"101000100",
87611=>"000000000",
87612=>"100110110",
87613=>"010000000",
87614=>"000000000",
87615=>"001011101",
87616=>"011001101",
87617=>"001111000",
87618=>"100001101",
87619=>"110011111",
87620=>"000000000",
87621=>"100001000",
87622=>"011001000",
87623=>"111111111",
87624=>"110100011",
87625=>"000001000",
87626=>"111101000",
87627=>"000010000",
87628=>"100010010",
87629=>"011011010",
87630=>"000111011",
87631=>"000110111",
87632=>"001010010",
87633=>"010010101",
87634=>"011111000",
87635=>"000001000",
87636=>"000100111",
87637=>"111100000",
87638=>"011011010",
87639=>"111101111",
87640=>"101000110",
87641=>"010000001",
87642=>"100100011",
87643=>"110111110",
87644=>"110000000",
87645=>"000001000",
87646=>"011000101",
87647=>"010100000",
87648=>"000111111",
87649=>"011000111",
87650=>"101111111",
87651=>"010000100",
87652=>"000111100",
87653=>"110000100",
87654=>"100000111",
87655=>"100000000",
87656=>"000101110",
87657=>"111100000",
87658=>"010000111",
87659=>"011010111",
87660=>"011000000",
87661=>"101110101",
87662=>"011101111",
87663=>"111110111",
87664=>"000011011",
87665=>"000000000",
87666=>"110011000",
87667=>"111011010",
87668=>"000111111",
87669=>"111000000",
87670=>"000000100",
87671=>"010111010",
87672=>"111000001",
87673=>"000010000",
87674=>"100010111",
87675=>"000000000",
87676=>"000100110",
87677=>"000100000",
87678=>"101101111",
87679=>"100001111",
87680=>"010000000",
87681=>"010000000",
87682=>"010000001",
87683=>"010001101",
87684=>"110010001",
87685=>"111101101",
87686=>"100011001",
87687=>"000000110",
87688=>"000110100",
87689=>"000111010",
87690=>"111000100",
87691=>"000110001",
87692=>"000000101",
87693=>"000010000",
87694=>"110000000",
87695=>"000000000",
87696=>"101000000",
87697=>"111000111",
87698=>"000000000",
87699=>"011000000",
87700=>"010011111",
87701=>"000101100",
87702=>"010111110",
87703=>"000010011",
87704=>"111111000",
87705=>"111011111",
87706=>"010111111",
87707=>"001001111",
87708=>"011000000",
87709=>"110000111",
87710=>"101000000",
87711=>"000111000",
87712=>"101011010",
87713=>"111101111",
87714=>"111001111",
87715=>"111000111",
87716=>"111111000",
87717=>"100011011",
87718=>"001010110",
87719=>"110000000",
87720=>"110111100",
87721=>"000000110",
87722=>"101000111",
87723=>"110110000",
87724=>"000110000",
87725=>"000000000",
87726=>"111001100",
87727=>"111111111",
87728=>"000000000",
87729=>"000000001",
87730=>"000001000",
87731=>"011001000",
87732=>"110111101",
87733=>"010000000",
87734=>"000111100",
87735=>"000000100",
87736=>"001011111",
87737=>"011110011",
87738=>"110110111",
87739=>"111000000",
87740=>"011110111",
87741=>"101101011",
87742=>"100100100",
87743=>"111011011",
87744=>"000000100",
87745=>"000000000",
87746=>"000100000",
87747=>"100000000",
87748=>"111111111",
87749=>"110110000",
87750=>"111111000",
87751=>"000000000",
87752=>"000011110",
87753=>"000000000",
87754=>"010000000",
87755=>"000111111",
87756=>"011010000",
87757=>"000011010",
87758=>"110100111",
87759=>"101101000",
87760=>"000110111",
87761=>"000111011",
87762=>"010000110",
87763=>"011111111",
87764=>"000000000",
87765=>"011000000",
87766=>"000010111",
87767=>"001000001",
87768=>"001101101",
87769=>"010100000",
87770=>"000101101",
87771=>"101000000",
87772=>"110011001",
87773=>"000010111",
87774=>"111011000",
87775=>"001011000",
87776=>"011100001",
87777=>"111111011",
87778=>"111000101",
87779=>"010001001",
87780=>"101100100",
87781=>"000000001",
87782=>"010111111",
87783=>"010011111",
87784=>"110100111",
87785=>"000100111",
87786=>"001010000",
87787=>"010000000",
87788=>"000000101",
87789=>"000000000",
87790=>"000000010",
87791=>"010000010",
87792=>"111000000",
87793=>"011011000",
87794=>"010111010",
87795=>"111111000",
87796=>"010010101",
87797=>"011001011",
87798=>"000000010",
87799=>"101110000",
87800=>"000000000",
87801=>"001001101",
87802=>"111101100",
87803=>"000000011",
87804=>"000111011",
87805=>"000000000",
87806=>"010100001",
87807=>"000111000",
87808=>"101011001",
87809=>"010101111",
87810=>"100000000",
87811=>"000000001",
87812=>"000100100",
87813=>"000000001",
87814=>"000000000",
87815=>"000111011",
87816=>"000000010",
87817=>"000100111",
87818=>"001000000",
87819=>"000000001",
87820=>"000000101",
87821=>"100111001",
87822=>"100000110",
87823=>"000000000",
87824=>"111001010",
87825=>"000000010",
87826=>"000111010",
87827=>"110111110",
87828=>"100101111",
87829=>"000100000",
87830=>"111011100",
87831=>"111111111",
87832=>"100100000",
87833=>"111001000",
87834=>"110000000",
87835=>"000001111",
87836=>"011101111",
87837=>"000000000",
87838=>"110111001",
87839=>"000010011",
87840=>"111101101",
87841=>"010001111",
87842=>"000000000",
87843=>"111101110",
87844=>"100100100",
87845=>"111110111",
87846=>"001000000",
87847=>"000000101",
87848=>"111001111",
87849=>"011001000",
87850=>"110000001",
87851=>"000000010",
87852=>"110100010",
87853=>"111010111",
87854=>"100000001",
87855=>"111110110",
87856=>"111000000",
87857=>"010100110",
87858=>"111110111",
87859=>"100101000",
87860=>"000000001",
87861=>"000000001",
87862=>"100110100",
87863=>"100110010",
87864=>"111010000",
87865=>"000000000",
87866=>"000000111",
87867=>"101111111",
87868=>"001001011",
87869=>"111111111",
87870=>"000000000",
87871=>"110111011",
87872=>"110100000",
87873=>"111001111",
87874=>"101000000",
87875=>"011011111",
87876=>"111110010",
87877=>"000000000",
87878=>"011001001",
87879=>"111111010",
87880=>"101011110",
87881=>"010000011",
87882=>"000001001",
87883=>"000000000",
87884=>"111111011",
87885=>"001001011",
87886=>"000000001",
87887=>"111110100",
87888=>"101101111",
87889=>"110111111",
87890=>"001110111",
87891=>"011000001",
87892=>"000000000",
87893=>"001001110",
87894=>"000000101",
87895=>"001111111",
87896=>"101101111",
87897=>"001101111",
87898=>"011011111",
87899=>"100000101",
87900=>"111111010",
87901=>"010001011",
87902=>"110111110",
87903=>"100100101",
87904=>"111000000",
87905=>"010000100",
87906=>"000000001",
87907=>"110010100",
87908=>"110110110",
87909=>"000001000",
87910=>"010111010",
87911=>"111110010",
87912=>"000010011",
87913=>"110101000",
87914=>"011100010",
87915=>"011001111",
87916=>"100000000",
87917=>"000001001",
87918=>"000000000",
87919=>"000000111",
87920=>"000100100",
87921=>"001000111",
87922=>"111111000",
87923=>"100000000",
87924=>"000111010",
87925=>"100000000",
87926=>"011111111",
87927=>"101001001",
87928=>"011000010",
87929=>"000011011",
87930=>"110110111",
87931=>"100110111",
87932=>"100110101",
87933=>"110000000",
87934=>"000000001",
87935=>"000000111",
87936=>"111001000",
87937=>"000101110",
87938=>"000011111",
87939=>"001110010",
87940=>"010100000",
87941=>"000000001",
87942=>"100110011",
87943=>"110010010",
87944=>"110111111",
87945=>"111000000",
87946=>"000000000",
87947=>"101101111",
87948=>"101010000",
87949=>"101000001",
87950=>"000000000",
87951=>"001000000",
87952=>"111001001",
87953=>"111110110",
87954=>"000011000",
87955=>"000000000",
87956=>"000000110",
87957=>"001000111",
87958=>"011111010",
87959=>"010100001",
87960=>"011000010",
87961=>"000110111",
87962=>"000011010",
87963=>"101100100",
87964=>"111100000",
87965=>"000110111",
87966=>"101001111",
87967=>"111001111",
87968=>"101111111",
87969=>"010111111",
87970=>"100110100",
87971=>"111000101",
87972=>"000100111",
87973=>"101001000",
87974=>"001001001",
87975=>"110111111",
87976=>"010001000",
87977=>"000011111",
87978=>"111000000",
87979=>"111000000",
87980=>"111110000",
87981=>"000000101",
87982=>"011111110",
87983=>"000000000",
87984=>"111111111",
87985=>"011001000",
87986=>"010000000",
87987=>"000000000",
87988=>"011011101",
87989=>"001000101",
87990=>"000000100",
87991=>"111100011",
87992=>"000000100",
87993=>"000110111",
87994=>"000010111",
87995=>"111010010",
87996=>"111011110",
87997=>"000010111",
87998=>"000111000",
87999=>"010111011",
88000=>"001000000",
88001=>"000000111",
88002=>"111001010",
88003=>"001001001",
88004=>"000000000",
88005=>"111000101",
88006=>"110111100",
88007=>"111111111",
88008=>"000010111",
88009=>"000001000",
88010=>"110011111",
88011=>"000000000",
88012=>"000011011",
88013=>"111111101",
88014=>"011000000",
88015=>"011110001",
88016=>"000111111",
88017=>"001001000",
88018=>"000001001",
88019=>"010101111",
88020=>"001000101",
88021=>"110110000",
88022=>"101111111",
88023=>"000000010",
88024=>"000111111",
88025=>"000111010",
88026=>"101101110",
88027=>"101000001",
88028=>"110000000",
88029=>"100010011",
88030=>"000000000",
88031=>"000001111",
88032=>"111000000",
88033=>"111101001",
88034=>"000000000",
88035=>"011010110",
88036=>"111000000",
88037=>"111001000",
88038=>"000111111",
88039=>"100111000",
88040=>"100000101",
88041=>"010111000",
88042=>"000000000",
88043=>"111000000",
88044=>"000000011",
88045=>"101001101",
88046=>"101001001",
88047=>"000000110",
88048=>"100110101",
88049=>"111100110",
88050=>"011011011",
88051=>"100000011",
88052=>"001111110",
88053=>"000000000",
88054=>"000000110",
88055=>"100010000",
88056=>"001111111",
88057=>"000000011",
88058=>"111100111",
88059=>"000000010",
88060=>"111111010",
88061=>"111101100",
88062=>"001011001",
88063=>"100000000",
88064=>"001000111",
88065=>"110100111",
88066=>"001000111",
88067=>"010101100",
88068=>"110100100",
88069=>"111111111",
88070=>"000101001",
88071=>"011001111",
88072=>"000101101",
88073=>"000011011",
88074=>"111110001",
88075=>"001011001",
88076=>"111111010",
88077=>"000000101",
88078=>"101111000",
88079=>"000001111",
88080=>"111011110",
88081=>"010010010",
88082=>"010111010",
88083=>"111110101",
88084=>"100101101",
88085=>"011011111",
88086=>"010111010",
88087=>"010111011",
88088=>"110100100",
88089=>"001111110",
88090=>"100100111",
88091=>"000011111",
88092=>"010011100",
88093=>"100101001",
88094=>"111101111",
88095=>"010111000",
88096=>"011100111",
88097=>"001011011",
88098=>"011000011",
88099=>"101101100",
88100=>"111111010",
88101=>"100111111",
88102=>"100000000",
88103=>"000011000",
88104=>"100100101",
88105=>"000101000",
88106=>"100110011",
88107=>"010000000",
88108=>"110111110",
88109=>"111111010",
88110=>"000001100",
88111=>"111101101",
88112=>"000110010",
88113=>"011011110",
88114=>"000000010",
88115=>"011000010",
88116=>"011000010",
88117=>"100010000",
88118=>"100000001",
88119=>"010111001",
88120=>"011000000",
88121=>"010000000",
88122=>"010001000",
88123=>"000000000",
88124=>"100011100",
88125=>"111111011",
88126=>"000010000",
88127=>"010111001",
88128=>"000000111",
88129=>"101011000",
88130=>"111111000",
88131=>"110111000",
88132=>"101100000",
88133=>"000000000",
88134=>"000000000",
88135=>"111010111",
88136=>"100000100",
88137=>"011010100",
88138=>"000000000",
88139=>"111101100",
88140=>"111111010",
88141=>"111100011",
88142=>"011011001",
88143=>"111010111",
88144=>"011001000",
88145=>"111111100",
88146=>"011000110",
88147=>"011011000",
88148=>"101101101",
88149=>"110100111",
88150=>"011000000",
88151=>"000111000",
88152=>"100111100",
88153=>"111111110",
88154=>"110110000",
88155=>"011111001",
88156=>"010010000",
88157=>"000000001",
88158=>"000111000",
88159=>"011111011",
88160=>"000100000",
88161=>"010110010",
88162=>"101100101",
88163=>"000110100",
88164=>"010011110",
88165=>"111010111",
88166=>"001011000",
88167=>"101111010",
88168=>"010010011",
88169=>"011000100",
88170=>"000011011",
88171=>"111000111",
88172=>"011111001",
88173=>"011011000",
88174=>"000011000",
88175=>"110000000",
88176=>"001001000",
88177=>"010101100",
88178=>"011000110",
88179=>"111101111",
88180=>"101100110",
88181=>"000000010",
88182=>"100101000",
88183=>"001100000",
88184=>"000001001",
88185=>"010110000",
88186=>"000010111",
88187=>"001001000",
88188=>"111111111",
88189=>"000110010",
88190=>"010011010",
88191=>"010111010",
88192=>"100000110",
88193=>"111111011",
88194=>"000001010",
88195=>"000000001",
88196=>"000000111",
88197=>"000010000",
88198=>"000010011",
88199=>"011001000",
88200=>"000011000",
88201=>"010000100",
88202=>"010000000",
88203=>"011111111",
88204=>"000001000",
88205=>"000010000",
88206=>"101111111",
88207=>"000001011",
88208=>"110110111",
88209=>"000100000",
88210=>"110011011",
88211=>"111100101",
88212=>"000000000",
88213=>"000000000",
88214=>"111101000",
88215=>"010100011",
88216=>"011011000",
88217=>"000101111",
88218=>"101100100",
88219=>"000111111",
88220=>"000011011",
88221=>"100100110",
88222=>"101000010",
88223=>"101000000",
88224=>"000011001",
88225=>"101001010",
88226=>"000011011",
88227=>"100010011",
88228=>"100000000",
88229=>"100100100",
88230=>"010111011",
88231=>"000000000",
88232=>"000011000",
88233=>"100101111",
88234=>"111011010",
88235=>"000010000",
88236=>"010010011",
88237=>"101100111",
88238=>"111110100",
88239=>"000111001",
88240=>"000010111",
88241=>"110001110",
88242=>"111100100",
88243=>"000100010",
88244=>"000011010",
88245=>"000010010",
88246=>"110100000",
88247=>"000010100",
88248=>"000010001",
88249=>"001000011",
88250=>"111011000",
88251=>"111111011",
88252=>"000011011",
88253=>"111111110",
88254=>"001011111",
88255=>"010000000",
88256=>"000000000",
88257=>"010111011",
88258=>"001111111",
88259=>"100100111",
88260=>"000000101",
88261=>"110110110",
88262=>"000101111",
88263=>"000000100",
88264=>"101000000",
88265=>"100000000",
88266=>"000000010",
88267=>"000011011",
88268=>"010000000",
88269=>"100111011",
88270=>"111010011",
88271=>"000011010",
88272=>"000100000",
88273=>"011000000",
88274=>"000101000",
88275=>"111011000",
88276=>"000111111",
88277=>"110110110",
88278=>"000000000",
88279=>"011010000",
88280=>"001101111",
88281=>"000010111",
88282=>"000110010",
88283=>"000000000",
88284=>"001100011",
88285=>"101101011",
88286=>"000000011",
88287=>"111110000",
88288=>"111111111",
88289=>"101010101",
88290=>"000100101",
88291=>"001011011",
88292=>"000100000",
88293=>"111100111",
88294=>"011000000",
88295=>"011010010",
88296=>"101100100",
88297=>"000100110",
88298=>"111001000",
88299=>"000000000",
88300=>"000000110",
88301=>"111010000",
88302=>"111111010",
88303=>"010000111",
88304=>"000100100",
88305=>"111001001",
88306=>"100000000",
88307=>"010011000",
88308=>"000000000",
88309=>"000110100",
88310=>"000111110",
88311=>"010100000",
88312=>"000010010",
88313=>"000100000",
88314=>"000111011",
88315=>"111001111",
88316=>"111101111",
88317=>"100100111",
88318=>"001000001",
88319=>"000011011",
88320=>"001100101",
88321=>"000000000",
88322=>"101000001",
88323=>"101000000",
88324=>"000100001",
88325=>"010000100",
88326=>"010001111",
88327=>"001011000",
88328=>"101111000",
88329=>"111000111",
88330=>"000111111",
88331=>"111000000",
88332=>"111111011",
88333=>"000000010",
88334=>"000100100",
88335=>"001111000",
88336=>"100100111",
88337=>"000111111",
88338=>"101000000",
88339=>"111110000",
88340=>"000000000",
88341=>"010010000",
88342=>"100110100",
88343=>"100111111",
88344=>"000000101",
88345=>"110111111",
88346=>"010111111",
88347=>"000010000",
88348=>"000111111",
88349=>"000010111",
88350=>"100110011",
88351=>"011011000",
88352=>"111101100",
88353=>"101000101",
88354=>"000000000",
88355=>"101100000",
88356=>"001010011",
88357=>"111011110",
88358=>"011111001",
88359=>"101000100",
88360=>"000001101",
88361=>"101001100",
88362=>"111111100",
88363=>"111101101",
88364=>"111110110",
88365=>"110000111",
88366=>"000000111",
88367=>"010111000",
88368=>"000000101",
88369=>"100111011",
88370=>"000010111",
88371=>"111010001",
88372=>"000011000",
88373=>"111111110",
88374=>"110011011",
88375=>"110011010",
88376=>"010011010",
88377=>"000000000",
88378=>"000000000",
88379=>"000000000",
88380=>"111111001",
88381=>"111111111",
88382=>"101000000",
88383=>"010011001",
88384=>"111111001",
88385=>"011111111",
88386=>"000101000",
88387=>"001000110",
88388=>"010000000",
88389=>"000010000",
88390=>"111111001",
88391=>"000010111",
88392=>"001010000",
88393=>"000000000",
88394=>"000000000",
88395=>"000000111",
88396=>"100011011",
88397=>"110111111",
88398=>"001111001",
88399=>"000001000",
88400=>"011011011",
88401=>"010111111",
88402=>"111111100",
88403=>"000000100",
88404=>"011111000",
88405=>"101111111",
88406=>"000011011",
88407=>"111100111",
88408=>"011111011",
88409=>"100011010",
88410=>"101111001",
88411=>"111111011",
88412=>"111111010",
88413=>"000010110",
88414=>"101000100",
88415=>"101001011",
88416=>"011111001",
88417=>"100000000",
88418=>"111101111",
88419=>"110111001",
88420=>"001000001",
88421=>"111010000",
88422=>"000000000",
88423=>"100101101",
88424=>"000000000",
88425=>"000110111",
88426=>"111011011",
88427=>"111111101",
88428=>"000000001",
88429=>"000100000",
88430=>"000011010",
88431=>"000010111",
88432=>"011011011",
88433=>"111111110",
88434=>"011110110",
88435=>"000001011",
88436=>"000010010",
88437=>"001000000",
88438=>"000010001",
88439=>"000111000",
88440=>"000000000",
88441=>"101000100",
88442=>"000001111",
88443=>"001000000",
88444=>"111111000",
88445=>"000000000",
88446=>"101000101",
88447=>"010010000",
88448=>"111110101",
88449=>"000011011",
88450=>"000010000",
88451=>"000000111",
88452=>"011111111",
88453=>"111111111",
88454=>"111111101",
88455=>"111101111",
88456=>"110110110",
88457=>"101101101",
88458=>"000100111",
88459=>"100011100",
88460=>"000000000",
88461=>"111000000",
88462=>"111011100",
88463=>"001000010",
88464=>"010111110",
88465=>"101010000",
88466=>"001100110",
88467=>"001011001",
88468=>"111011011",
88469=>"100100000",
88470=>"111111000",
88471=>"111000001",
88472=>"000000101",
88473=>"000000000",
88474=>"010111010",
88475=>"111000100",
88476=>"010011111",
88477=>"111000000",
88478=>"110111101",
88479=>"010111011",
88480=>"100010010",
88481=>"111111000",
88482=>"000000000",
88483=>"101111111",
88484=>"111111011",
88485=>"110111110",
88486=>"110111110",
88487=>"101100000",
88488=>"110001111",
88489=>"010000000",
88490=>"000011000",
88491=>"000010011",
88492=>"101000100",
88493=>"011101100",
88494=>"101111110",
88495=>"101100100",
88496=>"101010000",
88497=>"111010000",
88498=>"000100100",
88499=>"001010011",
88500=>"001011001",
88501=>"000011000",
88502=>"000000000",
88503=>"100101100",
88504=>"111111011",
88505=>"001010011",
88506=>"001011111",
88507=>"111111111",
88508=>"011001111",
88509=>"000010011",
88510=>"000110100",
88511=>"000011011",
88512=>"101100000",
88513=>"100100000",
88514=>"010010011",
88515=>"110111011",
88516=>"010100111",
88517=>"000001101",
88518=>"011111001",
88519=>"111101111",
88520=>"000010000",
88521=>"010111111",
88522=>"000000010",
88523=>"001001011",
88524=>"100000000",
88525=>"011101011",
88526=>"110000111",
88527=>"100010111",
88528=>"100010000",
88529=>"100100100",
88530=>"111111101",
88531=>"111111111",
88532=>"000001001",
88533=>"100010000",
88534=>"000000000",
88535=>"000010010",
88536=>"111111000",
88537=>"011000000",
88538=>"001001000",
88539=>"001100101",
88540=>"001111100",
88541=>"010010110",
88542=>"010001011",
88543=>"111111111",
88544=>"000111111",
88545=>"000101011",
88546=>"111111100",
88547=>"001011011",
88548=>"000000000",
88549=>"111111000",
88550=>"111111010",
88551=>"111011011",
88552=>"011110010",
88553=>"000110111",
88554=>"111011000",
88555=>"010110010",
88556=>"110111111",
88557=>"101101010",
88558=>"111101101",
88559=>"011000000",
88560=>"000011000",
88561=>"100100111",
88562=>"000000100",
88563=>"001000000",
88564=>"110000110",
88565=>"010010111",
88566=>"111010100",
88567=>"100100111",
88568=>"111001010",
88569=>"001000000",
88570=>"000010010",
88571=>"010010000",
88572=>"000000000",
88573=>"000100000",
88574=>"101111111",
88575=>"101011001",
88576=>"100101100",
88577=>"000000000",
88578=>"111001000",
88579=>"011110101",
88580=>"000101011",
88581=>"101100010",
88582=>"000010110",
88583=>"001011111",
88584=>"000001111",
88585=>"000000010",
88586=>"000110111",
88587=>"000111011",
88588=>"100100000",
88589=>"110110000",
88590=>"110101101",
88591=>"001100000",
88592=>"110111011",
88593=>"111000000",
88594=>"000100000",
88595=>"101001000",
88596=>"000010000",
88597=>"110111011",
88598=>"000100000",
88599=>"111000100",
88600=>"010000000",
88601=>"000110010",
88602=>"000111111",
88603=>"000000111",
88604=>"101101001",
88605=>"011111000",
88606=>"000000011",
88607=>"111000000",
88608=>"111000000",
88609=>"000000101",
88610=>"000000000",
88611=>"001101100",
88612=>"001101111",
88613=>"000100111",
88614=>"111000111",
88615=>"000000110",
88616=>"111010110",
88617=>"000000111",
88618=>"100000111",
88619=>"100110000",
88620=>"010110101",
88621=>"010111101",
88622=>"110011010",
88623=>"010111100",
88624=>"011111001",
88625=>"000100101",
88626=>"000010001",
88627=>"000000111",
88628=>"001101110",
88629=>"000000101",
88630=>"001000000",
88631=>"000000111",
88632=>"001110111",
88633=>"101000011",
88634=>"111101100",
88635=>"000000000",
88636=>"001001111",
88637=>"000010111",
88638=>"000000000",
88639=>"000010011",
88640=>"000000110",
88641=>"000100111",
88642=>"111101101",
88643=>"100110110",
88644=>"010111000",
88645=>"000000000",
88646=>"000110000",
88647=>"010101101",
88648=>"001110111",
88649=>"000111010",
88650=>"011011111",
88651=>"111100000",
88652=>"101000010",
88653=>"110111011",
88654=>"000000100",
88655=>"101111111",
88656=>"111001001",
88657=>"111111111",
88658=>"101111111",
88659=>"000101000",
88660=>"111000000",
88661=>"011001110",
88662=>"000100100",
88663=>"000000010",
88664=>"010001000",
88665=>"010011110",
88666=>"011000100",
88667=>"100110101",
88668=>"101000111",
88669=>"010000000",
88670=>"111111110",
88671=>"011011011",
88672=>"000000000",
88673=>"110111010",
88674=>"111100000",
88675=>"111000000",
88676=>"011011101",
88677=>"000011011",
88678=>"111111110",
88679=>"000011111",
88680=>"000010011",
88681=>"111110000",
88682=>"000111111",
88683=>"111111111",
88684=>"010011111",
88685=>"111000000",
88686=>"000000000",
88687=>"000101100",
88688=>"111111101",
88689=>"000010111",
88690=>"110000000",
88691=>"110100000",
88692=>"000111101",
88693=>"000000001",
88694=>"110000000",
88695=>"000000010",
88696=>"111000010",
88697=>"111111010",
88698=>"101011001",
88699=>"000101001",
88700=>"010110000",
88701=>"110101000",
88702=>"111110000",
88703=>"111101111",
88704=>"000000000",
88705=>"000111000",
88706=>"000011011",
88707=>"000011111",
88708=>"000011110",
88709=>"000000001",
88710=>"000001111",
88711=>"000000011",
88712=>"110110100",
88713=>"000011111",
88714=>"000011100",
88715=>"100100000",
88716=>"110000000",
88717=>"100000100",
88718=>"000100111",
88719=>"000000000",
88720=>"010011111",
88721=>"000100000",
88722=>"111110010",
88723=>"111111111",
88724=>"000010001",
88725=>"111110010",
88726=>"111111111",
88727=>"000001011",
88728=>"101001101",
88729=>"110111011",
88730=>"000001000",
88731=>"111101000",
88732=>"000110111",
88733=>"000101011",
88734=>"000111011",
88735=>"010101011",
88736=>"110110110",
88737=>"000000101",
88738=>"110111111",
88739=>"110010000",
88740=>"111010011",
88741=>"000100100",
88742=>"100101001",
88743=>"010111011",
88744=>"100001000",
88745=>"000000100",
88746=>"010101000",
88747=>"101000000",
88748=>"001101101",
88749=>"000100010",
88750=>"011011000",
88751=>"111101000",
88752=>"001111111",
88753=>"011010100",
88754=>"100001000",
88755=>"000000110",
88756=>"010011101",
88757=>"100100100",
88758=>"000000000",
88759=>"100100000",
88760=>"000110011",
88761=>"000010111",
88762=>"000111111",
88763=>"010111111",
88764=>"011110010",
88765=>"111100000",
88766=>"000100110",
88767=>"000000010",
88768=>"110110010",
88769=>"100000010",
88770=>"101011001",
88771=>"111111011",
88772=>"000000111",
88773=>"111100101",
88774=>"000000110",
88775=>"000111011",
88776=>"111110110",
88777=>"101000110",
88778=>"111000000",
88779=>"111001011",
88780=>"000111111",
88781=>"000001011",
88782=>"010000000",
88783=>"100000111",
88784=>"101001010",
88785=>"000011000",
88786=>"000000011",
88787=>"000010100",
88788=>"000010000",
88789=>"111001001",
88790=>"001111111",
88791=>"000110010",
88792=>"111010110",
88793=>"000001000",
88794=>"000001000",
88795=>"111101000",
88796=>"001001011",
88797=>"100100001",
88798=>"000000000",
88799=>"001110111",
88800=>"001001011",
88801=>"011111100",
88802=>"111011000",
88803=>"011111000",
88804=>"111110110",
88805=>"000110111",
88806=>"101100111",
88807=>"000000000",
88808=>"000110011",
88809=>"010010001",
88810=>"000011111",
88811=>"111101100",
88812=>"000000011",
88813=>"000001011",
88814=>"000001000",
88815=>"001111111",
88816=>"000101111",
88817=>"000001101",
88818=>"000111010",
88819=>"000101001",
88820=>"000001110",
88821=>"111000100",
88822=>"110100000",
88823=>"000111000",
88824=>"000000000",
88825=>"011111000",
88826=>"000010010",
88827=>"110100101",
88828=>"101111111",
88829=>"110000111",
88830=>"000110111",
88831=>"010100001",
88832=>"111011011",
88833=>"111111101",
88834=>"101000101",
88835=>"110000101",
88836=>"011111001",
88837=>"110110101",
88838=>"000101010",
88839=>"000110000",
88840=>"000100111",
88841=>"111000101",
88842=>"100000000",
88843=>"000000111",
88844=>"011111111",
88845=>"000000000",
88846=>"111001100",
88847=>"000100000",
88848=>"010000000",
88849=>"000000000",
88850=>"000000111",
88851=>"011010000",
88852=>"111111110",
88853=>"000000010",
88854=>"110111111",
88855=>"100101101",
88856=>"001010000",
88857=>"111111111",
88858=>"011010100",
88859=>"110101101",
88860=>"101101101",
88861=>"001001010",
88862=>"000000011",
88863=>"001000001",
88864=>"111010101",
88865=>"110101111",
88866=>"101000111",
88867=>"010010000",
88868=>"000011011",
88869=>"111110110",
88870=>"000000000",
88871=>"001101111",
88872=>"111001101",
88873=>"001100010",
88874=>"000000000",
88875=>"010101111",
88876=>"111111011",
88877=>"101101100",
88878=>"110010101",
88879=>"000101110",
88880=>"110101001",
88881=>"011011101",
88882=>"000110000",
88883=>"110000010",
88884=>"000000010",
88885=>"010111011",
88886=>"001000000",
88887=>"000000111",
88888=>"101000100",
88889=>"000011011",
88890=>"011001010",
88891=>"111000100",
88892=>"110100101",
88893=>"111111000",
88894=>"000000001",
88895=>"100100100",
88896=>"000001111",
88897=>"111111101",
88898=>"101000111",
88899=>"011000001",
88900=>"000001000",
88901=>"001011010",
88902=>"100110010",
88903=>"001000101",
88904=>"110100010",
88905=>"010111111",
88906=>"000001101",
88907=>"001111110",
88908=>"000010010",
88909=>"010010111",
88910=>"000111010",
88911=>"001100100",
88912=>"000000000",
88913=>"111000110",
88914=>"010001000",
88915=>"011001000",
88916=>"100110101",
88917=>"101001101",
88918=>"111101000",
88919=>"111000000",
88920=>"100110111",
88921=>"000111111",
88922=>"111000000",
88923=>"001100110",
88924=>"010000000",
88925=>"010000000",
88926=>"010110010",
88927=>"100000100",
88928=>"100111111",
88929=>"000111011",
88930=>"000000001",
88931=>"111101010",
88932=>"101000000",
88933=>"111100111",
88934=>"110110010",
88935=>"000000111",
88936=>"111001011",
88937=>"000000010",
88938=>"000111111",
88939=>"010011101",
88940=>"111111001",
88941=>"000010010",
88942=>"001000100",
88943=>"000011111",
88944=>"101001011",
88945=>"000000110",
88946=>"100000000",
88947=>"000010000",
88948=>"010100100",
88949=>"101000001",
88950=>"111101010",
88951=>"000000111",
88952=>"101101101",
88953=>"111111111",
88954=>"011111110",
88955=>"010111110",
88956=>"010010100",
88957=>"110100100",
88958=>"001010111",
88959=>"101001001",
88960=>"010110000",
88961=>"111111111",
88962=>"101100000",
88963=>"000111111",
88964=>"010111111",
88965=>"111101001",
88966=>"110011001",
88967=>"000100011",
88968=>"001110110",
88969=>"111010000",
88970=>"000111101",
88971=>"000000000",
88972=>"000110110",
88973=>"001000001",
88974=>"101000101",
88975=>"000000000",
88976=>"001110110",
88977=>"111101101",
88978=>"000110000",
88979=>"000111111",
88980=>"111111000",
88981=>"110110000",
88982=>"010011111",
88983=>"000100110",
88984=>"101111000",
88985=>"000111101",
88986=>"010100111",
88987=>"000101111",
88988=>"110111011",
88989=>"010101101",
88990=>"000001100",
88991=>"000111011",
88992=>"000000111",
88993=>"101000101",
88994=>"000001000",
88995=>"000100000",
88996=>"000101100",
88997=>"000110010",
88998=>"001010110",
88999=>"000000000",
89000=>"111111100",
89001=>"000001101",
89002=>"111000001",
89003=>"111101000",
89004=>"000010111",
89005=>"101001101",
89006=>"110011111",
89007=>"000101111",
89008=>"011011101",
89009=>"001111110",
89010=>"010001000",
89011=>"000001000",
89012=>"000001011",
89013=>"101111111",
89014=>"000111011",
89015=>"111111010",
89016=>"011001100",
89017=>"001011110",
89018=>"000000101",
89019=>"010010111",
89020=>"111010000",
89021=>"111111111",
89022=>"000010100",
89023=>"000100111",
89024=>"000000000",
89025=>"011000100",
89026=>"111101101",
89027=>"000010011",
89028=>"111010000",
89029=>"001110100",
89030=>"010110111",
89031=>"111001000",
89032=>"000000000",
89033=>"000011110",
89034=>"110000011",
89035=>"100100111",
89036=>"000000100",
89037=>"001001011",
89038=>"010000000",
89039=>"111111110",
89040=>"001000000",
89041=>"011111110",
89042=>"000111111",
89043=>"001101010",
89044=>"010000000",
89045=>"000000111",
89046=>"110000100",
89047=>"000101101",
89048=>"011101000",
89049=>"001111101",
89050=>"100000001",
89051=>"100000000",
89052=>"110111001",
89053=>"101000101",
89054=>"100111111",
89055=>"111000111",
89056=>"111100100",
89057=>"111001000",
89058=>"111111110",
89059=>"111111011",
89060=>"000000000",
89061=>"110111000",
89062=>"111101101",
89063=>"100100111",
89064=>"010101010",
89065=>"000000001",
89066=>"111110000",
89067=>"001000000",
89068=>"000010011",
89069=>"101111010",
89070=>"000000011",
89071=>"000000000",
89072=>"110111100",
89073=>"111111100",
89074=>"010001111",
89075=>"000100010",
89076=>"110110110",
89077=>"101000000",
89078=>"000000000",
89079=>"111101111",
89080=>"010000000",
89081=>"100101101",
89082=>"000000000",
89083=>"000111111",
89084=>"101100111",
89085=>"110100100",
89086=>"010000110",
89087=>"111000000",
89088=>"100001001",
89089=>"111000000",
89090=>"000000000",
89091=>"110111011",
89092=>"100110111",
89093=>"001000111",
89094=>"100111111",
89095=>"101001011",
89096=>"001101101",
89097=>"000111111",
89098=>"000110110",
89099=>"101101000",
89100=>"000000001",
89101=>"100100000",
89102=>"111011110",
89103=>"001001000",
89104=>"100111110",
89105=>"000001000",
89106=>"000110000",
89107=>"000011111",
89108=>"111111101",
89109=>"101101000",
89110=>"111111111",
89111=>"000000010",
89112=>"110101000",
89113=>"111111111",
89114=>"100101001",
89115=>"100111011",
89116=>"101101000",
89117=>"010000010",
89118=>"001011111",
89119=>"001001001",
89120=>"000000101",
89121=>"000110011",
89122=>"111011000",
89123=>"101001111",
89124=>"110110000",
89125=>"011111111",
89126=>"111111111",
89127=>"011111000",
89128=>"011000000",
89129=>"100111010",
89130=>"000111111",
89131=>"111111000",
89132=>"011010110",
89133=>"110111100",
89134=>"110110111",
89135=>"000000111",
89136=>"111000000",
89137=>"110110011",
89138=>"000001010",
89139=>"101011110",
89140=>"001000000",
89141=>"110000110",
89142=>"111110110",
89143=>"101000000",
89144=>"111000000",
89145=>"000000100",
89146=>"000011111",
89147=>"110000010",
89148=>"001000100",
89149=>"011011111",
89150=>"000000100",
89151=>"110110111",
89152=>"101101000",
89153=>"001111100",
89154=>"111111110",
89155=>"000000100",
89156=>"000000000",
89157=>"000000111",
89158=>"001011001",
89159=>"111111110",
89160=>"011011010",
89161=>"001111111",
89162=>"100000000",
89163=>"100000011",
89164=>"100001001",
89165=>"110011011",
89166=>"011000010",
89167=>"011111111",
89168=>"000010010",
89169=>"010111011",
89170=>"011001000",
89171=>"011001111",
89172=>"000101101",
89173=>"001001111",
89174=>"010011001",
89175=>"001001001",
89176=>"000110110",
89177=>"111110001",
89178=>"100001000",
89179=>"110111110",
89180=>"001001101",
89181=>"010011000",
89182=>"100101101",
89183=>"000001011",
89184=>"000000000",
89185=>"000000100",
89186=>"101101100",
89187=>"101111110",
89188=>"111111110",
89189=>"110010100",
89190=>"101101000",
89191=>"101000000",
89192=>"001011001",
89193=>"111111111",
89194=>"101111111",
89195=>"101001001",
89196=>"001000000",
89197=>"101101000",
89198=>"001000101",
89199=>"100000010",
89200=>"011001111",
89201=>"101111000",
89202=>"111001011",
89203=>"011000000",
89204=>"000000000",
89205=>"000000100",
89206=>"111111111",
89207=>"000000000",
89208=>"000111101",
89209=>"111111101",
89210=>"101100001",
89211=>"011000111",
89212=>"001000011",
89213=>"010100100",
89214=>"000010000",
89215=>"000111111",
89216=>"111101000",
89217=>"000111111",
89218=>"100100100",
89219=>"111010010",
89220=>"010000101",
89221=>"111111110",
89222=>"100111111",
89223=>"100000110",
89224=>"110000000",
89225=>"111011010",
89226=>"011101000",
89227=>"101101000",
89228=>"101101111",
89229=>"101101101",
89230=>"010111111",
89231=>"000100101",
89232=>"011010100",
89233=>"000101101",
89234=>"101101111",
89235=>"001001100",
89236=>"111110100",
89237=>"000101001",
89238=>"000010010",
89239=>"110101001",
89240=>"010101111",
89241=>"101001001",
89242=>"000000010",
89243=>"001111111",
89244=>"100011000",
89245=>"000100000",
89246=>"111111100",
89247=>"000101001",
89248=>"110100010",
89249=>"001101100",
89250=>"001010011",
89251=>"101000000",
89252=>"010010111",
89253=>"111011010",
89254=>"111001000",
89255=>"000010111",
89256=>"010100111",
89257=>"000001011",
89258=>"101000011",
89259=>"001111001",
89260=>"000100000",
89261=>"000000000",
89262=>"000000000",
89263=>"101100100",
89264=>"001001101",
89265=>"001001011",
89266=>"111000110",
89267=>"011010010",
89268=>"100111100",
89269=>"111110001",
89270=>"100000100",
89271=>"001101101",
89272=>"100000101",
89273=>"001001011",
89274=>"111101111",
89275=>"001100100",
89276=>"111110111",
89277=>"101111111",
89278=>"111001111",
89279=>"001100000",
89280=>"000000100",
89281=>"010011100",
89282=>"000000001",
89283=>"010010010",
89284=>"111111110",
89285=>"011111100",
89286=>"000100101",
89287=>"010010010",
89288=>"101100111",
89289=>"011001000",
89290=>"000101011",
89291=>"101100110",
89292=>"000001111",
89293=>"000100111",
89294=>"000000101",
89295=>"000000101",
89296=>"110010110",
89297=>"010111001",
89298=>"100010001",
89299=>"101111000",
89300=>"000000111",
89301=>"001000000",
89302=>"000101101",
89303=>"010011111",
89304=>"101001111",
89305=>"111101001",
89306=>"011001100",
89307=>"110110010",
89308=>"111111111",
89309=>"110001100",
89310=>"111111110",
89311=>"111110111",
89312=>"000001111",
89313=>"000111100",
89314=>"110011111",
89315=>"010110110",
89316=>"100001101",
89317=>"101001010",
89318=>"101000100",
89319=>"000000000",
89320=>"100101111",
89321=>"000110101",
89322=>"000001000",
89323=>"001000000",
89324=>"000000001",
89325=>"101000111",
89326=>"111111000",
89327=>"111001101",
89328=>"011011011",
89329=>"111010001",
89330=>"001000000",
89331=>"000001001",
89332=>"011110110",
89333=>"111111111",
89334=>"010001101",
89335=>"000000010",
89336=>"100101111",
89337=>"110110010",
89338=>"111111111",
89339=>"111111111",
89340=>"000010010",
89341=>"111011111",
89342=>"110111011",
89343=>"010010110",
89344=>"011001100",
89345=>"000000101",
89346=>"000000101",
89347=>"000000001",
89348=>"101111000",
89349=>"001100000",
89350=>"000000001",
89351=>"000000010",
89352=>"001001101",
89353=>"000001000",
89354=>"000110001",
89355=>"111111111",
89356=>"001000000",
89357=>"000111110",
89358=>"101001001",
89359=>"001110010",
89360=>"101111110",
89361=>"000000001",
89362=>"000101111",
89363=>"000000000",
89364=>"000000111",
89365=>"110010010",
89366=>"110101011",
89367=>"000101011",
89368=>"000101111",
89369=>"001100111",
89370=>"000101111",
89371=>"111111000",
89372=>"000100101",
89373=>"110110111",
89374=>"111111000",
89375=>"111000010",
89376=>"000000101",
89377=>"111110110",
89378=>"000000000",
89379=>"000000000",
89380=>"110000000",
89381=>"100110111",
89382=>"111101000",
89383=>"001111111",
89384=>"010110100",
89385=>"111111111",
89386=>"001011111",
89387=>"010000010",
89388=>"111111110",
89389=>"000101111",
89390=>"000111111",
89391=>"001000001",
89392=>"000000111",
89393=>"010011011",
89394=>"111011101",
89395=>"111111111",
89396=>"111111011",
89397=>"110010000",
89398=>"011011000",
89399=>"101000111",
89400=>"111000000",
89401=>"111000000",
89402=>"000000000",
89403=>"000000100",
89404=>"010111000",
89405=>"011011000",
89406=>"100000000",
89407=>"000000000",
89408=>"111111000",
89409=>"100111101",
89410=>"111101011",
89411=>"100100100",
89412=>"010000000",
89413=>"000111111",
89414=>"101001001",
89415=>"111110010",
89416=>"011111111",
89417=>"001111110",
89418=>"101000110",
89419=>"000000111",
89420=>"001000001",
89421=>"100100000",
89422=>"000111100",
89423=>"111011000",
89424=>"111000000",
89425=>"000111011",
89426=>"000000000",
89427=>"001001000",
89428=>"000000000",
89429=>"111111111",
89430=>"011001001",
89431=>"000010111",
89432=>"010001110",
89433=>"011011000",
89434=>"111000001",
89435=>"100010100",
89436=>"111000000",
89437=>"001001001",
89438=>"111111011",
89439=>"011011001",
89440=>"101000000",
89441=>"001010000",
89442=>"000000101",
89443=>"101100101",
89444=>"111111110",
89445=>"110100111",
89446=>"000110101",
89447=>"010000111",
89448=>"111101000",
89449=>"000000000",
89450=>"111011000",
89451=>"111111001",
89452=>"000010011",
89453=>"011010110",
89454=>"000000000",
89455=>"100101111",
89456=>"111111011",
89457=>"010110111",
89458=>"110110000",
89459=>"000000011",
89460=>"000010000",
89461=>"000101000",
89462=>"111111111",
89463=>"000000000",
89464=>"010010000",
89465=>"010000001",
89466=>"101111111",
89467=>"000000001",
89468=>"100110011",
89469=>"100100000",
89470=>"010111100",
89471=>"010010111",
89472=>"000001011",
89473=>"000100000",
89474=>"100010111",
89475=>"111100100",
89476=>"000100000",
89477=>"101001100",
89478=>"100011001",
89479=>"001000000",
89480=>"101111101",
89481=>"010010111",
89482=>"101100111",
89483=>"110101101",
89484=>"111000000",
89485=>"111011111",
89486=>"100001111",
89487=>"000000000",
89488=>"111011111",
89489=>"111011000",
89490=>"001000010",
89491=>"101010000",
89492=>"101101000",
89493=>"001111011",
89494=>"111111111",
89495=>"001011111",
89496=>"111110011",
89497=>"010010111",
89498=>"101000000",
89499=>"101100011",
89500=>"000000000",
89501=>"111101111",
89502=>"101111111",
89503=>"000001000",
89504=>"110111111",
89505=>"111101111",
89506=>"110111111",
89507=>"000000010",
89508=>"100001000",
89509=>"110000000",
89510=>"010110010",
89511=>"111111111",
89512=>"000110111",
89513=>"010110111",
89514=>"111001000",
89515=>"111110010",
89516=>"010000010",
89517=>"010000000",
89518=>"111111110",
89519=>"011000001",
89520=>"000000000",
89521=>"110001111",
89522=>"111111000",
89523=>"101110110",
89524=>"011011110",
89525=>"100100101",
89526=>"101000000",
89527=>"110110101",
89528=>"001001001",
89529=>"111101001",
89530=>"000110111",
89531=>"000011111",
89532=>"010010010",
89533=>"111111011",
89534=>"000001001",
89535=>"000000010",
89536=>"000000001",
89537=>"000000000",
89538=>"110100010",
89539=>"111001001",
89540=>"000000111",
89541=>"100100101",
89542=>"000001111",
89543=>"111000000",
89544=>"011101100",
89545=>"010000000",
89546=>"000000000",
89547=>"000000110",
89548=>"111111110",
89549=>"011011111",
89550=>"000000000",
89551=>"000000000",
89552=>"101000111",
89553=>"100111111",
89554=>"000011010",
89555=>"111110110",
89556=>"101001111",
89557=>"100100110",
89558=>"110110000",
89559=>"001000111",
89560=>"000010110",
89561=>"000111111",
89562=>"111111100",
89563=>"000101101",
89564=>"111110110",
89565=>"000001001",
89566=>"111110010",
89567=>"000111010",
89568=>"000000000",
89569=>"100000011",
89570=>"110110010",
89571=>"000100110",
89572=>"001000000",
89573=>"000110110",
89574=>"101101111",
89575=>"101101101",
89576=>"111111000",
89577=>"000001111",
89578=>"000011001",
89579=>"101000000",
89580=>"110111000",
89581=>"000000000",
89582=>"000010000",
89583=>"111100000",
89584=>"111111110",
89585=>"100001001",
89586=>"000001000",
89587=>"100100100",
89588=>"110101001",
89589=>"010010111",
89590=>"000000000",
89591=>"101000000",
89592=>"010110111",
89593=>"111000010",
89594=>"110010000",
89595=>"000000000",
89596=>"111101000",
89597=>"000000000",
89598=>"011101000",
89599=>"000000000",
89600=>"010000111",
89601=>"110110111",
89602=>"100100101",
89603=>"111000111",
89604=>"100000100",
89605=>"001101100",
89606=>"101100101",
89607=>"000000111",
89608=>"111010000",
89609=>"000000100",
89610=>"110110111",
89611=>"111100000",
89612=>"001000111",
89613=>"010010000",
89614=>"000000000",
89615=>"000000000",
89616=>"000000000",
89617=>"110100000",
89618=>"011000000",
89619=>"100001000",
89620=>"011111111",
89621=>"011111111",
89622=>"001111011",
89623=>"000111111",
89624=>"101100111",
89625=>"111111101",
89626=>"111011000",
89627=>"100101000",
89628=>"010011010",
89629=>"011010000",
89630=>"110111111",
89631=>"011111000",
89632=>"111101111",
89633=>"100011110",
89634=>"000111111",
89635=>"001011011",
89636=>"011100000",
89637=>"110010010",
89638=>"011011010",
89639=>"000000111",
89640=>"110000011",
89641=>"000000001",
89642=>"110101100",
89643=>"000000000",
89644=>"111111011",
89645=>"011000000",
89646=>"010001111",
89647=>"011100100",
89648=>"001111000",
89649=>"000000100",
89650=>"000000010",
89651=>"111000011",
89652=>"000010000",
89653=>"111110000",
89654=>"001010000",
89655=>"000000101",
89656=>"000000111",
89657=>"111101000",
89658=>"010111010",
89659=>"111111011",
89660=>"011011111",
89661=>"000011011",
89662=>"000000000",
89663=>"000000000",
89664=>"101001000",
89665=>"000111101",
89666=>"000111010",
89667=>"000100000",
89668=>"111111001",
89669=>"000100100",
89670=>"111101011",
89671=>"100111011",
89672=>"010010110",
89673=>"011101101",
89674=>"100100001",
89675=>"101100000",
89676=>"000000000",
89677=>"011000000",
89678=>"110100001",
89679=>"010110011",
89680=>"000010000",
89681=>"111111111",
89682=>"011111000",
89683=>"001001001",
89684=>"011010000",
89685=>"011011110",
89686=>"001100011",
89687=>"001010011",
89688=>"111111111",
89689=>"010011111",
89690=>"101001000",
89691=>"000000000",
89692=>"000000000",
89693=>"011001010",
89694=>"111000101",
89695=>"001001101",
89696=>"111101000",
89697=>"001000011",
89698=>"111000011",
89699=>"100110100",
89700=>"111000000",
89701=>"100011111",
89702=>"100011001",
89703=>"011000101",
89704=>"101011111",
89705=>"101111111",
89706=>"001000111",
89707=>"111101000",
89708=>"111000001",
89709=>"111101000",
89710=>"100110110",
89711=>"000101101",
89712=>"101000100",
89713=>"100100101",
89714=>"111011000",
89715=>"101000000",
89716=>"101101000",
89717=>"111000010",
89718=>"111100000",
89719=>"010010010",
89720=>"001111010",
89721=>"000011111",
89722=>"111101110",
89723=>"010000111",
89724=>"100100010",
89725=>"011110110",
89726=>"100000111",
89727=>"100110000",
89728=>"111000000",
89729=>"100100110",
89730=>"000000110",
89731=>"001000111",
89732=>"011101001",
89733=>"100000010",
89734=>"000011001",
89735=>"010010000",
89736=>"100000100",
89737=>"000010000",
89738=>"111111000",
89739=>"111100111",
89740=>"101101100",
89741=>"111101101",
89742=>"000101111",
89743=>"111000000",
89744=>"010000000",
89745=>"100100000",
89746=>"100000010",
89747=>"111111000",
89748=>"011010000",
89749=>"100100000",
89750=>"111110101",
89751=>"011000000",
89752=>"111101000",
89753=>"000011010",
89754=>"110111111",
89755=>"000000100",
89756=>"000000000",
89757=>"111101111",
89758=>"000000000",
89759=>"000100000",
89760=>"000011101",
89761=>"001111111",
89762=>"011000000",
89763=>"000111111",
89764=>"101011110",
89765=>"100001000",
89766=>"010001011",
89767=>"000000000",
89768=>"010000110",
89769=>"111010000",
89770=>"110101001",
89771=>"010111101",
89772=>"000110110",
89773=>"100000100",
89774=>"010110101",
89775=>"000000001",
89776=>"010000000",
89777=>"111111001",
89778=>"111100000",
89779=>"001000001",
89780=>"000101000",
89781=>"010111011",
89782=>"111011100",
89783=>"000111111",
89784=>"001011011",
89785=>"100010011",
89786=>"111011111",
89787=>"100101110",
89788=>"111000010",
89789=>"111100111",
89790=>"110100010",
89791=>"000000000",
89792=>"011011000",
89793=>"110101000",
89794=>"100000000",
89795=>"111000100",
89796=>"101111101",
89797=>"001100111",
89798=>"111101101",
89799=>"000011110",
89800=>"010000101",
89801=>"000011111",
89802=>"000101111",
89803=>"101101111",
89804=>"010000000",
89805=>"110010000",
89806=>"110111111",
89807=>"111000101",
89808=>"111011001",
89809=>"010100101",
89810=>"111000011",
89811=>"000101000",
89812=>"101101101",
89813=>"011110000",
89814=>"111111000",
89815=>"111111000",
89816=>"000011000",
89817=>"010000000",
89818=>"000111110",
89819=>"101100100",
89820=>"110111110",
89821=>"110010010",
89822=>"111100000",
89823=>"000101100",
89824=>"000111001",
89825=>"111101111",
89826=>"011010111",
89827=>"011001100",
89828=>"100000000",
89829=>"111101101",
89830=>"110000000",
89831=>"000010101",
89832=>"111100000",
89833=>"000000000",
89834=>"001111110",
89835=>"011111111",
89836=>"000000111",
89837=>"011000000",
89838=>"000000010",
89839=>"110111010",
89840=>"111111010",
89841=>"000110001",
89842=>"100101111",
89843=>"010110110",
89844=>"011101110",
89845=>"001111101",
89846=>"100000000",
89847=>"000000000",
89848=>"000100011",
89849=>"000001010",
89850=>"000011111",
89851=>"101111010",
89852=>"101101000",
89853=>"010110010",
89854=>"100000000",
89855=>"111100111",
89856=>"011001011",
89857=>"111110011",
89858=>"000100100",
89859=>"000000011",
89860=>"100011001",
89861=>"010110100",
89862=>"111011011",
89863=>"111001011",
89864=>"100110100",
89865=>"000000000",
89866=>"000111111",
89867=>"011101110",
89868=>"000000000",
89869=>"000000000",
89870=>"100100111",
89871=>"110010010",
89872=>"100000001",
89873=>"101111100",
89874=>"010000000",
89875=>"100110011",
89876=>"101111000",
89877=>"101111101",
89878=>"000101111",
89879=>"100000111",
89880=>"000000000",
89881=>"011111011",
89882=>"000011010",
89883=>"111100100",
89884=>"101100011",
89885=>"111010001",
89886=>"111111010",
89887=>"000111110",
89888=>"000100101",
89889=>"110110111",
89890=>"000001000",
89891=>"000000000",
89892=>"001000000",
89893=>"100000011",
89894=>"111011011",
89895=>"000100000",
89896=>"100111101",
89897=>"001010111",
89898=>"000000011",
89899=>"001000010",
89900=>"110001011",
89901=>"011110111",
89902=>"110110100",
89903=>"000101100",
89904=>"000001011",
89905=>"011010110",
89906=>"111100000",
89907=>"000111011",
89908=>"101111111",
89909=>"000011011",
89910=>"111011111",
89911=>"000001000",
89912=>"010010000",
89913=>"111100110",
89914=>"011000000",
89915=>"000011000",
89916=>"111001000",
89917=>"111111110",
89918=>"101100100",
89919=>"110111111",
89920=>"111111011",
89921=>"000100110",
89922=>"110000001",
89923=>"001111011",
89924=>"000000001",
89925=>"011000000",
89926=>"001011011",
89927=>"011011111",
89928=>"111110100",
89929=>"100000011",
89930=>"000100100",
89931=>"000100000",
89932=>"100100100",
89933=>"111111101",
89934=>"001111111",
89935=>"000011111",
89936=>"000000000",
89937=>"111100100",
89938=>"000101011",
89939=>"000001011",
89940=>"100100100",
89941=>"111110010",
89942=>"000100110",
89943=>"101000000",
89944=>"000000000",
89945=>"000000001",
89946=>"000000011",
89947=>"110110111",
89948=>"000000000",
89949=>"011000010",
89950=>"000011111",
89951=>"110110001",
89952=>"000011011",
89953=>"000000001",
89954=>"000000100",
89955=>"001000001",
89956=>"110110011",
89957=>"110110111",
89958=>"100100010",
89959=>"110100000",
89960=>"011111011",
89961=>"011011111",
89962=>"011010000",
89963=>"100101111",
89964=>"100100110",
89965=>"001011101",
89966=>"110110100",
89967=>"000000000",
89968=>"000000000",
89969=>"111000000",
89970=>"011111111",
89971=>"111100100",
89972=>"000000000",
89973=>"100100100",
89974=>"001011000",
89975=>"000011011",
89976=>"000010001",
89977=>"100000011",
89978=>"011100110",
89979=>"000000001",
89980=>"001100000",
89981=>"000000000",
89982=>"111100111",
89983=>"111100100",
89984=>"100000011",
89985=>"011011100",
89986=>"000001000",
89987=>"000001010",
89988=>"100110111",
89989=>"100111111",
89990=>"010110110",
89991=>"010000000",
89992=>"110111101",
89993=>"000001000",
89994=>"110000010",
89995=>"011000000",
89996=>"000000000",
89997=>"100111000",
89998=>"000001011",
89999=>"000000000",
90000=>"000000000",
90001=>"000100111",
90002=>"001100100",
90003=>"111100101",
90004=>"110111100",
90005=>"111101000",
90006=>"000011110",
90007=>"110011011",
90008=>"000111011",
90009=>"111100001",
90010=>"100100101",
90011=>"000010011",
90012=>"000000000",
90013=>"110111011",
90014=>"000001011",
90015=>"100100111",
90016=>"000100000",
90017=>"100110000",
90018=>"010011001",
90019=>"100011011",
90020=>"101100100",
90021=>"100010011",
90022=>"110010011",
90023=>"010011011",
90024=>"011100000",
90025=>"001011111",
90026=>"000110111",
90027=>"100110111",
90028=>"010011100",
90029=>"010100001",
90030=>"100100100",
90031=>"011011011",
90032=>"010100100",
90033=>"001100100",
90034=>"100010111",
90035=>"001100000",
90036=>"000001001",
90037=>"011011000",
90038=>"000001011",
90039=>"000000000",
90040=>"010010000",
90041=>"010010111",
90042=>"001001111",
90043=>"000001011",
90044=>"111001000",
90045=>"011111110",
90046=>"000001000",
90047=>"011001000",
90048=>"011111111",
90049=>"000011011",
90050=>"000011011",
90051=>"100100110",
90052=>"010100000",
90053=>"011010110",
90054=>"000000010",
90055=>"111111000",
90056=>"100000011",
90057=>"110001010",
90058=>"000011011",
90059=>"111111111",
90060=>"100011010",
90061=>"100111110",
90062=>"011011000",
90063=>"100110110",
90064=>"000100110",
90065=>"001111111",
90066=>"001000100",
90067=>"000111011",
90068=>"000100100",
90069=>"011010000",
90070=>"011100110",
90071=>"110010111",
90072=>"011000101",
90073=>"010000000",
90074=>"100111111",
90075=>"110100000",
90076=>"101111111",
90077=>"011011110",
90078=>"000011011",
90079=>"100110011",
90080=>"000000000",
90081=>"111110000",
90082=>"101111110",
90083=>"000000101",
90084=>"111100100",
90085=>"000111101",
90086=>"111110000",
90087=>"011111000",
90088=>"111100100",
90089=>"011100100",
90090=>"111001101",
90091=>"000011011",
90092=>"000000000",
90093=>"011100100",
90094=>"011000000",
90095=>"100100000",
90096=>"111100100",
90097=>"101001100",
90098=>"011000000",
90099=>"101110111",
90100=>"010011010",
90101=>"010000100",
90102=>"001000001",
90103=>"110110100",
90104=>"000001111",
90105=>"110010011",
90106=>"001001001",
90107=>"011011111",
90108=>"111000111",
90109=>"110100100",
90110=>"000011011",
90111=>"100111011",
90112=>"001000000",
90113=>"000001101",
90114=>"101000101",
90115=>"011000011",
90116=>"000011111",
90117=>"111101101",
90118=>"111000101",
90119=>"111011101",
90120=>"011000000",
90121=>"100000100",
90122=>"100111001",
90123=>"110010010",
90124=>"011001011",
90125=>"111111000",
90126=>"100111100",
90127=>"011010000",
90128=>"000100111",
90129=>"101101001",
90130=>"000001110",
90131=>"101000001",
90132=>"111111111",
90133=>"000111000",
90134=>"110000111",
90135=>"111111110",
90136=>"000000100",
90137=>"001000100",
90138=>"110111011",
90139=>"000111111",
90140=>"000000101",
90141=>"000000101",
90142=>"111100111",
90143=>"000000000",
90144=>"001000011",
90145=>"101111010",
90146=>"100101001",
90147=>"101000101",
90148=>"001111111",
90149=>"100001000",
90150=>"010000000",
90151=>"000111101",
90152=>"100010100",
90153=>"001001001",
90154=>"010111011",
90155=>"001000111",
90156=>"000111110",
90157=>"111110011",
90158=>"111001100",
90159=>"001000000",
90160=>"000101000",
90161=>"111010000",
90162=>"000000000",
90163=>"100000100",
90164=>"111011000",
90165=>"101111001",
90166=>"101101100",
90167=>"111111000",
90168=>"111010010",
90169=>"101111111",
90170=>"000010010",
90171=>"000111000",
90172=>"011111011",
90173=>"000000001",
90174=>"000000101",
90175=>"011111011",
90176=>"101101101",
90177=>"000000101",
90178=>"000000000",
90179=>"011011001",
90180=>"111111010",
90181=>"001000000",
90182=>"011010000",
90183=>"000010011",
90184=>"111111111",
90185=>"010111010",
90186=>"010001001",
90187=>"010001000",
90188=>"111000000",
90189=>"111111011",
90190=>"001000111",
90191=>"000111111",
90192=>"000000000",
90193=>"111111111",
90194=>"111111000",
90195=>"011001000",
90196=>"101101000",
90197=>"001011110",
90198=>"001100011",
90199=>"111101101",
90200=>"000000011",
90201=>"000011010",
90202=>"100011010",
90203=>"000100100",
90204=>"000101101",
90205=>"000100110",
90206=>"011000010",
90207=>"110110101",
90208=>"000000100",
90209=>"001010000",
90210=>"111001111",
90211=>"000111010",
90212=>"000001010",
90213=>"011010000",
90214=>"010110111",
90215=>"111111010",
90216=>"010011001",
90217=>"010010110",
90218=>"110000110",
90219=>"111111111",
90220=>"000000111",
90221=>"001111110",
90222=>"001001000",
90223=>"010101110",
90224=>"001110000",
90225=>"000010110",
90226=>"101101001",
90227=>"000000000",
90228=>"111100000",
90229=>"010000000",
90230=>"000011111",
90231=>"111000100",
90232=>"000000111",
90233=>"000111011",
90234=>"100111000",
90235=>"010111111",
90236=>"001001101",
90237=>"010100000",
90238=>"000111000",
90239=>"000111000",
90240=>"110111001",
90241=>"010000010",
90242=>"000111101",
90243=>"000000100",
90244=>"111111111",
90245=>"111110001",
90246=>"001000011",
90247=>"000001100",
90248=>"100011010",
90249=>"001000000",
90250=>"011111010",
90251=>"000010111",
90252=>"100001101",
90253=>"001101101",
90254=>"101010111",
90255=>"000000000",
90256=>"111111000",
90257=>"001111000",
90258=>"111110000",
90259=>"100000111",
90260=>"101000011",
90261=>"101000101",
90262=>"000010111",
90263=>"010000100",
90264=>"000011000",
90265=>"100000001",
90266=>"111111000",
90267=>"000000111",
90268=>"111111110",
90269=>"100000110",
90270=>"110010011",
90271=>"101000110",
90272=>"100010001",
90273=>"111101101",
90274=>"000000010",
90275=>"010111010",
90276=>"010110011",
90277=>"101000000",
90278=>"010001100",
90279=>"101111101",
90280=>"100100100",
90281=>"110111001",
90282=>"111000001",
90283=>"111101101",
90284=>"001101011",
90285=>"110000000",
90286=>"000000000",
90287=>"111000010",
90288=>"100000101",
90289=>"001000111",
90290=>"000010000",
90291=>"001001011",
90292=>"111111011",
90293=>"000001001",
90294=>"000000000",
90295=>"101110010",
90296=>"100111110",
90297=>"000000110",
90298=>"111000000",
90299=>"011000111",
90300=>"000000000",
90301=>"111111100",
90302=>"110011000",
90303=>"000000000",
90304=>"111000000",
90305=>"000001001",
90306=>"111110001",
90307=>"111010000",
90308=>"001111000",
90309=>"111001101",
90310=>"011000010",
90311=>"001001101",
90312=>"110110000",
90313=>"010100000",
90314=>"000000001",
90315=>"001000000",
90316=>"000001000",
90317=>"000100101",
90318=>"000000101",
90319=>"000001111",
90320=>"000110000",
90321=>"111110100",
90322=>"100110111",
90323=>"010011000",
90324=>"101001111",
90325=>"100000011",
90326=>"010011111",
90327=>"010010111",
90328=>"001011001",
90329=>"000000010",
90330=>"000000000",
90331=>"000010000",
90332=>"010101011",
90333=>"110111110",
90334=>"000000010",
90335=>"101110010",
90336=>"111000000",
90337=>"111100001",
90338=>"100110001",
90339=>"001111111",
90340=>"000000000",
90341=>"111111001",
90342=>"001011111",
90343=>"001001000",
90344=>"000010111",
90345=>"101011111",
90346=>"001111100",
90347=>"000000001",
90348=>"000000000",
90349=>"000010010",
90350=>"000000000",
90351=>"010101111",
90352=>"111110000",
90353=>"111110000",
90354=>"111101111",
90355=>"111110110",
90356=>"000111011",
90357=>"000000000",
90358=>"000000100",
90359=>"100111001",
90360=>"011001011",
90361=>"011011000",
90362=>"000011000",
90363=>"000101101",
90364=>"010000101",
90365=>"000001000",
90366=>"101111110",
90367=>"011010001",
90368=>"011101111",
90369=>"001000000",
90370=>"000000000",
90371=>"000100110",
90372=>"111011001",
90373=>"000001111",
90374=>"101100000",
90375=>"111111010",
90376=>"001001111",
90377=>"000001000",
90378=>"011100100",
90379=>"000000000",
90380=>"000000111",
90381=>"000000100",
90382=>"110111111",
90383=>"101111101",
90384=>"100111111",
90385=>"000000111",
90386=>"111111000",
90387=>"000000000",
90388=>"110110000",
90389=>"100000010",
90390=>"101111111",
90391=>"111111011",
90392=>"000001001",
90393=>"000000111",
90394=>"000000111",
90395=>"000000001",
90396=>"101111101",
90397=>"000011111",
90398=>"111111111",
90399=>"000110110",
90400=>"000000010",
90401=>"000000000",
90402=>"111011100",
90403=>"000000000",
90404=>"111001001",
90405=>"101001001",
90406=>"000000001",
90407=>"111011100",
90408=>"111010000",
90409=>"000001010",
90410=>"111001111",
90411=>"111111111",
90412=>"001101111",
90413=>"011000000",
90414=>"111111101",
90415=>"110111111",
90416=>"000000000",
90417=>"111111011",
90418=>"000000001",
90419=>"101111100",
90420=>"000111110",
90421=>"111110111",
90422=>"000000010",
90423=>"011011111",
90424=>"111111001",
90425=>"010001000",
90426=>"000000111",
90427=>"100000010",
90428=>"001001001",
90429=>"111111111",
90430=>"000000111",
90431=>"111001001",
90432=>"010001000",
90433=>"010000000",
90434=>"000111111",
90435=>"111110110",
90436=>"110000000",
90437=>"101111100",
90438=>"111110110",
90439=>"010100100",
90440=>"010101101",
90441=>"111101101",
90442=>"111101111",
90443=>"000101111",
90444=>"000001000",
90445=>"111111010",
90446=>"100110110",
90447=>"100000110",
90448=>"000100111",
90449=>"111111000",
90450=>"000000111",
90451=>"001000000",
90452=>"111000000",
90453=>"000100100",
90454=>"001011110",
90455=>"000000010",
90456=>"011000111",
90457=>"001001001",
90458=>"110000011",
90459=>"000100111",
90460=>"001001111",
90461=>"101000001",
90462=>"111111000",
90463=>"111101110",
90464=>"111111111",
90465=>"000100110",
90466=>"000000000",
90467=>"111010000",
90468=>"100000100",
90469=>"000000000",
90470=>"000101001",
90471=>"111011010",
90472=>"010000000",
90473=>"100001101",
90474=>"111000000",
90475=>"000000000",
90476=>"000111011",
90477=>"000000000",
90478=>"000000000",
90479=>"000000101",
90480=>"100000110",
90481=>"000000111",
90482=>"010000000",
90483=>"000101111",
90484=>"100101101",
90485=>"000101101",
90486=>"000000000",
90487=>"110101100",
90488=>"111100000",
90489=>"000001111",
90490=>"011000001",
90491=>"111110000",
90492=>"110110100",
90493=>"100000001",
90494=>"111111010",
90495=>"000000111",
90496=>"000001000",
90497=>"111111111",
90498=>"110111111",
90499=>"001011100",
90500=>"100110110",
90501=>"101100011",
90502=>"000000100",
90503=>"000000000",
90504=>"011001011",
90505=>"110111111",
90506=>"111111011",
90507=>"000000100",
90508=>"000000000",
90509=>"001101110",
90510=>"011110000",
90511=>"000000000",
90512=>"011011001",
90513=>"111000100",
90514=>"000001000",
90515=>"111110010",
90516=>"000111111",
90517=>"000000100",
90518=>"111111111",
90519=>"001001011",
90520=>"000001110",
90521=>"111111100",
90522=>"011111000",
90523=>"000110000",
90524=>"100000000",
90525=>"000000001",
90526=>"101110110",
90527=>"101111111",
90528=>"001000001",
90529=>"101110111",
90530=>"111001111",
90531=>"000100000",
90532=>"101111011",
90533=>"001001101",
90534=>"100100111",
90535=>"111111111",
90536=>"000111111",
90537=>"011110000",
90538=>"000000000",
90539=>"001000000",
90540=>"011010001",
90541=>"000000001",
90542=>"011010110",
90543=>"011010000",
90544=>"111000000",
90545=>"101000101",
90546=>"000100110",
90547=>"000000100",
90548=>"011111101",
90549=>"111111111",
90550=>"010000000",
90551=>"000000000",
90552=>"110000101",
90553=>"001010010",
90554=>"001000101",
90555=>"011010100",
90556=>"000010000",
90557=>"000101000",
90558=>"101100100",
90559=>"000101111",
90560=>"111010010",
90561=>"011001111",
90562=>"000111010",
90563=>"001001001",
90564=>"000111000",
90565=>"000000000",
90566=>"011101111",
90567=>"110111111",
90568=>"111110000",
90569=>"010001001",
90570=>"110000000",
90571=>"000000000",
90572=>"011111010",
90573=>"111011011",
90574=>"000000000",
90575=>"000001011",
90576=>"000111111",
90577=>"110111111",
90578=>"000000000",
90579=>"101111111",
90580=>"000000000",
90581=>"001001001",
90582=>"101000001",
90583=>"000111011",
90584=>"111111110",
90585=>"011111010",
90586=>"100000110",
90587=>"000001000",
90588=>"010111101",
90589=>"000000100",
90590=>"000010110",
90591=>"001101111",
90592=>"000000000",
90593=>"000000000",
90594=>"111000000",
90595=>"100111111",
90596=>"001001011",
90597=>"100001100",
90598=>"000000000",
90599=>"111100100",
90600=>"000000111",
90601=>"000000010",
90602=>"110001001",
90603=>"000000100",
90604=>"000000000",
90605=>"000000000",
90606=>"000000001",
90607=>"001000000",
90608=>"000100111",
90609=>"000000100",
90610=>"001101100",
90611=>"111111111",
90612=>"100101001",
90613=>"110111101",
90614=>"000000100",
90615=>"000001011",
90616=>"111110010",
90617=>"000110100",
90618=>"111111111",
90619=>"000010010",
90620=>"111111010",
90621=>"000000000",
90622=>"110110110",
90623=>"111111111",
90624=>"110010111",
90625=>"011110110",
90626=>"001001111",
90627=>"000010111",
90628=>"010011110",
90629=>"000011011",
90630=>"100110100",
90631=>"100110001",
90632=>"010000001",
90633=>"011000011",
90634=>"110101001",
90635=>"111111011",
90636=>"011001011",
90637=>"001001001",
90638=>"100010000",
90639=>"101100000",
90640=>"100100001",
90641=>"000100100",
90642=>"001001000",
90643=>"001100100",
90644=>"110110100",
90645=>"011011011",
90646=>"110000110",
90647=>"001100101",
90648=>"100000001",
90649=>"101001001",
90650=>"001000110",
90651=>"000100110",
90652=>"111101110",
90653=>"011011011",
90654=>"100000011",
90655=>"001001000",
90656=>"001001101",
90657=>"100101101",
90658=>"111001011",
90659=>"001011001",
90660=>"010000000",
90661=>"111101100",
90662=>"111110010",
90663=>"000100001",
90664=>"010111111",
90665=>"100110001",
90666=>"110100100",
90667=>"000001111",
90668=>"111111110",
90669=>"110110101",
90670=>"010000110",
90671=>"001001000",
90672=>"100100000",
90673=>"010011110",
90674=>"000000000",
90675=>"101101000",
90676=>"000000001",
90677=>"110111110",
90678=>"011011000",
90679=>"110011000",
90680=>"000111011",
90681=>"110000011",
90682=>"001001110",
90683=>"000100100",
90684=>"011010010",
90685=>"111011111",
90686=>"001001001",
90687=>"000110000",
90688=>"101101011",
90689=>"001010111",
90690=>"011001000",
90691=>"001011101",
90692=>"010011010",
90693=>"000000100",
90694=>"000000100",
90695=>"011111011",
90696=>"111111011",
90697=>"110100110",
90698=>"100100000",
90699=>"011000001",
90700=>"001000100",
90701=>"111011001",
90702=>"111000101",
90703=>"101111100",
90704=>"010000100",
90705=>"000011011",
90706=>"001100101",
90707=>"101111000",
90708=>"100100010",
90709=>"000000000",
90710=>"100000010",
90711=>"101001111",
90712=>"110110111",
90713=>"110111001",
90714=>"100101111",
90715=>"011001000",
90716=>"101101101",
90717=>"010011100",
90718=>"001111111",
90719=>"010000011",
90720=>"011011011",
90721=>"010001000",
90722=>"001001001",
90723=>"000010000",
90724=>"000001010",
90725=>"011011001",
90726=>"111110101",
90727=>"111011011",
90728=>"100101011",
90729=>"101101111",
90730=>"100000100",
90731=>"110011001",
90732=>"011001110",
90733=>"110100100",
90734=>"101000011",
90735=>"001111100",
90736=>"010000001",
90737=>"100000000",
90738=>"000001001",
90739=>"000011000",
90740=>"001001001",
90741=>"000001010",
90742=>"001001010",
90743=>"000011000",
90744=>"110111110",
90745=>"000000110",
90746=>"100100101",
90747=>"000010000",
90748=>"101011011",
90749=>"001001000",
90750=>"000100011",
90751=>"011011001",
90752=>"001101100",
90753=>"010010001",
90754=>"011001101",
90755=>"010011111",
90756=>"101101101",
90757=>"011011111",
90758=>"100111110",
90759=>"100111001",
90760=>"000000001",
90761=>"011000000",
90762=>"001100000",
90763=>"000000100",
90764=>"001110001",
90765=>"010011111",
90766=>"000110100",
90767=>"111001000",
90768=>"110011011",
90769=>"100011110",
90770=>"001100000",
90771=>"111011001",
90772=>"111110100",
90773=>"001000100",
90774=>"110110100",
90775=>"000010000",
90776=>"111111011",
90777=>"011100110",
90778=>"011011001",
90779=>"001011011",
90780=>"111111001",
90781=>"000000001",
90782=>"100100111",
90783=>"011101111",
90784=>"111100001",
90785=>"100100001",
90786=>"000010110",
90787=>"001011010",
90788=>"100100101",
90789=>"100000000",
90790=>"100001001",
90791=>"111110111",
90792=>"011100100",
90793=>"100100000",
90794=>"001001111",
90795=>"001001001",
90796=>"001001100",
90797=>"000001001",
90798=>"111111000",
90799=>"101011001",
90800=>"001000000",
90801=>"110100011",
90802=>"101011110",
90803=>"101001001",
90804=>"010110110",
90805=>"011110110",
90806=>"101001011",
90807=>"100111110",
90808=>"000000000",
90809=>"000000000",
90810=>"000011011",
90811=>"110111100",
90812=>"101001111",
90813=>"001001011",
90814=>"001000000",
90815=>"010010000",
90816=>"011001100",
90817=>"000100001",
90818=>"100011100",
90819=>"011010000",
90820=>"100100100",
90821=>"010001000",
90822=>"001101100",
90823=>"011011110",
90824=>"100110000",
90825=>"011000000",
90826=>"011111011",
90827=>"111110011",
90828=>"110111001",
90829=>"110010000",
90830=>"000001011",
90831=>"001111001",
90832=>"101111001",
90833=>"010111011",
90834=>"111011001",
90835=>"001000000",
90836=>"001001001",
90837=>"110110110",
90838=>"100001001",
90839=>"100100100",
90840=>"100110100",
90841=>"100001000",
90842=>"011000000",
90843=>"100101100",
90844=>"000110000",
90845=>"000010000",
90846=>"110010000",
90847=>"000001111",
90848=>"110001000",
90849=>"100001010",
90850=>"100100110",
90851=>"001000001",
90852=>"011000100",
90853=>"011111011",
90854=>"111011011",
90855=>"000111110",
90856=>"111011111",
90857=>"000110110",
90858=>"000100110",
90859=>"111100110",
90860=>"011011001",
90861=>"101101110",
90862=>"000001110",
90863=>"110000100",
90864=>"110000100",
90865=>"111111111",
90866=>"100000100",
90867=>"110110000",
90868=>"011010001",
90869=>"100111110",
90870=>"000000100",
90871=>"110010110",
90872=>"100100001",
90873=>"100011000",
90874=>"011011111",
90875=>"100010100",
90876=>"011110100",
90877=>"001010011",
90878=>"110011111",
90879=>"000001110",
90880=>"000111000",
90881=>"010000011",
90882=>"101100001",
90883=>"111111010",
90884=>"100110100",
90885=>"100000111",
90886=>"111000100",
90887=>"010000000",
90888=>"110010000",
90889=>"010000001",
90890=>"111101100",
90891=>"000111000",
90892=>"101000101",
90893=>"111111011",
90894=>"000000000",
90895=>"000000000",
90896=>"011111111",
90897=>"111110110",
90898=>"101100111",
90899=>"001000000",
90900=>"100000111",
90901=>"111101100",
90902=>"111111100",
90903=>"110110111",
90904=>"000001111",
90905=>"000001100",
90906=>"000000000",
90907=>"110111001",
90908=>"111111011",
90909=>"010000010",
90910=>"101011000",
90911=>"111111111",
90912=>"111111000",
90913=>"001000000",
90914=>"000000110",
90915=>"000000000",
90916=>"000000000",
90917=>"110100000",
90918=>"000000000",
90919=>"111111111",
90920=>"111000111",
90921=>"000010010",
90922=>"111111111",
90923=>"000111110",
90924=>"111110111",
90925=>"000000000",
90926=>"000111111",
90927=>"000100000",
90928=>"000110000",
90929=>"000111110",
90930=>"000001111",
90931=>"111110010",
90932=>"101100111",
90933=>"010111010",
90934=>"011001110",
90935=>"001001011",
90936=>"111000000",
90937=>"000000000",
90938=>"100110111",
90939=>"000000011",
90940=>"100110110",
90941=>"111111111",
90942=>"000000000",
90943=>"111111101",
90944=>"011000001",
90945=>"010110000",
90946=>"000000000",
90947=>"110101100",
90948=>"000010000",
90949=>"001001100",
90950=>"101001000",
90951=>"001000111",
90952=>"000000000",
90953=>"110111010",
90954=>"001000000",
90955=>"111110111",
90956=>"000000000",
90957=>"111001110",
90958=>"000001001",
90959=>"011010111",
90960=>"111111111",
90961=>"110110111",
90962=>"000000000",
90963=>"001001000",
90964=>"111110110",
90965=>"100011011",
90966=>"001001000",
90967=>"111111111",
90968=>"000000111",
90969=>"000001110",
90970=>"001001000",
90971=>"111111111",
90972=>"000000000",
90973=>"001100010",
90974=>"001001000",
90975=>"111111111",
90976=>"111110110",
90977=>"111010010",
90978=>"101000000",
90979=>"000111100",
90980=>"100000110",
90981=>"000111111",
90982=>"111111110",
90983=>"000000000",
90984=>"111111000",
90985=>"000000000",
90986=>"100000111",
90987=>"010000000",
90988=>"000000000",
90989=>"110110000",
90990=>"111111000",
90991=>"110000000",
90992=>"111111011",
90993=>"000000010",
90994=>"000110010",
90995=>"000001101",
90996=>"000001001",
90997=>"001001001",
90998=>"011111111",
90999=>"011111111",
91000=>"111111111",
91001=>"110010010",
91002=>"000111001",
91003=>"000000100",
91004=>"111110000",
91005=>"110110000",
91006=>"111111001",
91007=>"111111110",
91008=>"001101000",
91009=>"111111100",
91010=>"000110000",
91011=>"000000000",
91012=>"111101000",
91013=>"000011111",
91014=>"011011001",
91015=>"010010110",
91016=>"011111011",
91017=>"000000001",
91018=>"010011111",
91019=>"001000000",
91020=>"000001000",
91021=>"111111111",
91022=>"000111100",
91023=>"101001001",
91024=>"000001011",
91025=>"111000000",
91026=>"111111000",
91027=>"111111000",
91028=>"011111111",
91029=>"111111011",
91030=>"011111001",
91031=>"010011010",
91032=>"111111111",
91033=>"101000000",
91034=>"111111001",
91035=>"110111111",
91036=>"010010000",
91037=>"010111000",
91038=>"011111111",
91039=>"000111111",
91040=>"000000000",
91041=>"010110010",
91042=>"111111000",
91043=>"000000001",
91044=>"100010111",
91045=>"100010010",
91046=>"000000000",
91047=>"000100100",
91048=>"010000010",
91049=>"000100101",
91050=>"000000000",
91051=>"110110110",
91052=>"101101111",
91053=>"101000000",
91054=>"111111110",
91055=>"000000001",
91056=>"000000101",
91057=>"000000111",
91058=>"000110100",
91059=>"100000001",
91060=>"000010011",
91061=>"011001111",
91062=>"000000110",
91063=>"000001101",
91064=>"000011111",
91065=>"110110010",
91066=>"000010111",
91067=>"110111010",
91068=>"101010011",
91069=>"111111110",
91070=>"100110111",
91071=>"000000111",
91072=>"111000101",
91073=>"010011011",
91074=>"011010000",
91075=>"111010111",
91076=>"000000000",
91077=>"110000000",
91078=>"010000000",
91079=>"110100000",
91080=>"000101111",
91081=>"000111010",
91082=>"000101000",
91083=>"111111001",
91084=>"011011011",
91085=>"111001000",
91086=>"000000000",
91087=>"010110000",
91088=>"111111000",
91089=>"110110010",
91090=>"010001000",
91091=>"000000000",
91092=>"010001100",
91093=>"000000000",
91094=>"101101101",
91095=>"111111111",
91096=>"000000001",
91097=>"110010101",
91098=>"000010001",
91099=>"111111101",
91100=>"001111110",
91101=>"000000100",
91102=>"000000000",
91103=>"100001000",
91104=>"000000000",
91105=>"000000001",
91106=>"000000000",
91107=>"011111011",
91108=>"000011101",
91109=>"000000000",
91110=>"001111101",
91111=>"011011010",
91112=>"110000000",
91113=>"111110100",
91114=>"111001001",
91115=>"000111111",
91116=>"000111111",
91117=>"111101000",
91118=>"110110000",
91119=>"000000110",
91120=>"000000001",
91121=>"011001000",
91122=>"000000011",
91123=>"000110000",
91124=>"000111011",
91125=>"111111001",
91126=>"111000010",
91127=>"000000000",
91128=>"110111001",
91129=>"000000000",
91130=>"000110000",
91131=>"000000010",
91132=>"111111000",
91133=>"000000000",
91134=>"001100011",
91135=>"001111111",
91136=>"100001001",
91137=>"100100111",
91138=>"100000100",
91139=>"010001100",
91140=>"111111011",
91141=>"110101110",
91142=>"111010011",
91143=>"000000000",
91144=>"010011011",
91145=>"100100110",
91146=>"000100000",
91147=>"100100100",
91148=>"110000110",
91149=>"110100000",
91150=>"100110111",
91151=>"000001000",
91152=>"111000001",
91153=>"000000111",
91154=>"010110111",
91155=>"100110000",
91156=>"110000110",
91157=>"000100111",
91158=>"101000111",
91159=>"111100101",
91160=>"100000110",
91161=>"100100111",
91162=>"110100100",
91163=>"011001000",
91164=>"100001111",
91165=>"010010000",
91166=>"101100100",
91167=>"011011011",
91168=>"111001000",
91169=>"111100011",
91170=>"000000001",
91171=>"000000000",
91172=>"001001001",
91173=>"000000000",
91174=>"000011011",
91175=>"011010000",
91176=>"110100000",
91177=>"000000011",
91178=>"100100100",
91179=>"111110110",
91180=>"111010111",
91181=>"100011011",
91182=>"001100110",
91183=>"101111010",
91184=>"001011010",
91185=>"100110111",
91186=>"001011011",
91187=>"011111110",
91188=>"110100110",
91189=>"000010011",
91190=>"000110111",
91191=>"011011011",
91192=>"011111000",
91193=>"100100100",
91194=>"010110110",
91195=>"000000100",
91196=>"000010010",
91197=>"011011010",
91198=>"010000100",
91199=>"101001000",
91200=>"110100100",
91201=>"000000000",
91202=>"000001011",
91203=>"110110111",
91204=>"011111000",
91205=>"000000000",
91206=>"101101111",
91207=>"101111000",
91208=>"000011011",
91209=>"000000110",
91210=>"010000000",
91211=>"100100110",
91212=>"001000100",
91213=>"111011111",
91214=>"011000000",
91215=>"001011011",
91216=>"000000001",
91217=>"100000000",
91218=>"100110111",
91219=>"101000000",
91220=>"100100000",
91221=>"000000011",
91222=>"110001001",
91223=>"000100100",
91224=>"110100000",
91225=>"001111111",
91226=>"001000000",
91227=>"111110110",
91228=>"000011011",
91229=>"000101100",
91230=>"000001011",
91231=>"100000001",
91232=>"001011011",
91233=>"011011000",
91234=>"100100100",
91235=>"111111111",
91236=>"010010010",
91237=>"111111100",
91238=>"100100110",
91239=>"011000000",
91240=>"011011000",
91241=>"001010100",
91242=>"000000111",
91243=>"110110100",
91244=>"011011011",
91245=>"100100111",
91246=>"001000000",
91247=>"000100110",
91248=>"001001001",
91249=>"011110110",
91250=>"111011011",
91251=>"011111001",
91252=>"100110011",
91253=>"100100010",
91254=>"111100100",
91255=>"000000001",
91256=>"111100111",
91257=>"011011011",
91258=>"000110111",
91259=>"110100110",
91260=>"011100100",
91261=>"010010000",
91262=>"111011000",
91263=>"000100111",
91264=>"000110000",
91265=>"000000000",
91266=>"010000011",
91267=>"011011001",
91268=>"100100100",
91269=>"010011011",
91270=>"100100011",
91271=>"011100101",
91272=>"100011110",
91273=>"001000010",
91274=>"101100111",
91275=>"011011010",
91276=>"000011011",
91277=>"100111111",
91278=>"011011011",
91279=>"100000010",
91280=>"000000000",
91281=>"010110110",
91282=>"111110110",
91283=>"011110111",
91284=>"011011000",
91285=>"110100100",
91286=>"000001001",
91287=>"000000001",
91288=>"000000000",
91289=>"000101011",
91290=>"011011110",
91291=>"000000000",
91292=>"001110110",
91293=>"101001101",
91294=>"111110010",
91295=>"001000100",
91296=>"010100101",
91297=>"100100110",
91298=>"010001011",
91299=>"010111000",
91300=>"100100100",
91301=>"011000110",
91302=>"111111000",
91303=>"011111011",
91304=>"101011111",
91305=>"000011011",
91306=>"000110100",
91307=>"110100000",
91308=>"011011000",
91309=>"111001001",
91310=>"110110111",
91311=>"111011011",
91312=>"001100010",
91313=>"001001001",
91314=>"111111100",
91315=>"110010110",
91316=>"010001001",
91317=>"000000000",
91318=>"011011100",
91319=>"001100100",
91320=>"110100100",
91321=>"001011000",
91322=>"110100000",
91323=>"011001000",
91324=>"000100001",
91325=>"000011011",
91326=>"011011001",
91327=>"000000000",
91328=>"100100100",
91329=>"000100000",
91330=>"000000011",
91331=>"001101011",
91332=>"011111111",
91333=>"001011010",
91334=>"011011001",
91335=>"111100100",
91336=>"011001010",
91337=>"111011001",
91338=>"011011101",
91339=>"000000111",
91340=>"111000011",
91341=>"001000110",
91342=>"011111101",
91343=>"011011010",
91344=>"110100100",
91345=>"100111111",
91346=>"010100100",
91347=>"111000011",
91348=>"011100000",
91349=>"111111111",
91350=>"000000110",
91351=>"110000000",
91352=>"110000000",
91353=>"011000000",
91354=>"000010110",
91355=>"100100100",
91356=>"011010100",
91357=>"011111001",
91358=>"010000010",
91359=>"000000000",
91360=>"010110100",
91361=>"100110100",
91362=>"100100100",
91363=>"011001010",
91364=>"100100100",
91365=>"011000000",
91366=>"111100100",
91367=>"001011011",
91368=>"110100100",
91369=>"011000100",
91370=>"100100110",
91371=>"101100101",
91372=>"010010010",
91373=>"111100100",
91374=>"000000000",
91375=>"011101011",
91376=>"001000000",
91377=>"111111001",
91378=>"111000000",
91379=>"001110100",
91380=>"010010010",
91381=>"000000001",
91382=>"110100000",
91383=>"000001000",
91384=>"100100100",
91385=>"111100011",
91386=>"010010110",
91387=>"111011011",
91388=>"011011011",
91389=>"001011010",
91390=>"000000000",
91391=>"000000100",
91392=>"011101000",
91393=>"000000000",
91394=>"000101111",
91395=>"110110111",
91396=>"000011100",
91397=>"000001000",
91398=>"011010100",
91399=>"110110000",
91400=>"010111111",
91401=>"011111111",
91402=>"011111110",
91403=>"000000000",
91404=>"111111111",
91405=>"010000001",
91406=>"001111011",
91407=>"111101111",
91408=>"001011111",
91409=>"111101101",
91410=>"100010010",
91411=>"111011000",
91412=>"010000000",
91413=>"111001000",
91414=>"011100111",
91415=>"000111111",
91416=>"001000001",
91417=>"000101111",
91418=>"101111111",
91419=>"000100000",
91420=>"100001001",
91421=>"011111111",
91422=>"111010010",
91423=>"000010100",
91424=>"000100000",
91425=>"000000000",
91426=>"111111101",
91427=>"100101111",
91428=>"001111001",
91429=>"110100100",
91430=>"111111000",
91431=>"001011111",
91432=>"000111000",
91433=>"100010000",
91434=>"111001011",
91435=>"011111011",
91436=>"111111111",
91437=>"011111111",
91438=>"111100000",
91439=>"010001001",
91440=>"001011000",
91441=>"100100000",
91442=>"110001111",
91443=>"110110110",
91444=>"000011001",
91445=>"110000000",
91446=>"000001001",
91447=>"000000001",
91448=>"100111110",
91449=>"101000001",
91450=>"101111111",
91451=>"111111111",
91452=>"000000001",
91453=>"111111111",
91454=>"111001000",
91455=>"000101110",
91456=>"100000000",
91457=>"000000010",
91458=>"000000000",
91459=>"000000100",
91460=>"111010000",
91461=>"111011000",
91462=>"110000000",
91463=>"111111111",
91464=>"111111001",
91465=>"101101101",
91466=>"101000000",
91467=>"101000000",
91468=>"001000101",
91469=>"110100100",
91470=>"000011011",
91471=>"111111110",
91472=>"000000000",
91473=>"000111000",
91474=>"111011111",
91475=>"111111001",
91476=>"010001011",
91477=>"000100001",
91478=>"110111101",
91479=>"000111111",
91480=>"111111101",
91481=>"001110010",
91482=>"001000001",
91483=>"100111001",
91484=>"010010111",
91485=>"011011001",
91486=>"000000000",
91487=>"000001001",
91488=>"000110110",
91489=>"000011111",
91490=>"101001000",
91491=>"100100110",
91492=>"111111111",
91493=>"011111111",
91494=>"110010000",
91495=>"111111111",
91496=>"101000001",
91497=>"101010000",
91498=>"001000000",
91499=>"111101000",
91500=>"000000000",
91501=>"001000000",
91502=>"001001101",
91503=>"010000000",
91504=>"000001000",
91505=>"010011111",
91506=>"000100100",
91507=>"011111111",
91508=>"010000111",
91509=>"001000111",
91510=>"110000000",
91511=>"010000000",
91512=>"000111001",
91513=>"000000111",
91514=>"000000101",
91515=>"110010011",
91516=>"110110110",
91517=>"111110100",
91518=>"110111111",
91519=>"110110101",
91520=>"111001000",
91521=>"000000000",
91522=>"000000000",
91523=>"000000011",
91524=>"100011111",
91525=>"101010000",
91526=>"011001000",
91527=>"011011011",
91528=>"100000001",
91529=>"101010000",
91530=>"010110100",
91531=>"111111000",
91532=>"000000010",
91533=>"000100000",
91534=>"000000101",
91535=>"111001101",
91536=>"111111110",
91537=>"101000000",
91538=>"011101111",
91539=>"111011111",
91540=>"110011111",
91541=>"000000000",
91542=>"111111111",
91543=>"011001000",
91544=>"000000000",
91545=>"000111111",
91546=>"111111111",
91547=>"000111111",
91548=>"000000000",
91549=>"000000000",
91550=>"011111000",
91551=>"010000000",
91552=>"001001000",
91553=>"011111100",
91554=>"011001100",
91555=>"101111111",
91556=>"011000001",
91557=>"110111111",
91558=>"111111111",
91559=>"000001001",
91560=>"011111010",
91561=>"100110110",
91562=>"101101101",
91563=>"010000000",
91564=>"110010010",
91565=>"110000000",
91566=>"111111000",
91567=>"111110000",
91568=>"000000000",
91569=>"011101100",
91570=>"100110000",
91571=>"100000000",
91572=>"011110010",
91573=>"011111011",
91574=>"111111110",
91575=>"110100001",
91576=>"001000000",
91577=>"010110110",
91578=>"111001111",
91579=>"000001101",
91580=>"111111111",
91581=>"000000000",
91582=>"000111111",
91583=>"011011011",
91584=>"111111111",
91585=>"111111001",
91586=>"111000000",
91587=>"011111101",
91588=>"010011010",
91589=>"100101000",
91590=>"111011110",
91591=>"000000001",
91592=>"111110000",
91593=>"110000011",
91594=>"111111001",
91595=>"111111111",
91596=>"111100000",
91597=>"011111111",
91598=>"000100111",
91599=>"101000000",
91600=>"110100000",
91601=>"001011011",
91602=>"111111111",
91603=>"011111111",
91604=>"110111111",
91605=>"100100100",
91606=>"100110111",
91607=>"010011110",
91608=>"110111111",
91609=>"000000011",
91610=>"100100000",
91611=>"000000111",
91612=>"010001100",
91613=>"000000011",
91614=>"111111011",
91615=>"111111111",
91616=>"110011011",
91617=>"110110100",
91618=>"010111011",
91619=>"010111110",
91620=>"111100110",
91621=>"000000000",
91622=>"000000000",
91623=>"100100100",
91624=>"000000101",
91625=>"111101111",
91626=>"110111111",
91627=>"111101111",
91628=>"000010010",
91629=>"110111111",
91630=>"111110000",
91631=>"111101111",
91632=>"000001111",
91633=>"001010000",
91634=>"111100111",
91635=>"111111111",
91636=>"010011011",
91637=>"001110111",
91638=>"101101111",
91639=>"010100100",
91640=>"000000000",
91641=>"111111110",
91642=>"000001001",
91643=>"010100100",
91644=>"000111111",
91645=>"001000000",
91646=>"001001001",
91647=>"000100000",
91648=>"110110111",
91649=>"000000101",
91650=>"111011001",
91651=>"101101111",
91652=>"111000101",
91653=>"000001001",
91654=>"000001010",
91655=>"111111101",
91656=>"111101111",
91657=>"010000011",
91658=>"000010000",
91659=>"100011110",
91660=>"101000101",
91661=>"111111111",
91662=>"100010010",
91663=>"111111110",
91664=>"111111111",
91665=>"111111111",
91666=>"010110000",
91667=>"000001111",
91668=>"111101111",
91669=>"110000111",
91670=>"000000000",
91671=>"000111000",
91672=>"110000000",
91673=>"000011000",
91674=>"100000000",
91675=>"101100100",
91676=>"000100110",
91677=>"101111111",
91678=>"011111101",
91679=>"101000111",
91680=>"101110111",
91681=>"010111011",
91682=>"000000000",
91683=>"010001111",
91684=>"000111111",
91685=>"011101110",
91686=>"100111000",
91687=>"000000011",
91688=>"101111000",
91689=>"111111001",
91690=>"000101000",
91691=>"011000111",
91692=>"000111011",
91693=>"110111001",
91694=>"000111000",
91695=>"110000110",
91696=>"111110000",
91697=>"001110000",
91698=>"010000000",
91699=>"011111111",
91700=>"000010000",
91701=>"010011111",
91702=>"100000000",
91703=>"111010111",
91704=>"101000111",
91705=>"001000110",
91706=>"000000000",
91707=>"000010011",
91708=>"001111110",
91709=>"001000000",
91710=>"111111110",
91711=>"000001010",
91712=>"111111100",
91713=>"001000011",
91714=>"010100010",
91715=>"010100100",
91716=>"101001110",
91717=>"111000101",
91718=>"000001011",
91719=>"101110111",
91720=>"001111010",
91721=>"100011101",
91722=>"111001000",
91723=>"111001000",
91724=>"110010110",
91725=>"001111111",
91726=>"010111010",
91727=>"000101101",
91728=>"111110111",
91729=>"101111101",
91730=>"001101111",
91731=>"101111000",
91732=>"001000010",
91733=>"100000000",
91734=>"000000010",
91735=>"111101100",
91736=>"011011110",
91737=>"110100000",
91738=>"000000110",
91739=>"111011000",
91740=>"101101110",
91741=>"100100001",
91742=>"101101111",
91743=>"010000001",
91744=>"000000000",
91745=>"011000100",
91746=>"011000110",
91747=>"000001001",
91748=>"011001100",
91749=>"000111010",
91750=>"000000001",
91751=>"000001111",
91752=>"000100111",
91753=>"000000000",
91754=>"000100001",
91755=>"001000101",
91756=>"000111000",
91757=>"111111011",
91758=>"110000111",
91759=>"000111001",
91760=>"110000000",
91761=>"111000000",
91762=>"010010000",
91763=>"000100001",
91764=>"100000010",
91765=>"101000000",
91766=>"001000001",
91767=>"111001101",
91768=>"101111001",
91769=>"011111000",
91770=>"000001011",
91771=>"110111000",
91772=>"011011110",
91773=>"000001000",
91774=>"111111011",
91775=>"000000011",
91776=>"111111000",
91777=>"000011001",
91778=>"000000110",
91779=>"101100010",
91780=>"001101000",
91781=>"000010000",
91782=>"111001011",
91783=>"000001110",
91784=>"011000000",
91785=>"000000000",
91786=>"111111111",
91787=>"000010011",
91788=>"011001111",
91789=>"110010110",
91790=>"111000000",
91791=>"000000000",
91792=>"000101100",
91793=>"010000000",
91794=>"011111000",
91795=>"100101001",
91796=>"101000101",
91797=>"110111111",
91798=>"000111011",
91799=>"111100000",
91800=>"011111101",
91801=>"111100011",
91802=>"110111111",
91803=>"111001000",
91804=>"101101101",
91805=>"111110000",
91806=>"000110111",
91807=>"000111110",
91808=>"000000000",
91809=>"111111111",
91810=>"101111110",
91811=>"011110111",
91812=>"000111000",
91813=>"011011000",
91814=>"111001001",
91815=>"010000100",
91816=>"111111111",
91817=>"111001001",
91818=>"111100001",
91819=>"000010111",
91820=>"111100001",
91821=>"111100100",
91822=>"111111111",
91823=>"100101000",
91824=>"111000100",
91825=>"001011011",
91826=>"000111010",
91827=>"000000000",
91828=>"010111000",
91829=>"101010101",
91830=>"011001000",
91831=>"001000010",
91832=>"100111011",
91833=>"001001011",
91834=>"000000000",
91835=>"011000000",
91836=>"100000011",
91837=>"000001100",
91838=>"011000110",
91839=>"010010000",
91840=>"000101101",
91841=>"000000000",
91842=>"110100111",
91843=>"000000000",
91844=>"110000000",
91845=>"000111111",
91846=>"010111000",
91847=>"000011101",
91848=>"010010011",
91849=>"001000000",
91850=>"111010111",
91851=>"101001000",
91852=>"001000010",
91853=>"111110111",
91854=>"010010110",
91855=>"110000101",
91856=>"111101000",
91857=>"010011001",
91858=>"111111111",
91859=>"101001110",
91860=>"111000111",
91861=>"000000011",
91862=>"101001111",
91863=>"001111110",
91864=>"001111011",
91865=>"111001110",
91866=>"000000000",
91867=>"011110000",
91868=>"000000000",
91869=>"110000111",
91870=>"000110000",
91871=>"001100001",
91872=>"101000001",
91873=>"001111111",
91874=>"000001011",
91875=>"111101001",
91876=>"101000000",
91877=>"111010011",
91878=>"101100111",
91879=>"111110111",
91880=>"001000010",
91881=>"101000101",
91882=>"010010110",
91883=>"001000111",
91884=>"111000100",
91885=>"000000000",
91886=>"111000000",
91887=>"110000110",
91888=>"000000000",
91889=>"001100111",
91890=>"000101101",
91891=>"101111110",
91892=>"000100101",
91893=>"000000000",
91894=>"110000110",
91895=>"001011011",
91896=>"011111111",
91897=>"000010001",
91898=>"111111000",
91899=>"100000000",
91900=>"010111111",
91901=>"101101010",
91902=>"000001011",
91903=>"111111110",
91904=>"001101001",
91905=>"010000010",
91906=>"111100100",
91907=>"000100111",
91908=>"111011001",
91909=>"111001010",
91910=>"100101100",
91911=>"101101010",
91912=>"100110111",
91913=>"000111000",
91914=>"111100001",
91915=>"000000000",
91916=>"101000000",
91917=>"111101101",
91918=>"000111111",
91919=>"101011100",
91920=>"011000110",
91921=>"000010011",
91922=>"101000111",
91923=>"000000010",
91924=>"111101111",
91925=>"000000000",
91926=>"100100100",
91927=>"110011010",
91928=>"111100001",
91929=>"000111011",
91930=>"000000100",
91931=>"100100101",
91932=>"000010011",
91933=>"000000100",
91934=>"001000000",
91935=>"100100101",
91936=>"010010000",
91937=>"010011000",
91938=>"000000100",
91939=>"100011011",
91940=>"010000010",
91941=>"110111111",
91942=>"010000000",
91943=>"101010111",
91944=>"011011011",
91945=>"010111010",
91946=>"000011000",
91947=>"111000101",
91948=>"000100000",
91949=>"101000011",
91950=>"110100100",
91951=>"010110010",
91952=>"111100000",
91953=>"101111111",
91954=>"000011100",
91955=>"011011010",
91956=>"111000000",
91957=>"111111110",
91958=>"100110000",
91959=>"010111011",
91960=>"111111110",
91961=>"000000000",
91962=>"011101111",
91963=>"000010011",
91964=>"000111110",
91965=>"111111001",
91966=>"100000100",
91967=>"110011000",
91968=>"001010011",
91969=>"010011000",
91970=>"010111110",
91971=>"010110100",
91972=>"000010000",
91973=>"000000000",
91974=>"000111000",
91975=>"111101100",
91976=>"100000100",
91977=>"100100111",
91978=>"101101101",
91979=>"011001100",
91980=>"000111111",
91981=>"101111111",
91982=>"000111111",
91983=>"111001011",
91984=>"000000101",
91985=>"110111100",
91986=>"111110100",
91987=>"011001000",
91988=>"011000000",
91989=>"010110100",
91990=>"000111011",
91991=>"000000000",
91992=>"101110101",
91993=>"100100000",
91994=>"100110100",
91995=>"011100111",
91996=>"000000010",
91997=>"110101101",
91998=>"111111100",
91999=>"011011000",
92000=>"000110010",
92001=>"100100110",
92002=>"100000110",
92003=>"011001000",
92004=>"000111010",
92005=>"000100000",
92006=>"110000100",
92007=>"000111011",
92008=>"111000000",
92009=>"111101111",
92010=>"111000001",
92011=>"111011011",
92012=>"111000000",
92013=>"111000111",
92014=>"000011011",
92015=>"111000011",
92016=>"101110010",
92017=>"011000011",
92018=>"001000000",
92019=>"100100000",
92020=>"000010011",
92021=>"010000000",
92022=>"000010010",
92023=>"011111011",
92024=>"011000000",
92025=>"100100100",
92026=>"100000100",
92027=>"111111111",
92028=>"000110110",
92029=>"011000000",
92030=>"111101100",
92031=>"100000000",
92032=>"011000000",
92033=>"100100000",
92034=>"010011011",
92035=>"111100111",
92036=>"111001000",
92037=>"000100000",
92038=>"011111110",
92039=>"000011011",
92040=>"100001110",
92041=>"000000000",
92042=>"111101100",
92043=>"111111010",
92044=>"000111010",
92045=>"100011111",
92046=>"000010000",
92047=>"111101001",
92048=>"111111010",
92049=>"000000010",
92050=>"010010011",
92051=>"001000000",
92052=>"000001011",
92053=>"011010010",
92054=>"110110000",
92055=>"100011011",
92056=>"011011001",
92057=>"000100100",
92058=>"011011000",
92059=>"111100100",
92060=>"000100100",
92061=>"011011110",
92062=>"001000000",
92063=>"100100100",
92064=>"111001100",
92065=>"011101100",
92066=>"111101010",
92067=>"111000100",
92068=>"011000011",
92069=>"100011111",
92070=>"000011011",
92071=>"010011111",
92072=>"011010001",
92073=>"101000111",
92074=>"011011000",
92075=>"110000111",
92076=>"011001000",
92077=>"100110111",
92078=>"010000000",
92079=>"000100000",
92080=>"011001010",
92081=>"010000000",
92082=>"101100110",
92083=>"000110011",
92084=>"001100111",
92085=>"101111001",
92086=>"011011011",
92087=>"000011011",
92088=>"000011011",
92089=>"000011011",
92090=>"100011011",
92091=>"111111000",
92092=>"111111111",
92093=>"011011011",
92094=>"011011000",
92095=>"010000100",
92096=>"011000111",
92097=>"000011111",
92098=>"000000000",
92099=>"101101101",
92100=>"011011111",
92101=>"110000000",
92102=>"010001111",
92103=>"100011001",
92104=>"000101111",
92105=>"011000000",
92106=>"111111111",
92107=>"111001000",
92108=>"000011011",
92109=>"000001010",
92110=>"000010000",
92111=>"011000011",
92112=>"100111011",
92113=>"010110110",
92114=>"000010010",
92115=>"010111011",
92116=>"111111010",
92117=>"000000011",
92118=>"100000100",
92119=>"100100000",
92120=>"111101000",
92121=>"111100111",
92122=>"111100010",
92123=>"111101111",
92124=>"100100100",
92125=>"000000101",
92126=>"011111111",
92127=>"011001001",
92128=>"100100100",
92129=>"101100100",
92130=>"011101111",
92131=>"111100000",
92132=>"111100000",
92133=>"010000010",
92134=>"011000111",
92135=>"011000000",
92136=>"111101110",
92137=>"010000100",
92138=>"100100100",
92139=>"110000111",
92140=>"001001000",
92141=>"000011011",
92142=>"000000000",
92143=>"000000010",
92144=>"000000000",
92145=>"000000100",
92146=>"010001101",
92147=>"101111111",
92148=>"000100100",
92149=>"111100000",
92150=>"000001011",
92151=>"100101100",
92152=>"011000000",
92153=>"111011110",
92154=>"111100100",
92155=>"000000101",
92156=>"000000000",
92157=>"011000000",
92158=>"011111100",
92159=>"101100100",
92160=>"000010001",
92161=>"000000010",
92162=>"010011100",
92163=>"010001001",
92164=>"101100000",
92165=>"000001001",
92166=>"011001100",
92167=>"011010011",
92168=>"010000000",
92169=>"000010010",
92170=>"010000000",
92171=>"010001000",
92172=>"001001001",
92173=>"101101001",
92174=>"100001000",
92175=>"111011001",
92176=>"010010000",
92177=>"011011000",
92178=>"000100110",
92179=>"000000011",
92180=>"011001001",
92181=>"000001111",
92182=>"010011101",
92183=>"001111011",
92184=>"001100100",
92185=>"111111100",
92186=>"011001001",
92187=>"111001001",
92188=>"011101111",
92189=>"000100000",
92190=>"011101001",
92191=>"010010000",
92192=>"011001001",
92193=>"000100101",
92194=>"111001000",
92195=>"110011011",
92196=>"100110100",
92197=>"010000101",
92198=>"010110010",
92199=>"101101000",
92200=>"110110011",
92201=>"010010000",
92202=>"100111011",
92203=>"000000001",
92204=>"111111110",
92205=>"001001100",
92206=>"011111100",
92207=>"100100010",
92208=>"111001000",
92209=>"110100000",
92210=>"011000000",
92211=>"111110011",
92212=>"011001000",
92213=>"010001010",
92214=>"100000100",
92215=>"001101000",
92216=>"000100100",
92217=>"001100100",
92218=>"000100100",
92219=>"001010000",
92220=>"000000011",
92221=>"110110010",
92222=>"011001001",
92223=>"000100110",
92224=>"001001101",
92225=>"011000100",
92226=>"110110011",
92227=>"000001001",
92228=>"000111001",
92229=>"001001000",
92230=>"110110010",
92231=>"111111111",
92232=>"000100011",
92233=>"111010010",
92234=>"011001001",
92235=>"001110110",
92236=>"000000100",
92237=>"101110010",
92238=>"000000110",
92239=>"111010011",
92240=>"000001000",
92241=>"110110110",
92242=>"011001001",
92243=>"000011010",
92244=>"010111111",
92245=>"111000000",
92246=>"000100111",
92247=>"010010111",
92248=>"011111111",
92249=>"000110000",
92250=>"101000010",
92251=>"110100110",
92252=>"011001000",
92253=>"000000100",
92254=>"111111011",
92255=>"011010000",
92256=>"100100000",
92257=>"011001001",
92258=>"100011111",
92259=>"000101101",
92260=>"110110110",
92261=>"100100000",
92262=>"111111000",
92263=>"110110010",
92264=>"110010101",
92265=>"100100111",
92266=>"000111011",
92267=>"111111011",
92268=>"110011111",
92269=>"101101111",
92270=>"000000000",
92271=>"010100100",
92272=>"101110010",
92273=>"010100100",
92274=>"110011010",
92275=>"011000000",
92276=>"110100110",
92277=>"000101001",
92278=>"111110011",
92279=>"000110110",
92280=>"011001001",
92281=>"011000110",
92282=>"100101011",
92283=>"001001111",
92284=>"101100110",
92285=>"111001001",
92286=>"010000111",
92287=>"000011000",
92288=>"010110001",
92289=>"100100101",
92290=>"001001001",
92291=>"000100000",
92292=>"000110101",
92293=>"110111000",
92294=>"001000100",
92295=>"010010000",
92296=>"110100101",
92297=>"001010000",
92298=>"001111000",
92299=>"111001000",
92300=>"100000011",
92301=>"100011011",
92302=>"011011110",
92303=>"001000001",
92304=>"000110110",
92305=>"000010011",
92306=>"000110000",
92307=>"100000000",
92308=>"000110010",
92309=>"011000001",
92310=>"010110111",
92311=>"000000000",
92312=>"111000010",
92313=>"110000010",
92314=>"110100000",
92315=>"110100000",
92316=>"001001001",
92317=>"000001010",
92318=>"011001110",
92319=>"100101111",
92320=>"000100000",
92321=>"011000001",
92322=>"110100100",
92323=>"010011001",
92324=>"110111111",
92325=>"101011001",
92326=>"111000000",
92327=>"110111001",
92328=>"011011011",
92329=>"001100100",
92330=>"100000000",
92331=>"000000001",
92332=>"001011111",
92333=>"110100010",
92334=>"011000000",
92335=>"111011001",
92336=>"000000111",
92337=>"011001110",
92338=>"000101100",
92339=>"000100110",
92340=>"100110011",
92341=>"111100010",
92342=>"000100110",
92343=>"010000000",
92344=>"000100000",
92345=>"111000110",
92346=>"011011001",
92347=>"000100011",
92348=>"100100000",
92349=>"110110011",
92350=>"101110011",
92351=>"011011100",
92352=>"011001000",
92353=>"011011000",
92354=>"011100110",
92355=>"010110000",
92356=>"001100100",
92357=>"111111100",
92358=>"010100111",
92359=>"011010001",
92360=>"000000001",
92361=>"000100000",
92362=>"100110110",
92363=>"011011010",
92364=>"000011011",
92365=>"110000101",
92366=>"001000000",
92367=>"010100000",
92368=>"100110111",
92369=>"001000010",
92370=>"000010000",
92371=>"111011011",
92372=>"100000101",
92373=>"011101000",
92374=>"001000100",
92375=>"010001000",
92376=>"101110010",
92377=>"111000111",
92378=>"101001110",
92379=>"101001001",
92380=>"111100100",
92381=>"000110111",
92382=>"001111111",
92383=>"011000001",
92384=>"011011001",
92385=>"101001001",
92386=>"100111011",
92387=>"100110110",
92388=>"010000001",
92389=>"110110100",
92390=>"111000111",
92391=>"100100111",
92392=>"111101111",
92393=>"011100000",
92394=>"111100010",
92395=>"100110011",
92396=>"011001001",
92397=>"000000000",
92398=>"000001001",
92399=>"000000100",
92400=>"100011011",
92401=>"000000100",
92402=>"011001001",
92403=>"110101110",
92404=>"111001001",
92405=>"100110011",
92406=>"000001000",
92407=>"100100110",
92408=>"001001001",
92409=>"100000000",
92410=>"011001000",
92411=>"100110110",
92412=>"011010110",
92413=>"110100011",
92414=>"100100111",
92415=>"011110111",
92416=>"000000011",
92417=>"001000111",
92418=>"000010111",
92419=>"000000100",
92420=>"000111111",
92421=>"101001100",
92422=>"110100010",
92423=>"000111010",
92424=>"010000000",
92425=>"010011001",
92426=>"111111110",
92427=>"000000000",
92428=>"001000000",
92429=>"000000110",
92430=>"011100100",
92431=>"110110101",
92432=>"000111011",
92433=>"010110110",
92434=>"000000101",
92435=>"111111111",
92436=>"000000111",
92437=>"000000000",
92438=>"100000100",
92439=>"011111111",
92440=>"000000011",
92441=>"000000001",
92442=>"011000000",
92443=>"000000111",
92444=>"110010010",
92445=>"010101111",
92446=>"000010010",
92447=>"001000000",
92448=>"000010000",
92449=>"001111111",
92450=>"000000111",
92451=>"111101111",
92452=>"111100100",
92453=>"000101000",
92454=>"000111011",
92455=>"000111111",
92456=>"000111111",
92457=>"011100000",
92458=>"000000000",
92459=>"100000101",
92460=>"100110111",
92461=>"111010110",
92462=>"000110111",
92463=>"001001000",
92464=>"110111111",
92465=>"101111011",
92466=>"000101000",
92467=>"010010000",
92468=>"001111111",
92469=>"011111101",
92470=>"000100011",
92471=>"000001101",
92472=>"111111001",
92473=>"001000111",
92474=>"111000000",
92475=>"010011000",
92476=>"011011111",
92477=>"101100101",
92478=>"110000000",
92479=>"100011111",
92480=>"111111000",
92481=>"000110000",
92482=>"111000000",
92483=>"110011011",
92484=>"111000000",
92485=>"001010011",
92486=>"111011110",
92487=>"001000000",
92488=>"001001011",
92489=>"000111111",
92490=>"001100111",
92491=>"010011000",
92492=>"111000000",
92493=>"011111111",
92494=>"001111110",
92495=>"111101100",
92496=>"000000111",
92497=>"111000000",
92498=>"010000001",
92499=>"010101100",
92500=>"000010110",
92501=>"100110111",
92502=>"111011011",
92503=>"000111111",
92504=>"111000000",
92505=>"010000000",
92506=>"111000000",
92507=>"010000000",
92508=>"111111111",
92509=>"110110000",
92510=>"111111000",
92511=>"011110111",
92512=>"111001000",
92513=>"011000010",
92514=>"001000000",
92515=>"111011000",
92516=>"111101000",
92517=>"101100000",
92518=>"000111011",
92519=>"000000000",
92520=>"001111101",
92521=>"111111000",
92522=>"111111000",
92523=>"000000000",
92524=>"111111001",
92525=>"110111111",
92526=>"111101111",
92527=>"000000001",
92528=>"001100110",
92529=>"111000000",
92530=>"001001001",
92531=>"000101000",
92532=>"001101111",
92533=>"000000000",
92534=>"111101000",
92535=>"000011000",
92536=>"000000111",
92537=>"000000101",
92538=>"111101000",
92539=>"010111111",
92540=>"111100111",
92541=>"010100000",
92542=>"000101000",
92543=>"000000110",
92544=>"010001000",
92545=>"010011111",
92546=>"000001111",
92547=>"001000101",
92548=>"010110111",
92549=>"111000001",
92550=>"000110000",
92551=>"111100000",
92552=>"101001011",
92553=>"110011000",
92554=>"000100011",
92555=>"000000010",
92556=>"111000000",
92557=>"110000000",
92558=>"111000000",
92559=>"110110000",
92560=>"011101111",
92561=>"001001000",
92562=>"100000000",
92563=>"001000110",
92564=>"000001111",
92565=>"111110000",
92566=>"011000000",
92567=>"111110100",
92568=>"010000000",
92569=>"000000010",
92570=>"010011011",
92571=>"000100010",
92572=>"111000000",
92573=>"101110111",
92574=>"100000000",
92575=>"000000101",
92576=>"001101111",
92577=>"111010101",
92578=>"111101001",
92579=>"111000000",
92580=>"111111101",
92581=>"000000011",
92582=>"111100100",
92583=>"110000000",
92584=>"111110111",
92585=>"111111001",
92586=>"111000000",
92587=>"000000101",
92588=>"011000111",
92589=>"000111111",
92590=>"011011111",
92591=>"011000000",
92592=>"101001001",
92593=>"111100000",
92594=>"101111110",
92595=>"001000101",
92596=>"011111110",
92597=>"111001000",
92598=>"000100111",
92599=>"000110000",
92600=>"100110100",
92601=>"000010111",
92602=>"000000000",
92603=>"000011111",
92604=>"100011000",
92605=>"111111111",
92606=>"110100111",
92607=>"100000000",
92608=>"000010111",
92609=>"111000000",
92610=>"001101111",
92611=>"000100100",
92612=>"000111101",
92613=>"111000001",
92614=>"101111111",
92615=>"100000000",
92616=>"000000110",
92617=>"111001111",
92618=>"111001001",
92619=>"000010000",
92620=>"000010000",
92621=>"110011111",
92622=>"000000111",
92623=>"000000111",
92624=>"000111111",
92625=>"111011000",
92626=>"001001011",
92627=>"101000001",
92628=>"110000000",
92629=>"011011011",
92630=>"111100000",
92631=>"000000001",
92632=>"000111000",
92633=>"010111101",
92634=>"000000101",
92635=>"100000000",
92636=>"001011001",
92637=>"000100000",
92638=>"111000000",
92639=>"001110111",
92640=>"000000111",
92641=>"011000111",
92642=>"000111111",
92643=>"000101110",
92644=>"100000000",
92645=>"011000001",
92646=>"111010111",
92647=>"110110011",
92648=>"111111000",
92649=>"011000101",
92650=>"110110111",
92651=>"111100000",
92652=>"001111111",
92653=>"000111111",
92654=>"010010110",
92655=>"111101000",
92656=>"000001000",
92657=>"111000100",
92658=>"111001000",
92659=>"111001000",
92660=>"000000110",
92661=>"111000000",
92662=>"111000000",
92663=>"000000000",
92664=>"000111111",
92665=>"111111101",
92666=>"100000111",
92667=>"111110000",
92668=>"110000010",
92669=>"001000000",
92670=>"111011111",
92671=>"111111100",
92672=>"010101100",
92673=>"010011010",
92674=>"001000000",
92675=>"010001001",
92676=>"010110011",
92677=>"000101111",
92678=>"000010011",
92679=>"111101000",
92680=>"101000000",
92681=>"011011010",
92682=>"010111111",
92683=>"111001001",
92684=>"111001001",
92685=>"100000001",
92686=>"111111111",
92687=>"111111111",
92688=>"010010000",
92689=>"110010000",
92690=>"110100111",
92691=>"000000000",
92692=>"100001000",
92693=>"101000000",
92694=>"000000011",
92695=>"111100111",
92696=>"010100010",
92697=>"100111011",
92698=>"100100000",
92699=>"000001001",
92700=>"000101000",
92701=>"111111000",
92702=>"000001111",
92703=>"000000000",
92704=>"000000000",
92705=>"010110010",
92706=>"110000000",
92707=>"100000000",
92708=>"000000000",
92709=>"110111001",
92710=>"101000000",
92711=>"100111110",
92712=>"000001000",
92713=>"101001000",
92714=>"011001000",
92715=>"000000100",
92716=>"111110010",
92717=>"111101101",
92718=>"000000111",
92719=>"000110110",
92720=>"000000000",
92721=>"001011000",
92722=>"000001111",
92723=>"100010110",
92724=>"000111111",
92725=>"011000000",
92726=>"111010001",
92727=>"101101100",
92728=>"111111101",
92729=>"101000111",
92730=>"001000000",
92731=>"000111001",
92732=>"111001011",
92733=>"010111011",
92734=>"000000000",
92735=>"111111111",
92736=>"000000111",
92737=>"100110110",
92738=>"010000111",
92739=>"111111110",
92740=>"111100000",
92741=>"000100001",
92742=>"000000000",
92743=>"000000000",
92744=>"001101001",
92745=>"000111011",
92746=>"101000101",
92747=>"111111001",
92748=>"111000000",
92749=>"000000000",
92750=>"100011100",
92751=>"101000000",
92752=>"001001000",
92753=>"110111111",
92754=>"000000001",
92755=>"001001000",
92756=>"000111010",
92757=>"001000100",
92758=>"110110110",
92759=>"111000110",
92760=>"101101011",
92761=>"011111110",
92762=>"110010000",
92763=>"111111111",
92764=>"000010111",
92765=>"000000100",
92766=>"000111110",
92767=>"111111011",
92768=>"111101000",
92769=>"110111111",
92770=>"000111011",
92771=>"111111010",
92772=>"011001011",
92773=>"011111111",
92774=>"110111000",
92775=>"001111011",
92776=>"111001000",
92777=>"111111010",
92778=>"000110111",
92779=>"100101001",
92780=>"110000001",
92781=>"011111111",
92782=>"000000000",
92783=>"111000110",
92784=>"010110110",
92785=>"111111111",
92786=>"010000000",
92787=>"010110110",
92788=>"100001000",
92789=>"101101101",
92790=>"111111111",
92791=>"111111011",
92792=>"000000000",
92793=>"000000010",
92794=>"000111111",
92795=>"101000111",
92796=>"111011101",
92797=>"100000010",
92798=>"000000000",
92799=>"101111111",
92800=>"111000010",
92801=>"111110000",
92802=>"010010011",
92803=>"000000000",
92804=>"101111111",
92805=>"100000000",
92806=>"011011100",
92807=>"110010011",
92808=>"100011000",
92809=>"111011000",
92810=>"000000000",
92811=>"001000000",
92812=>"000111111",
92813=>"001010010",
92814=>"111001011",
92815=>"101000000",
92816=>"000110110",
92817=>"001101111",
92818=>"111111001",
92819=>"000010000",
92820=>"111001001",
92821=>"010010010",
92822=>"111111010",
92823=>"110100100",
92824=>"001101001",
92825=>"111011000",
92826=>"000000000",
92827=>"000000000",
92828=>"000000000",
92829=>"101000000",
92830=>"111101000",
92831=>"111000111",
92832=>"001001001",
92833=>"110011110",
92834=>"000000000",
92835=>"000000111",
92836=>"000000110",
92837=>"000000110",
92838=>"111001000",
92839=>"100000000",
92840=>"010111011",
92841=>"111100100",
92842=>"000000000",
92843=>"111110110",
92844=>"110110100",
92845=>"010100101",
92846=>"111111111",
92847=>"000000010",
92848=>"000000101",
92849=>"000110110",
92850=>"000011011",
92851=>"000100111",
92852=>"000101111",
92853=>"100000000",
92854=>"001000000",
92855=>"010110000",
92856=>"010011111",
92857=>"111011011",
92858=>"000111111",
92859=>"000000000",
92860=>"000011111",
92861=>"111111111",
92862=>"100101111",
92863=>"111110110",
92864=>"010010111",
92865=>"000000100",
92866=>"001001001",
92867=>"001000000",
92868=>"000000001",
92869=>"111100000",
92870=>"000000001",
92871=>"000000111",
92872=>"101100010",
92873=>"111000000",
92874=>"000000101",
92875=>"101000000",
92876=>"010111111",
92877=>"110110100",
92878=>"000010010",
92879=>"000101111",
92880=>"010110000",
92881=>"011011011",
92882=>"000010101",
92883=>"011111111",
92884=>"001111111",
92885=>"000000000",
92886=>"101000101",
92887=>"111010000",
92888=>"000000001",
92889=>"000110010",
92890=>"011000010",
92891=>"101000110",
92892=>"000000010",
92893=>"001100111",
92894=>"010111110",
92895=>"010111011",
92896=>"000010010",
92897=>"100110111",
92898=>"000111111",
92899=>"011111110",
92900=>"011111110",
92901=>"000111000",
92902=>"101001011",
92903=>"000111111",
92904=>"101011011",
92905=>"000100000",
92906=>"011111111",
92907=>"111111111",
92908=>"111101001",
92909=>"100001000",
92910=>"000000100",
92911=>"000001111",
92912=>"111101111",
92913=>"101001000",
92914=>"001000111",
92915=>"110001111",
92916=>"000010111",
92917=>"000010000",
92918=>"010111000",
92919=>"001000111",
92920=>"000110111",
92921=>"111000000",
92922=>"111101111",
92923=>"111110100",
92924=>"001000001",
92925=>"010111111",
92926=>"000000000",
92927=>"111000000",
92928=>"000110111",
92929=>"000000000",
92930=>"111000001",
92931=>"111011111",
92932=>"111011110",
92933=>"100000111",
92934=>"000000000",
92935=>"010111010",
92936=>"111111000",
92937=>"000000001",
92938=>"100101111",
92939=>"100101000",
92940=>"001101111",
92941=>"010100101",
92942=>"000010111",
92943=>"000000111",
92944=>"010111111",
92945=>"100100001",
92946=>"100010111",
92947=>"110000000",
92948=>"010111110",
92949=>"110010110",
92950=>"101101001",
92951=>"001111101",
92952=>"101110011",
92953=>"011100110",
92954=>"000001011",
92955=>"111000101",
92956=>"000011110",
92957=>"000100000",
92958=>"101101111",
92959=>"000000000",
92960=>"101100100",
92961=>"011101110",
92962=>"000000101",
92963=>"000111111",
92964=>"110110011",
92965=>"101101001",
92966=>"100101111",
92967=>"000100000",
92968=>"101111111",
92969=>"000101000",
92970=>"001100001",
92971=>"000010101",
92972=>"111111010",
92973=>"101010111",
92974=>"000101111",
92975=>"110110000",
92976=>"011110011",
92977=>"111000100",
92978=>"000001000",
92979=>"000111110",
92980=>"000000101",
92981=>"001101011",
92982=>"000110100",
92983=>"000110000",
92984=>"111111000",
92985=>"000001111",
92986=>"000000000",
92987=>"101000010",
92988=>"000000101",
92989=>"111010010",
92990=>"000000101",
92991=>"110100101",
92992=>"100000000",
92993=>"100101011",
92994=>"000000000",
92995=>"111111111",
92996=>"100101111",
92997=>"000000101",
92998=>"001111000",
92999=>"010000000",
93000=>"000100010",
93001=>"010111010",
93002=>"000101000",
93003=>"001110101",
93004=>"100000111",
93005=>"001100110",
93006=>"110100011",
93007=>"010000111",
93008=>"100110100",
93009=>"111010110",
93010=>"100010001",
93011=>"000000011",
93012=>"000000100",
93013=>"001000000",
93014=>"000010011",
93015=>"010110111",
93016=>"101111110",
93017=>"001000001",
93018=>"011001011",
93019=>"001010010",
93020=>"100111110",
93021=>"101000101",
93022=>"111000111",
93023=>"101101111",
93024=>"000000000",
93025=>"000100000",
93026=>"000000001",
93027=>"111110111",
93028=>"000010010",
93029=>"000100000",
93030=>"110110000",
93031=>"111101011",
93032=>"010011011",
93033=>"100111010",
93034=>"100101010",
93035=>"101100111",
93036=>"001100111",
93037=>"101111111",
93038=>"000000000",
93039=>"111111111",
93040=>"110100100",
93041=>"101001011",
93042=>"000111110",
93043=>"101000000",
93044=>"111010010",
93045=>"000100100",
93046=>"010000000",
93047=>"010110100",
93048=>"100100111",
93049=>"111100110",
93050=>"000000101",
93051=>"111111101",
93052=>"000000001",
93053=>"001001111",
93054=>"000000011",
93055=>"000000011",
93056=>"000000010",
93057=>"101001111",
93058=>"010011000",
93059=>"111000000",
93060=>"111111111",
93061=>"000001001",
93062=>"100011100",
93063=>"000100001",
93064=>"001110010",
93065=>"011010010",
93066=>"100111110",
93067=>"100100000",
93068=>"100000000",
93069=>"000100100",
93070=>"100000010",
93071=>"000000000",
93072=>"110001000",
93073=>"111100100",
93074=>"000101111",
93075=>"001010101",
93076=>"111111010",
93077=>"011000101",
93078=>"101011001",
93079=>"000100100",
93080=>"000000010",
93081=>"100100100",
93082=>"011000000",
93083=>"010000000",
93084=>"000000100",
93085=>"011010000",
93086=>"111100111",
93087=>"100000010",
93088=>"111101011",
93089=>"111111111",
93090=>"010101111",
93091=>"011111111",
93092=>"011010101",
93093=>"000010111",
93094=>"100111000",
93095=>"111000000",
93096=>"000000001",
93097=>"000000000",
93098=>"011100100",
93099=>"000101101",
93100=>"110110111",
93101=>"000010001",
93102=>"000111011",
93103=>"001111111",
93104=>"011010100",
93105=>"000000000",
93106=>"100000000",
93107=>"101010011",
93108=>"011011111",
93109=>"001000000",
93110=>"000000100",
93111=>"000000000",
93112=>"000100101",
93113=>"000010110",
93114=>"010000011",
93115=>"010010111",
93116=>"101011111",
93117=>"111000000",
93118=>"000000000",
93119=>"010111000",
93120=>"100100000",
93121=>"100000010",
93122=>"010010000",
93123=>"011001000",
93124=>"000011001",
93125=>"001111010",
93126=>"010111000",
93127=>"110100011",
93128=>"000101011",
93129=>"001101101",
93130=>"010010010",
93131=>"100111111",
93132=>"011011000",
93133=>"000000100",
93134=>"100111000",
93135=>"011111111",
93136=>"111110010",
93137=>"001101111",
93138=>"101111011",
93139=>"100110111",
93140=>"111100101",
93141=>"000100100",
93142=>"100000101",
93143=>"100000000",
93144=>"111110000",
93145=>"001011011",
93146=>"111110011",
93147=>"101000000",
93148=>"001100100",
93149=>"001101101",
93150=>"100000100",
93151=>"000001111",
93152=>"111110111",
93153=>"000100000",
93154=>"111111111",
93155=>"100010011",
93156=>"101000010",
93157=>"011011000",
93158=>"101011111",
93159=>"110100110",
93160=>"100100111",
93161=>"110001000",
93162=>"100110111",
93163=>"000111111",
93164=>"111000000",
93165=>"000101111",
93166=>"100000000",
93167=>"111011100",
93168=>"101111111",
93169=>"101101111",
93170=>"000000001",
93171=>"110010100",
93172=>"000000111",
93173=>"101101010",
93174=>"100000111",
93175=>"111010100",
93176=>"111000000",
93177=>"010001011",
93178=>"001101111",
93179=>"000001000",
93180=>"000011111",
93181=>"000110000",
93182=>"110111011",
93183=>"111111010",
93184=>"001000111",
93185=>"111000000",
93186=>"100110111",
93187=>"110110111",
93188=>"101101000",
93189=>"110110110",
93190=>"100110111",
93191=>"010111001",
93192=>"100000100",
93193=>"100100110",
93194=>"010010101",
93195=>"011011001",
93196=>"100000100",
93197=>"111000000",
93198=>"111101100",
93199=>"011001001",
93200=>"000001001",
93201=>"001111011",
93202=>"000100011",
93203=>"011001001",
93204=>"110110110",
93205=>"111110110",
93206=>"100100110",
93207=>"000111011",
93208=>"110000010",
93209=>"011011000",
93210=>"011001001",
93211=>"100110111",
93212=>"000000000",
93213=>"001011001",
93214=>"100110100",
93215=>"011001001",
93216=>"100110111",
93217=>"100110100",
93218=>"001000011",
93219=>"011011000",
93220=>"101111001",
93221=>"011001000",
93222=>"001001001",
93223=>"101011000",
93224=>"001011011",
93225=>"111000001",
93226=>"011000010",
93227=>"000000001",
93228=>"101110001",
93229=>"110001011",
93230=>"111011111",
93231=>"000110011",
93232=>"001100000",
93233=>"000100001",
93234=>"001001011",
93235=>"100100001",
93236=>"011000011",
93237=>"011011010",
93238=>"110001110",
93239=>"111011010",
93240=>"110100111",
93241=>"110110111",
93242=>"100011000",
93243=>"000010000",
93244=>"111111001",
93245=>"010011010",
93246=>"110100100",
93247=>"101100100",
93248=>"000011101",
93249=>"001010001",
93250=>"100100111",
93251=>"101110000",
93252=>"000000010",
93253=>"110110110",
93254=>"001011000",
93255=>"000001000",
93256=>"110111011",
93257=>"010110111",
93258=>"110000011",
93259=>"011100010",
93260=>"010000000",
93261=>"101111111",
93262=>"000111111",
93263=>"011011100",
93264=>"111110110",
93265=>"001111111",
93266=>"110100111",
93267=>"001000000",
93268=>"000000100",
93269=>"000000010",
93270=>"001001001",
93271=>"100100110",
93272=>"000111001",
93273=>"000000000",
93274=>"100000000",
93275=>"001011010",
93276=>"100100011",
93277=>"000000011",
93278=>"001001100",
93279=>"110100111",
93280=>"110110111",
93281=>"001000000",
93282=>"100100111",
93283=>"000100000",
93284=>"110101000",
93285=>"001001010",
93286=>"010001000",
93287=>"011001001",
93288=>"100100101",
93289=>"000011101",
93290=>"001000011",
93291=>"001011000",
93292=>"100101111",
93293=>"011001000",
93294=>"000110011",
93295=>"000010011",
93296=>"110111001",
93297=>"010011000",
93298=>"101001100",
93299=>"001001000",
93300=>"001001000",
93301=>"011011010",
93302=>"100011001",
93303=>"001100110",
93304=>"110110010",
93305=>"000001010",
93306=>"000011111",
93307=>"111110111",
93308=>"101111011",
93309=>"001001001",
93310=>"100100110",
93311=>"110110110",
93312=>"011001010",
93313=>"011000100",
93314=>"011110110",
93315=>"101111001",
93316=>"111100000",
93317=>"111111000",
93318=>"001100000",
93319=>"000001000",
93320=>"100101111",
93321=>"000100110",
93322=>"111110011",
93323=>"011001100",
93324=>"110100110",
93325=>"110100010",
93326=>"110110011",
93327=>"001000001",
93328=>"000001100",
93329=>"110000100",
93330=>"011000000",
93331=>"100000111",
93332=>"000001001",
93333=>"100100100",
93334=>"100100101",
93335=>"011010001",
93336=>"011011000",
93337=>"000000010",
93338=>"111111000",
93339=>"110110110",
93340=>"011010101",
93341=>"110111100",
93342=>"000000100",
93343=>"100110100",
93344=>"011000001",
93345=>"111000010",
93346=>"010000100",
93347=>"110100000",
93348=>"111110000",
93349=>"011011001",
93350=>"000001000",
93351=>"011000010",
93352=>"111110011",
93353=>"110011011",
93354=>"110110110",
93355=>"100100110",
93356=>"111000100",
93357=>"100100100",
93358=>"110110001",
93359=>"010001000",
93360=>"111000100",
93361=>"000010111",
93362=>"111110111",
93363=>"000000000",
93364=>"011001001",
93365=>"001000111",
93366=>"001001001",
93367=>"001111010",
93368=>"000000010",
93369=>"001011011",
93370=>"001011001",
93371=>"111110110",
93372=>"011000000",
93373=>"110111010",
93374=>"110110111",
93375=>"011011000",
93376=>"000000011",
93377=>"110010011",
93378=>"100001100",
93379=>"001001001",
93380=>"001000000",
93381=>"101100100",
93382=>"001001000",
93383=>"100100111",
93384=>"001111011",
93385=>"011111000",
93386=>"011011001",
93387=>"111111111",
93388=>"011000001",
93389=>"110101110",
93390=>"111111110",
93391=>"111001100",
93392=>"111110110",
93393=>"011011000",
93394=>"001001001",
93395=>"100110000",
93396=>"000000100",
93397=>"111100000",
93398=>"110100110",
93399=>"111111111",
93400=>"001011000",
93401=>"011011011",
93402=>"111100110",
93403=>"110100111",
93404=>"110110110",
93405=>"011001111",
93406=>"011011010",
93407=>"101000000",
93408=>"110110111",
93409=>"110110111",
93410=>"111111110",
93411=>"000000001",
93412=>"110100110",
93413=>"101101000",
93414=>"011101100",
93415=>"001100110",
93416=>"001000111",
93417=>"111111000",
93418=>"010110110",
93419=>"100000000",
93420=>"110110110",
93421=>"011011000",
93422=>"000100000",
93423=>"011010000",
93424=>"001001000",
93425=>"001100110",
93426=>"000100110",
93427=>"011011000",
93428=>"110110101",
93429=>"110100110",
93430=>"000001000",
93431=>"000001000",
93432=>"000111011",
93433=>"100101111",
93434=>"011010001",
93435=>"010110001",
93436=>"001000000",
93437=>"101000110",
93438=>"010000001",
93439=>"110110110",
93440=>"011011100",
93441=>"000110111",
93442=>"000000110",
93443=>"000000000",
93444=>"000101000",
93445=>"001100100",
93446=>"010100100",
93447=>"010010010",
93448=>"001001111",
93449=>"000000000",
93450=>"001011110",
93451=>"100111101",
93452=>"111001001",
93453=>"100000011",
93454=>"100000001",
93455=>"000110010",
93456=>"001000001",
93457=>"001000110",
93458=>"101001110",
93459=>"001111000",
93460=>"010110111",
93461=>"101101111",
93462=>"011111011",
93463=>"110001000",
93464=>"100100000",
93465=>"110001001",
93466=>"000000111",
93467=>"100000010",
93468=>"100000000",
93469=>"011010011",
93470=>"101100011",
93471=>"010110101",
93472=>"000000101",
93473=>"100110110",
93474=>"000010010",
93475=>"000111011",
93476=>"001000100",
93477=>"101001000",
93478=>"000001111",
93479=>"100001010",
93480=>"011111111",
93481=>"110101100",
93482=>"000000000",
93483=>"000111000",
93484=>"110000110",
93485=>"111101111",
93486=>"111111101",
93487=>"100000111",
93488=>"111111100",
93489=>"111100100",
93490=>"001000001",
93491=>"101011000",
93492=>"000010000",
93493=>"111010110",
93494=>"100001011",
93495=>"000101111",
93496=>"010101111",
93497=>"000001011",
93498=>"000001001",
93499=>"001000000",
93500=>"000100101",
93501=>"111111010",
93502=>"000000010",
93503=>"111111111",
93504=>"110000000",
93505=>"010000010",
93506=>"010111001",
93507=>"100000001",
93508=>"000010010",
93509=>"110100000",
93510=>"000111111",
93511=>"101111111",
93512=>"010000100",
93513=>"111111111",
93514=>"000001110",
93515=>"111010000",
93516=>"000101101",
93517=>"100000010",
93518=>"110001001",
93519=>"001000010",
93520=>"000111111",
93521=>"101100000",
93522=>"111111010",
93523=>"011001000",
93524=>"000111110",
93525=>"001000000",
93526=>"000101001",
93527=>"000000010",
93528=>"001001111",
93529=>"011001011",
93530=>"000000100",
93531=>"010100111",
93532=>"000000100",
93533=>"000011010",
93534=>"010101011",
93535=>"100100101",
93536=>"000000000",
93537=>"010111111",
93538=>"101000010",
93539=>"011001011",
93540=>"110000000",
93541=>"001011000",
93542=>"101111100",
93543=>"000010000",
93544=>"010001000",
93545=>"111001000",
93546=>"101111101",
93547=>"110000000",
93548=>"111011000",
93549=>"111000111",
93550=>"000000000",
93551=>"011111111",
93552=>"000101111",
93553=>"100101110",
93554=>"000111110",
93555=>"111000000",
93556=>"110001111",
93557=>"100000000",
93558=>"111111000",
93559=>"000000000",
93560=>"000001000",
93561=>"000000000",
93562=>"111000000",
93563=>"111001101",
93564=>"101100000",
93565=>"111000000",
93566=>"010010111",
93567=>"111001111",
93568=>"100010010",
93569=>"110110111",
93570=>"101111011",
93571=>"110111111",
93572=>"010001011",
93573=>"010111000",
93574=>"111011010",
93575=>"100000000",
93576=>"100001011",
93577=>"010000000",
93578=>"101101001",
93579=>"000100111",
93580=>"000100100",
93581=>"111101010",
93582=>"000101111",
93583=>"001100100",
93584=>"111111001",
93585=>"000010111",
93586=>"010001111",
93587=>"100100011",
93588=>"000100010",
93589=>"001000000",
93590=>"111110010",
93591=>"111000001",
93592=>"111111000",
93593=>"011011000",
93594=>"000111111",
93595=>"000000100",
93596=>"000111000",
93597=>"001000000",
93598=>"010100110",
93599=>"101101110",
93600=>"001100111",
93601=>"000010111",
93602=>"000000111",
93603=>"000110111",
93604=>"101110010",
93605=>"001111111",
93606=>"111000110",
93607=>"000110111",
93608=>"101000010",
93609=>"110110000",
93610=>"101100110",
93611=>"100011110",
93612=>"100000000",
93613=>"000101111",
93614=>"001011110",
93615=>"001011111",
93616=>"000111111",
93617=>"001000101",
93618=>"001010000",
93619=>"011011111",
93620=>"011111101",
93621=>"000111000",
93622=>"100000011",
93623=>"110000011",
93624=>"010001101",
93625=>"001101010",
93626=>"001101000",
93627=>"000000000",
93628=>"111000111",
93629=>"111000110",
93630=>"100001101",
93631=>"000111111",
93632=>"000111011",
93633=>"100000000",
93634=>"000101110",
93635=>"000010111",
93636=>"000000000",
93637=>"001111100",
93638=>"111010010",
93639=>"000000110",
93640=>"111100101",
93641=>"000000111",
93642=>"000000001",
93643=>"011010011",
93644=>"000101010",
93645=>"101000100",
93646=>"000010011",
93647=>"111001000",
93648=>"000000111",
93649=>"110001101",
93650=>"010100000",
93651=>"001101110",
93652=>"111000000",
93653=>"000000000",
93654=>"000101000",
93655=>"000101000",
93656=>"010011001",
93657=>"001110111",
93658=>"111011110",
93659=>"101000000",
93660=>"111111111",
93661=>"100000101",
93662=>"110111110",
93663=>"101110000",
93664=>"011000100",
93665=>"001011111",
93666=>"000000001",
93667=>"001000111",
93668=>"000110000",
93669=>"111100100",
93670=>"101101111",
93671=>"000101101",
93672=>"111101111",
93673=>"111001010",
93674=>"100100011",
93675=>"101011010",
93676=>"000000000",
93677=>"001001101",
93678=>"001000100",
93679=>"001011000",
93680=>"100000000",
93681=>"100101011",
93682=>"001101100",
93683=>"100110110",
93684=>"111110001",
93685=>"101101111",
93686=>"001001000",
93687=>"000010000",
93688=>"000000000",
93689=>"110011011",
93690=>"111111111",
93691=>"111000000",
93692=>"101111000",
93693=>"001010011",
93694=>"101011010",
93695=>"001001000",
93696=>"000000000",
93697=>"000100101",
93698=>"000111111",
93699=>"111111111",
93700=>"001110111",
93701=>"111001000",
93702=>"001000000",
93703=>"011010000",
93704=>"011111110",
93705=>"010110101",
93706=>"011001001",
93707=>"000000001",
93708=>"101000111",
93709=>"000011000",
93710=>"110110011",
93711=>"101111111",
93712=>"111101000",
93713=>"111111111",
93714=>"110111010",
93715=>"001000001",
93716=>"000010100",
93717=>"010000010",
93718=>"100000100",
93719=>"000000000",
93720=>"000000000",
93721=>"000001101",
93722=>"111011000",
93723=>"000010011",
93724=>"000101101",
93725=>"000000000",
93726=>"111000000",
93727=>"011000001",
93728=>"010110100",
93729=>"010000000",
93730=>"010000100",
93731=>"000000110",
93732=>"011111110",
93733=>"000000000",
93734=>"111000000",
93735=>"110111111",
93736=>"111110000",
93737=>"101101101",
93738=>"101101111",
93739=>"111111111",
93740=>"001001001",
93741=>"010000000",
93742=>"111000001",
93743=>"000000000",
93744=>"000000000",
93745=>"111111111",
93746=>"111011100",
93747=>"000011011",
93748=>"001000100",
93749=>"111111111",
93750=>"111001000",
93751=>"000000110",
93752=>"111100000",
93753=>"000000100",
93754=>"000101101",
93755=>"000010111",
93756=>"001011111",
93757=>"000001001",
93758=>"011111101",
93759=>"111111011",
93760=>"111000000",
93761=>"100000000",
93762=>"111111001",
93763=>"111111111",
93764=>"000010000",
93765=>"000000111",
93766=>"111010010",
93767=>"011011111",
93768=>"000000000",
93769=>"111111010",
93770=>"000011101",
93771=>"010111000",
93772=>"000001111",
93773=>"111111111",
93774=>"111111010",
93775=>"000000000",
93776=>"111111001",
93777=>"110111111",
93778=>"111111110",
93779=>"001000000",
93780=>"111111111",
93781=>"000001011",
93782=>"000001000",
93783=>"101101111",
93784=>"011001101",
93785=>"101111001",
93786=>"000000100",
93787=>"000010011",
93788=>"111111000",
93789=>"001001001",
93790=>"000111111",
93791=>"111111111",
93792=>"110010000",
93793=>"111100000",
93794=>"000010000",
93795=>"000000000",
93796=>"000110100",
93797=>"000000001",
93798=>"110000000",
93799=>"000111111",
93800=>"111111100",
93801=>"000000001",
93802=>"111001000",
93803=>"000111001",
93804=>"101011000",
93805=>"000000000",
93806=>"011000000",
93807=>"000000000",
93808=>"110110100",
93809=>"000000101",
93810=>"011000110",
93811=>"111111111",
93812=>"101110110",
93813=>"000000000",
93814=>"111111111",
93815=>"101111111",
93816=>"000000001",
93817=>"000000101",
93818=>"000000111",
93819=>"101111000",
93820=>"100110110",
93821=>"100001001",
93822=>"111111110",
93823=>"111111110",
93824=>"000101010",
93825=>"111000000",
93826=>"111111111",
93827=>"101001101",
93828=>"110000110",
93829=>"001011000",
93830=>"001011001",
93831=>"100001011",
93832=>"011011011",
93833=>"111110100",
93834=>"011011000",
93835=>"001111111",
93836=>"111111001",
93837=>"011010010",
93838=>"000000000",
93839=>"111111100",
93840=>"011111111",
93841=>"110101000",
93842=>"111111111",
93843=>"000000000",
93844=>"000011111",
93845=>"101100111",
93846=>"111001000",
93847=>"110000000",
93848=>"100000000",
93849=>"000001111",
93850=>"010111111",
93851=>"000010000",
93852=>"010011001",
93853=>"000100000",
93854=>"111000000",
93855=>"000000000",
93856=>"000100000",
93857=>"000111111",
93858=>"111111111",
93859=>"010100001",
93860=>"010101101",
93861=>"001000000",
93862=>"001001111",
93863=>"001001000",
93864=>"111000001",
93865=>"001000010",
93866=>"000010000",
93867=>"111110101",
93868=>"101000101",
93869=>"111110111",
93870=>"011001000",
93871=>"011111101",
93872=>"111110000",
93873=>"011001000",
93874=>"001000000",
93875=>"000010110",
93876=>"100000111",
93877=>"100011111",
93878=>"100100000",
93879=>"100000111",
93880=>"000100011",
93881=>"001100111",
93882=>"111101000",
93883=>"001111111",
93884=>"000110111",
93885=>"111111111",
93886=>"111111110",
93887=>"010101000",
93888=>"001001111",
93889=>"011010000",
93890=>"100100111",
93891=>"000110110",
93892=>"000000000",
93893=>"000000001",
93894=>"110111000",
93895=>"010111011",
93896=>"001001110",
93897=>"000000000",
93898=>"001111010",
93899=>"000000111",
93900=>"111111011",
93901=>"000011011",
93902=>"000000000",
93903=>"011110010",
93904=>"000011111",
93905=>"011011001",
93906=>"111000000",
93907=>"011011111",
93908=>"111110010",
93909=>"111100001",
93910=>"101000000",
93911=>"001000111",
93912=>"010111111",
93913=>"000111111",
93914=>"000000000",
93915=>"000011011",
93916=>"011000110",
93917=>"000011111",
93918=>"010001111",
93919=>"011110110",
93920=>"111111000",
93921=>"011000001",
93922=>"110110110",
93923=>"111110110",
93924=>"111000000",
93925=>"101101111",
93926=>"000000001",
93927=>"011101000",
93928=>"111111011",
93929=>"110100111",
93930=>"110100000",
93931=>"000001111",
93932=>"111001000",
93933=>"001001111",
93934=>"010000000",
93935=>"000010010",
93936=>"000000100",
93937=>"000000001",
93938=>"000000101",
93939=>"001011100",
93940=>"110001000",
93941=>"111111111",
93942=>"111111011",
93943=>"000000011",
93944=>"000000001",
93945=>"000000000",
93946=>"000001100",
93947=>"000000010",
93948=>"011111010",
93949=>"101111011",
93950=>"100100000",
93951=>"000000100",
93952=>"101111011",
93953=>"000000000",
93954=>"010110110",
93955=>"111000000",
93956=>"001111111",
93957=>"000000110",
93958=>"000000001",
93959=>"011110111",
93960=>"000000000",
93961=>"001000111",
93962=>"011000100",
93963=>"111111111",
93964=>"010010000",
93965=>"111111001",
93966=>"111101111",
93967=>"000111110",
93968=>"111011000",
93969=>"101000110",
93970=>"000000110",
93971=>"000000001",
93972=>"111101111",
93973=>"000010010",
93974=>"000000111",
93975=>"111110110",
93976=>"000000111",
93977=>"000010000",
93978=>"101111111",
93979=>"110111111",
93980=>"100111011",
93981=>"101101000",
93982=>"101111011",
93983=>"000000000",
93984=>"101000111",
93985=>"111111011",
93986=>"110000000",
93987=>"000000000",
93988=>"111100101",
93989=>"111011111",
93990=>"110010010",
93991=>"110111111",
93992=>"101010010",
93993=>"100010111",
93994=>"111111111",
93995=>"000000000",
93996=>"100101111",
93997=>"000000000",
93998=>"110010111",
93999=>"011111111",
94000=>"111100110",
94001=>"101001001",
94002=>"000111000",
94003=>"101000000",
94004=>"101101101",
94005=>"000111101",
94006=>"000001001",
94007=>"111001001",
94008=>"111000010",
94009=>"000110111",
94010=>"101000000",
94011=>"000000000",
94012=>"111011001",
94013=>"111111111",
94014=>"000000100",
94015=>"100110101",
94016=>"000011111",
94017=>"101101111",
94018=>"100001010",
94019=>"011111111",
94020=>"000001000",
94021=>"000001000",
94022=>"110011101",
94023=>"001000000",
94024=>"111001111",
94025=>"111111000",
94026=>"111001001",
94027=>"000000000",
94028=>"101100100",
94029=>"001111111",
94030=>"111101001",
94031=>"111010101",
94032=>"100111111",
94033=>"111111111",
94034=>"000000001",
94035=>"100000101",
94036=>"000000110",
94037=>"000011111",
94038=>"000000010",
94039=>"110111101",
94040=>"001110000",
94041=>"001010000",
94042=>"111111111",
94043=>"001001001",
94044=>"111001000",
94045=>"100100100",
94046=>"101000000",
94047=>"110000011",
94048=>"000000011",
94049=>"001011001",
94050=>"000001101",
94051=>"011010011",
94052=>"011111111",
94053=>"000011101",
94054=>"110011101",
94055=>"111110110",
94056=>"001000000",
94057=>"111101110",
94058=>"111000110",
94059=>"111111111",
94060=>"111110000",
94061=>"111011010",
94062=>"011001000",
94063=>"001111000",
94064=>"001001001",
94065=>"111111111",
94066=>"011110100",
94067=>"000000000",
94068=>"111000000",
94069=>"000000000",
94070=>"010110000",
94071=>"000101111",
94072=>"000010111",
94073=>"000000000",
94074=>"000000000",
94075=>"111010000",
94076=>"101101101",
94077=>"111000101",
94078=>"111011000",
94079=>"101101000",
94080=>"010000000",
94081=>"000000000",
94082=>"111101111",
94083=>"100000010",
94084=>"111000000",
94085=>"000010111",
94086=>"100101111",
94087=>"100000000",
94088=>"110011001",
94089=>"001000000",
94090=>"111000101",
94091=>"111111010",
94092=>"101000100",
94093=>"100001110",
94094=>"000100111",
94095=>"011010000",
94096=>"100100100",
94097=>"010111111",
94098=>"110010000",
94099=>"111111000",
94100=>"110100101",
94101=>"001000111",
94102=>"011111111",
94103=>"000100100",
94104=>"010111111",
94105=>"010000101",
94106=>"010110110",
94107=>"000001111",
94108=>"001011111",
94109=>"001101111",
94110=>"111110001",
94111=>"011111110",
94112=>"110110110",
94113=>"000111111",
94114=>"111111000",
94115=>"110100111",
94116=>"000000111",
94117=>"000001100",
94118=>"001110110",
94119=>"000111111",
94120=>"001000000",
94121=>"000000000",
94122=>"110111111",
94123=>"011010010",
94124=>"000000000",
94125=>"111000000",
94126=>"111011000",
94127=>"111000000",
94128=>"011011000",
94129=>"101011100",
94130=>"101101100",
94131=>"101001101",
94132=>"001110110",
94133=>"101001000",
94134=>"000000001",
94135=>"111010001",
94136=>"010110000",
94137=>"001001100",
94138=>"010111101",
94139=>"000010000",
94140=>"101100010",
94141=>"111101101",
94142=>"000100000",
94143=>"100101110",
94144=>"111000000",
94145=>"110101111",
94146=>"111111111",
94147=>"101110001",
94148=>"100111110",
94149=>"111100001",
94150=>"111110000",
94151=>"101101101",
94152=>"101000001",
94153=>"000000000",
94154=>"110010011",
94155=>"000000000",
94156=>"000010111",
94157=>"101000001",
94158=>"000000100",
94159=>"000000000",
94160=>"010110111",
94161=>"100111110",
94162=>"000000000",
94163=>"011001000",
94164=>"101111111",
94165=>"000000110",
94166=>"111111111",
94167=>"111000001",
94168=>"111100001",
94169=>"000000001",
94170=>"000000011",
94171=>"111000000",
94172=>"011011111",
94173=>"011010010",
94174=>"000010000",
94175=>"111010000",
94176=>"000111011",
94177=>"100111001",
94178=>"111110100",
94179=>"111111000",
94180=>"101000010",
94181=>"111101000",
94182=>"100111111",
94183=>"100101000",
94184=>"000000111",
94185=>"000000000",
94186=>"111100100",
94187=>"001001000",
94188=>"000111010",
94189=>"001111000",
94190=>"000110100",
94191=>"111000100",
94192=>"111101000",
94193=>"111001110",
94194=>"111000000",
94195=>"101111111",
94196=>"101101100",
94197=>"101000000",
94198=>"000000000",
94199=>"111101111",
94200=>"000111111",
94201=>"111000000",
94202=>"101101101",
94203=>"101111111",
94204=>"010111111",
94205=>"101000000",
94206=>"000000110",
94207=>"111110111",
94208=>"011011000",
94209=>"000111110",
94210=>"101000110",
94211=>"000000100",
94212=>"110110000",
94213=>"100110000",
94214=>"111101110",
94215=>"000000100",
94216=>"110010000",
94217=>"001000101",
94218=>"001110111",
94219=>"010110111",
94220=>"000000001",
94221=>"000000001",
94222=>"100001010",
94223=>"111111111",
94224=>"110110010",
94225=>"100111111",
94226=>"000000010",
94227=>"100101000",
94228=>"111111111",
94229=>"111110000",
94230=>"100100110",
94231=>"000011110",
94232=>"110101111",
94233=>"111111010",
94234=>"000000001",
94235=>"100111111",
94236=>"000001111",
94237=>"011101111",
94238=>"111000000",
94239=>"000101100",
94240=>"000000010",
94241=>"000000101",
94242=>"111111101",
94243=>"101000000",
94244=>"000100100",
94245=>"010001011",
94246=>"000010111",
94247=>"111000000",
94248=>"010010110",
94249=>"110110110",
94250=>"111000011",
94251=>"110110110",
94252=>"011011111",
94253=>"101000000",
94254=>"011110000",
94255=>"010001000",
94256=>"010000000",
94257=>"000101001",
94258=>"010000000",
94259=>"111111011",
94260=>"001000100",
94261=>"010111111",
94262=>"111011011",
94263=>"011011001",
94264=>"111111110",
94265=>"011000110",
94266=>"100110000",
94267=>"111111000",
94268=>"011011001",
94269=>"101101111",
94270=>"000001101",
94271=>"111111111",
94272=>"000110111",
94273=>"101001010",
94274=>"000100000",
94275=>"011011000",
94276=>"000001111",
94277=>"000000000",
94278=>"000000000",
94279=>"000011101",
94280=>"001101111",
94281=>"011110010",
94282=>"000000000",
94283=>"111111000",
94284=>"111101101",
94285=>"011011000",
94286=>"000100100",
94287=>"111111111",
94288=>"101101101",
94289=>"101111111",
94290=>"000000111",
94291=>"001101010",
94292=>"010110010",
94293=>"101111111",
94294=>"000011001",
94295=>"001000111",
94296=>"010101111",
94297=>"001101011",
94298=>"101111111",
94299=>"110110111",
94300=>"001000101",
94301=>"001001111",
94302=>"111111000",
94303=>"010010000",
94304=>"111111111",
94305=>"001111000",
94306=>"111011000",
94307=>"111111100",
94308=>"110111111",
94309=>"000100100",
94310=>"010000000",
94311=>"110001000",
94312=>"111111110",
94313=>"000000011",
94314=>"111010110",
94315=>"110011111",
94316=>"111111111",
94317=>"111111010",
94318=>"001000100",
94319=>"011101111",
94320=>"011001000",
94321=>"000000111",
94322=>"111100110",
94323=>"111010110",
94324=>"100101010",
94325=>"100000000",
94326=>"111101110",
94327=>"110010001",
94328=>"010111111",
94329=>"110000000",
94330=>"010110111",
94331=>"100000000",
94332=>"111101111",
94333=>"110100000",
94334=>"011010000",
94335=>"101101000",
94336=>"010010010",
94337=>"000001000",
94338=>"111011011",
94339=>"000011011",
94340=>"001001000",
94341=>"011110101",
94342=>"101100100",
94343=>"010110010",
94344=>"000111001",
94345=>"111111111",
94346=>"111001000",
94347=>"010011000",
94348=>"100111011",
94349=>"110000000",
94350=>"000111001",
94351=>"101001011",
94352=>"110101000",
94353=>"000010111",
94354=>"001000111",
94355=>"000000111",
94356=>"000111111",
94357=>"000000001",
94358=>"111011010",
94359=>"001011011",
94360=>"111111111",
94361=>"111111111",
94362=>"101000000",
94363=>"110100000",
94364=>"111001000",
94365=>"111111010",
94366=>"000010100",
94367=>"010000001",
94368=>"001001111",
94369=>"111111111",
94370=>"000000111",
94371=>"111011111",
94372=>"111111000",
94373=>"010111110",
94374=>"011101111",
94375=>"000000001",
94376=>"111000010",
94377=>"000110111",
94378=>"000000000",
94379=>"000101110",
94380=>"111111101",
94381=>"101000000",
94382=>"111001011",
94383=>"010010000",
94384=>"000001101",
94385=>"011101111",
94386=>"001000111",
94387=>"000101110",
94388=>"100111111",
94389=>"000111110",
94390=>"010110100",
94391=>"000000000",
94392=>"111110001",
94393=>"000110111",
94394=>"110000111",
94395=>"000111111",
94396=>"010111100",
94397=>"100111111",
94398=>"111010000",
94399=>"010000100",
94400=>"110000110",
94401=>"000000011",
94402=>"000110111",
94403=>"100101010",
94404=>"110111001",
94405=>"110100101",
94406=>"000000111",
94407=>"001000001",
94408=>"110000000",
94409=>"000111001",
94410=>"000000001",
94411=>"110111110",
94412=>"111111010",
94413=>"010111110",
94414=>"111110010",
94415=>"000000000",
94416=>"111110000",
94417=>"111110011",
94418=>"111100110",
94419=>"000000101",
94420=>"101000000",
94421=>"100100110",
94422=>"000000000",
94423=>"000001111",
94424=>"000000111",
94425=>"000000000",
94426=>"000000101",
94427=>"101100000",
94428=>"011011101",
94429=>"010110010",
94430=>"110110010",
94431=>"011000000",
94432=>"001101101",
94433=>"001000000",
94434=>"000000100",
94435=>"101010000",
94436=>"000000000",
94437=>"000111101",
94438=>"010011000",
94439=>"010011000",
94440=>"000000010",
94441=>"000000001",
94442=>"100111110",
94443=>"000110111",
94444=>"000000111",
94445=>"000100101",
94446=>"000000000",
94447=>"001111000",
94448=>"000010010",
94449=>"011100111",
94450=>"111110011",
94451=>"111111111",
94452=>"100100100",
94453=>"111111101",
94454=>"000011011",
94455=>"111111111",
94456=>"010011111",
94457=>"101000110",
94458=>"111111111",
94459=>"000001001",
94460=>"000000000",
94461=>"000111110",
94462=>"100010000",
94463=>"000000101",
94464=>"111001001",
94465=>"110111000",
94466=>"001110000",
94467=>"001001000",
94468=>"000011010",
94469=>"011111000",
94470=>"111100110",
94471=>"100000011",
94472=>"011010000",
94473=>"000000001",
94474=>"111000000",
94475=>"000000000",
94476=>"001011000",
94477=>"001111010",
94478=>"101100001",
94479=>"001100000",
94480=>"111111011",
94481=>"000000111",
94482=>"110110100",
94483=>"000100010",
94484=>"100011111",
94485=>"010111010",
94486=>"110110111",
94487=>"111101111",
94488=>"101100101",
94489=>"101100100",
94490=>"011111011",
94491=>"111111100",
94492=>"101110110",
94493=>"100100110",
94494=>"111111101",
94495=>"000110011",
94496=>"000000000",
94497=>"011011000",
94498=>"101001000",
94499=>"110000100",
94500=>"011011011",
94501=>"011001000",
94502=>"010111010",
94503=>"111101000",
94504=>"010000000",
94505=>"110111100",
94506=>"000010000",
94507=>"000000000",
94508=>"111111011",
94509=>"101001011",
94510=>"101011001",
94511=>"000000000",
94512=>"000000111",
94513=>"100100000",
94514=>"111010001",
94515=>"010111111",
94516=>"011111111",
94517=>"000000000",
94518=>"100011011",
94519=>"001000001",
94520=>"001011110",
94521=>"000111010",
94522=>"000010000",
94523=>"010011011",
94524=>"011101100",
94525=>"110111111",
94526=>"000000001",
94527=>"100000110",
94528=>"011101111",
94529=>"111111111",
94530=>"010010000",
94531=>"001000010",
94532=>"111111111",
94533=>"000000100",
94534=>"111111010",
94535=>"000111011",
94536=>"000100000",
94537=>"000000000",
94538=>"000000001",
94539=>"111000000",
94540=>"111111111",
94541=>"101111111",
94542=>"011111101",
94543=>"111011000",
94544=>"001111111",
94545=>"110111111",
94546=>"111111111",
94547=>"111111111",
94548=>"111111101",
94549=>"101110111",
94550=>"111011101",
94551=>"001000000",
94552=>"000000000",
94553=>"011110110",
94554=>"100100101",
94555=>"010110010",
94556=>"000000100",
94557=>"111001001",
94558=>"111111111",
94559=>"101000011",
94560=>"111111111",
94561=>"111000000",
94562=>"010010010",
94563=>"111011101",
94564=>"111111111",
94565=>"111100001",
94566=>"000001000",
94567=>"110100111",
94568=>"000000000",
94569=>"111011000",
94570=>"010010110",
94571=>"111111000",
94572=>"111111111",
94573=>"100001000",
94574=>"011001000",
94575=>"111111111",
94576=>"101001001",
94577=>"100011000",
94578=>"000100110",
94579=>"100000111",
94580=>"000000011",
94581=>"000000001",
94582=>"000111100",
94583=>"001100001",
94584=>"010000000",
94585=>"111111000",
94586=>"011000111",
94587=>"000000110",
94588=>"011101111",
94589=>"001000000",
94590=>"000001111",
94591=>"101000111",
94592=>"111111101",
94593=>"000000000",
94594=>"111101000",
94595=>"111110000",
94596=>"111111011",
94597=>"011011111",
94598=>"110111000",
94599=>"111100110",
94600=>"100100100",
94601=>"111011111",
94602=>"100111100",
94603=>"001000000",
94604=>"000000011",
94605=>"000000100",
94606=>"100000110",
94607=>"011000001",
94608=>"000011110",
94609=>"000010010",
94610=>"111000011",
94611=>"001000011",
94612=>"111101001",
94613=>"000111011",
94614=>"011111011",
94615=>"000011011",
94616=>"000000000",
94617=>"111111000",
94618=>"000101001",
94619=>"101000000",
94620=>"000111111",
94621=>"111001011",
94622=>"000001111",
94623=>"010010000",
94624=>"000000000",
94625=>"000111101",
94626=>"110000101",
94627=>"111111000",
94628=>"011110101",
94629=>"010011011",
94630=>"100000100",
94631=>"111111101",
94632=>"111011011",
94633=>"000111010",
94634=>"000000000",
94635=>"000000000",
94636=>"100100110",
94637=>"011111111",
94638=>"101001001",
94639=>"111111110",
94640=>"000010000",
94641=>"000000000",
94642=>"110110100",
94643=>"111011011",
94644=>"100101000",
94645=>"000000000",
94646=>"011000000",
94647=>"100000000",
94648=>"100110101",
94649=>"111000001",
94650=>"001111011",
94651=>"111000000",
94652=>"100000001",
94653=>"010010010",
94654=>"111001001",
94655=>"000000000",
94656=>"101100100",
94657=>"101000011",
94658=>"111000011",
94659=>"110110111",
94660=>"011001001",
94661=>"111100000",
94662=>"011011000",
94663=>"100100000",
94664=>"110000100",
94665=>"000011011",
94666=>"010100000",
94667=>"111011000",
94668=>"101100000",
94669=>"111111111",
94670=>"000101111",
94671=>"000000000",
94672=>"111100111",
94673=>"010110110",
94674=>"000010101",
94675=>"010010000",
94676=>"101001111",
94677=>"100100110",
94678=>"010111111",
94679=>"101011111",
94680=>"000000000",
94681=>"010000010",
94682=>"100000000",
94683=>"000000000",
94684=>"111111110",
94685=>"100000000",
94686=>"000001001",
94687=>"001111101",
94688=>"100000100",
94689=>"000100101",
94690=>"000000101",
94691=>"110101001",
94692=>"111101000",
94693=>"100100110",
94694=>"001000000",
94695=>"101101100",
94696=>"110111101",
94697=>"111100111",
94698=>"110000000",
94699=>"000000010",
94700=>"000000001",
94701=>"000101101",
94702=>"111010110",
94703=>"001000101",
94704=>"000000000",
94705=>"101001011",
94706=>"111111000",
94707=>"011011011",
94708=>"111101101",
94709=>"000000011",
94710=>"111011010",
94711=>"111111101",
94712=>"011001000",
94713=>"000001011",
94714=>"000010000",
94715=>"101101101",
94716=>"000111111",
94717=>"111001111",
94718=>"110110010",
94719=>"110000000",
94720=>"011101100",
94721=>"100000011",
94722=>"000101111",
94723=>"000000110",
94724=>"011011111",
94725=>"110111011",
94726=>"111011010",
94727=>"110011111",
94728=>"010000101",
94729=>"111000001",
94730=>"011000000",
94731=>"011001111",
94732=>"110001111",
94733=>"011001000",
94734=>"011000010",
94735=>"110000110",
94736=>"111101000",
94737=>"101100000",
94738=>"000000000",
94739=>"111111000",
94740=>"010110111",
94741=>"001111110",
94742=>"000110110",
94743=>"111110100",
94744=>"000110000",
94745=>"111110010",
94746=>"000111111",
94747=>"001101011",
94748=>"110011010",
94749=>"000001100",
94750=>"000011011",
94751=>"010000000",
94752=>"000000000",
94753=>"000001110",
94754=>"010000000",
94755=>"110011000",
94756=>"100001000",
94757=>"100101110",
94758=>"000010110",
94759=>"110110000",
94760=>"111111111",
94761=>"001001011",
94762=>"010000000",
94763=>"000111000",
94764=>"010100011",
94765=>"110111111",
94766=>"111110111",
94767=>"100000111",
94768=>"000000000",
94769=>"111111111",
94770=>"000001001",
94771=>"111111000",
94772=>"001000000",
94773=>"111010110",
94774=>"100000101",
94775=>"111111000",
94776=>"100111111",
94777=>"110010000",
94778=>"111000000",
94779=>"111011011",
94780=>"110010110",
94781=>"111010010",
94782=>"001000000",
94783=>"001110110",
94784=>"111000011",
94785=>"100100110",
94786=>"000001000",
94787=>"001100111",
94788=>"010000000",
94789=>"011010000",
94790=>"110010000",
94791=>"010010101",
94792=>"010011110",
94793=>"010000010",
94794=>"101000000",
94795=>"111100000",
94796=>"000000001",
94797=>"001111111",
94798=>"111111110",
94799=>"000001100",
94800=>"001000111",
94801=>"101001000",
94802=>"011101000",
94803=>"001100000",
94804=>"010010001",
94805=>"100001011",
94806=>"100100100",
94807=>"110001011",
94808=>"101100111",
94809=>"011011011",
94810=>"001001110",
94811=>"110100100",
94812=>"000001111",
94813=>"001001001",
94814=>"000111111",
94815=>"100001111",
94816=>"000000111",
94817=>"000000100",
94818=>"000000111",
94819=>"100110110",
94820=>"111110100",
94821=>"000011001",
94822=>"001111110",
94823=>"010010000",
94824=>"011110011",
94825=>"010010010",
94826=>"100100111",
94827=>"110000001",
94828=>"000100111",
94829=>"111111000",
94830=>"001001000",
94831=>"010010000",
94832=>"011001011",
94833=>"111001000",
94834=>"111101001",
94835=>"110011000",
94836=>"000010010",
94837=>"101001000",
94838=>"110000100",
94839=>"000000001",
94840=>"000010110",
94841=>"111010000",
94842=>"111001001",
94843=>"001111101",
94844=>"110011011",
94845=>"100000000",
94846=>"101111111",
94847=>"111000101",
94848=>"000000000",
94849=>"101100111",
94850=>"010011111",
94851=>"000111111",
94852=>"011111111",
94853=>"000000100",
94854=>"101111010",
94855=>"000000000",
94856=>"111101100",
94857=>"000000000",
94858=>"111000000",
94859=>"000000110",
94860=>"111111111",
94861=>"000000000",
94862=>"001111000",
94863=>"001000000",
94864=>"011100110",
94865=>"111000110",
94866=>"111011011",
94867=>"010111101",
94868=>"101010100",
94869=>"101000000",
94870=>"111000111",
94871=>"100000001",
94872=>"011001000",
94873=>"000010111",
94874=>"001000111",
94875=>"001001111",
94876=>"010011011",
94877=>"001101101",
94878=>"010000010",
94879=>"111010000",
94880=>"110100111",
94881=>"101101000",
94882=>"101000000",
94883=>"101101110",
94884=>"001111000",
94885=>"110010000",
94886=>"110111010",
94887=>"000001001",
94888=>"111111111",
94889=>"000000110",
94890=>"001111111",
94891=>"001000000",
94892=>"000001000",
94893=>"000110000",
94894=>"101011011",
94895=>"111000000",
94896=>"001000101",
94897=>"111111011",
94898=>"000100000",
94899=>"000000010",
94900=>"110111011",
94901=>"111011010",
94902=>"111000000",
94903=>"110111000",
94904=>"011000001",
94905=>"010110000",
94906=>"000000111",
94907=>"111000010",
94908=>"101000010",
94909=>"101000111",
94910=>"000001111",
94911=>"000011000",
94912=>"010000000",
94913=>"111010000",
94914=>"000101010",
94915=>"011000100",
94916=>"000010000",
94917=>"100001111",
94918=>"011111011",
94919=>"111000001",
94920=>"111010011",
94921=>"111101100",
94922=>"100000000",
94923=>"000100111",
94924=>"011000010",
94925=>"011110110",
94926=>"111010000",
94927=>"110001111",
94928=>"010000000",
94929=>"011001011",
94930=>"011010010",
94931=>"011010000",
94932=>"010000111",
94933=>"101100110",
94934=>"001000111",
94935=>"000000000",
94936=>"110010000",
94937=>"001111001",
94938=>"001001000",
94939=>"101100001",
94940=>"000110110",
94941=>"000010111",
94942=>"111010000",
94943=>"101110101",
94944=>"000001101",
94945=>"100111110",
94946=>"000111111",
94947=>"100101010",
94948=>"110100000",
94949=>"011000000",
94950=>"010010000",
94951=>"101101001",
94952=>"000000000",
94953=>"010010101",
94954=>"000000001",
94955=>"101000000",
94956=>"000001111",
94957=>"000110000",
94958=>"011000001",
94959=>"111111000",
94960=>"111000000",
94961=>"000001111",
94962=>"010111111",
94963=>"111000000",
94964=>"110001011",
94965=>"011011111",
94966=>"111000000",
94967=>"110101111",
94968=>"000000000",
94969=>"000010000",
94970=>"001101000",
94971=>"011111110",
94972=>"011000000",
94973=>"001101111",
94974=>"110111101",
94975=>"100001000",
94976=>"100011010",
94977=>"000010110",
94978=>"011001001",
94979=>"111111001",
94980=>"101000011",
94981=>"000001110",
94982=>"111001011",
94983=>"000110110",
94984=>"000001110",
94985=>"011001011",
94986=>"100001000",
94987=>"000000100",
94988=>"000000100",
94989=>"000000000",
94990=>"100000111",
94991=>"011001000",
94992=>"000110110",
94993=>"011001001",
94994=>"110011000",
94995=>"011000000",
94996=>"001111100",
94997=>"111101100",
94998=>"011011010",
94999=>"111001110",
95000=>"010001001",
95001=>"011111100",
95002=>"100001001",
95003=>"100100100",
95004=>"011111001",
95005=>"010000001",
95006=>"100110110",
95007=>"100100000",
95008=>"100001000",
95009=>"001100110",
95010=>"111011001",
95011=>"001110100",
95012=>"100010101",
95013=>"010111001",
95014=>"000000000",
95015=>"100110000",
95016=>"011001111",
95017=>"010110110",
95018=>"011000010",
95019=>"111001001",
95020=>"100100101",
95021=>"100110101",
95022=>"110111000",
95023=>"011001000",
95024=>"111011010",
95025=>"000011011",
95026=>"011100000",
95027=>"110100001",
95028=>"011011001",
95029=>"111111101",
95030=>"000000000",
95031=>"100110100",
95032=>"100100000",
95033=>"000000110",
95034=>"000001000",
95035=>"001011111",
95036=>"011011111",
95037=>"000110001",
95038=>"000001001",
95039=>"101110110",
95040=>"011001100",
95041=>"000100110",
95042=>"010000100",
95043=>"010110110",
95044=>"000011000",
95045=>"000000011",
95046=>"111001001",
95047=>"011110100",
95048=>"111111110",
95049=>"100010000",
95050=>"000110110",
95051=>"111000111",
95052=>"110110100",
95053=>"000000000",
95054=>"000000000",
95055=>"111111101",
95056=>"110010011",
95057=>"100111111",
95058=>"001001100",
95059=>"010011000",
95060=>"000011001",
95061=>"111001111",
95062=>"010011100",
95063=>"000001011",
95064=>"111011100",
95065=>"001001110",
95066=>"110000000",
95067=>"100110110",
95068=>"100100000",
95069=>"100010000",
95070=>"111100001",
95071=>"110111111",
95072=>"000000000",
95073=>"110001011",
95074=>"111001001",
95075=>"101111011",
95076=>"000100110",
95077=>"001001000",
95078=>"100110000",
95079=>"111001001",
95080=>"100011000",
95081=>"110001000",
95082=>"001001100",
95083=>"110110000",
95084=>"110110000",
95085=>"011001011",
95086=>"110001001",
95087=>"000000100",
95088=>"100111111",
95089=>"100000100",
95090=>"000000110",
95091=>"000000011",
95092=>"110110000",
95093=>"010001000",
95094=>"010000100",
95095=>"001001000",
95096=>"111001001",
95097=>"110111110",
95098=>"111001001",
95099=>"000001111",
95100=>"011001100",
95101=>"100000100",
95102=>"101111011",
95103=>"100110001",
95104=>"110111001",
95105=>"000110110",
95106=>"111111100",
95107=>"010011110",
95108=>"100101100",
95109=>"000000111",
95110=>"000100010",
95111=>"000010110",
95112=>"000100000",
95113=>"110100000",
95114=>"011001001",
95115=>"011111011",
95116=>"111001001",
95117=>"011001001",
95118=>"111101101",
95119=>"011001011",
95120=>"100111101",
95121=>"100110010",
95122=>"011001011",
95123=>"110110000",
95124=>"110010100",
95125=>"111000010",
95126=>"100100100",
95127=>"000111100",
95128=>"111100100",
95129=>"000100110",
95130=>"011001001",
95131=>"011001001",
95132=>"110100000",
95133=>"111000001",
95134=>"110110010",
95135=>"000100110",
95136=>"011011111",
95137=>"001001011",
95138=>"000110110",
95139=>"000011110",
95140=>"100100000",
95141=>"101101100",
95142=>"010110000",
95143=>"010110000",
95144=>"011001000",
95145=>"010100111",
95146=>"011001001",
95147=>"000001000",
95148=>"111101001",
95149=>"110000000",
95150=>"001000000",
95151=>"101001011",
95152=>"101000000",
95153=>"110110001",
95154=>"110000111",
95155=>"010001101",
95156=>"100110101",
95157=>"001001011",
95158=>"000001001",
95159=>"010001001",
95160=>"100000011",
95161=>"011100101",
95162=>"111011011",
95163=>"110110100",
95164=>"110100001",
95165=>"011011111",
95166=>"001001000",
95167=>"101011000",
95168=>"111001001",
95169=>"111001000",
95170=>"110110100",
95171=>"010000000",
95172=>"010011111",
95173=>"011011001",
95174=>"000100110",
95175=>"001001011",
95176=>"011110001",
95177=>"001110110",
95178=>"011010000",
95179=>"000100000",
95180=>"010001000",
95181=>"011111111",
95182=>"001000000",
95183=>"111000000",
95184=>"100001000",
95185=>"010000100",
95186=>"000110100",
95187=>"100110000",
95188=>"000010011",
95189=>"100000000",
95190=>"000110100",
95191=>"001000111",
95192=>"110100000",
95193=>"000101000",
95194=>"001001001",
95195=>"011001001",
95196=>"100001000",
95197=>"111101001",
95198=>"001001000",
95199=>"000101111",
95200=>"101111111",
95201=>"110001001",
95202=>"111011010",
95203=>"011110110",
95204=>"011000011",
95205=>"100110110",
95206=>"110000001",
95207=>"000001011",
95208=>"101001110",
95209=>"011001011",
95210=>"111001001",
95211=>"011001001",
95212=>"000110110",
95213=>"110011000",
95214=>"000000110",
95215=>"000111111",
95216=>"000000001",
95217=>"011000001",
95218=>"010110110",
95219=>"000000100",
95220=>"110001011",
95221=>"100001001",
95222=>"010001010",
95223=>"101001000",
95224=>"100001111",
95225=>"110110111",
95226=>"110111111",
95227=>"010111101",
95228=>"111011101",
95229=>"001001000",
95230=>"000011110",
95231=>"111011101",
95232=>"111011111",
95233=>"000111111",
95234=>"000010000",
95235=>"110000000",
95236=>"010100001",
95237=>"011000000",
95238=>"010010101",
95239=>"111101001",
95240=>"000000101",
95241=>"111111000",
95242=>"110010100",
95243=>"101111010",
95244=>"001000000",
95245=>"010000000",
95246=>"001001011",
95247=>"000110110",
95248=>"101111111",
95249=>"000000000",
95250=>"000000111",
95251=>"111100111",
95252=>"110101001",
95253=>"000000000",
95254=>"111111111",
95255=>"010110111",
95256=>"100000010",
95257=>"010001101",
95258=>"111111111",
95259=>"111111000",
95260=>"100000100",
95261=>"010000000",
95262=>"111100010",
95263=>"011111010",
95264=>"000000000",
95265=>"000011001",
95266=>"001101000",
95267=>"011100000",
95268=>"000000100",
95269=>"101001111",
95270=>"000010110",
95271=>"111111111",
95272=>"110111111",
95273=>"100000001",
95274=>"101100010",
95275=>"000000000",
95276=>"111110000",
95277=>"110111111",
95278=>"111111101",
95279=>"000000000",
95280=>"111111111",
95281=>"011001110",
95282=>"000000101",
95283=>"101000000",
95284=>"000001001",
95285=>"000000000",
95286=>"100001001",
95287=>"111111110",
95288=>"101111001",
95289=>"000000110",
95290=>"000000100",
95291=>"010110000",
95292=>"011010011",
95293=>"111111111",
95294=>"000001111",
95295=>"011111011",
95296=>"111011011",
95297=>"100100111",
95298=>"111111110",
95299=>"001000101",
95300=>"111111111",
95301=>"111101000",
95302=>"100000111",
95303=>"101101101",
95304=>"011111110",
95305=>"000000000",
95306=>"000000000",
95307=>"001000101",
95308=>"101000100",
95309=>"000000000",
95310=>"000000000",
95311=>"111111111",
95312=>"011111011",
95313=>"000000000",
95314=>"001101110",
95315=>"111110110",
95316=>"000001001",
95317=>"110000111",
95318=>"110110001",
95319=>"010010000",
95320=>"110000000",
95321=>"100111110",
95322=>"001011111",
95323=>"110111111",
95324=>"101111111",
95325=>"000000011",
95326=>"000000000",
95327=>"110010111",
95328=>"111111111",
95329=>"111111011",
95330=>"001001000",
95331=>"010110110",
95332=>"000000111",
95333=>"101111111",
95334=>"111110100",
95335=>"000100100",
95336=>"111000010",
95337=>"000010010",
95338=>"111001011",
95339=>"111111101",
95340=>"000101011",
95341=>"000000000",
95342=>"111000000",
95343=>"110110100",
95344=>"110110111",
95345=>"000010011",
95346=>"001101100",
95347=>"111110000",
95348=>"101001111",
95349=>"000000000",
95350=>"011000000",
95351=>"011111000",
95352=>"110100000",
95353=>"100001100",
95354=>"010111011",
95355=>"000000000",
95356=>"000111011",
95357=>"100000000",
95358=>"000101001",
95359=>"000100111",
95360=>"101111011",
95361=>"010110000",
95362=>"111110110",
95363=>"100100111",
95364=>"100101111",
95365=>"000001110",
95366=>"101100100",
95367=>"100110000",
95368=>"001001110",
95369=>"001011010",
95370=>"000001100",
95371=>"001111101",
95372=>"000101010",
95373=>"011000000",
95374=>"000000111",
95375=>"111001011",
95376=>"000000011",
95377=>"000111111",
95378=>"000000111",
95379=>"000000000",
95380=>"010111010",
95381=>"001000000",
95382=>"000000110",
95383=>"000101110",
95384=>"011000000",
95385=>"101000000",
95386=>"000111101",
95387=>"000001000",
95388=>"111101000",
95389=>"110111010",
95390=>"100101001",
95391=>"000000001",
95392=>"010011111",
95393=>"000111010",
95394=>"000001110",
95395=>"010000111",
95396=>"111000010",
95397=>"011111111",
95398=>"111000110",
95399=>"110010100",
95400=>"111111000",
95401=>"000111100",
95402=>"111111111",
95403=>"000000000",
95404=>"000000000",
95405=>"010111111",
95406=>"011111011",
95407=>"100110001",
95408=>"000000111",
95409=>"000000000",
95410=>"000000000",
95411=>"000111111",
95412=>"110110100",
95413=>"000000000",
95414=>"110000011",
95415=>"000110111",
95416=>"111010000",
95417=>"111000000",
95418=>"111101111",
95419=>"111011101",
95420=>"000011101",
95421=>"000001010",
95422=>"110110110",
95423=>"000000001",
95424=>"010000000",
95425=>"011000010",
95426=>"111101111",
95427=>"101000101",
95428=>"000110111",
95429=>"111000000",
95430=>"100101000",
95431=>"111110010",
95432=>"111000001",
95433=>"100100111",
95434=>"100101111",
95435=>"000001101",
95436=>"000000000",
95437=>"101011111",
95438=>"101001001",
95439=>"111111011",
95440=>"111000000",
95441=>"011111111",
95442=>"111111101",
95443=>"111111000",
95444=>"000000101",
95445=>"001000111",
95446=>"111101111",
95447=>"000001010",
95448=>"000001111",
95449=>"000001011",
95450=>"000110011",
95451=>"000111000",
95452=>"111011011",
95453=>"110110010",
95454=>"000010011",
95455=>"110111011",
95456=>"001111100",
95457=>"001000111",
95458=>"111111101",
95459=>"001011111",
95460=>"101000001",
95461=>"111000011",
95462=>"000001000",
95463=>"010011001",
95464=>"010001000",
95465=>"000000000",
95466=>"010011000",
95467=>"011110000",
95468=>"111101001",
95469=>"000101111",
95470=>"010010000",
95471=>"000100010",
95472=>"000000000",
95473=>"110000111",
95474=>"111111001",
95475=>"000000001",
95476=>"111100100",
95477=>"000000010",
95478=>"011100001",
95479=>"111111111",
95480=>"101001111",
95481=>"100001011",
95482=>"010001111",
95483=>"111011000",
95484=>"101111111",
95485=>"000001011",
95486=>"110001101",
95487=>"011011111",
95488=>"000010001",
95489=>"110010010",
95490=>"000100000",
95491=>"000000000",
95492=>"111111111",
95493=>"110110000",
95494=>"011111111",
95495=>"000011111",
95496=>"000000110",
95497=>"000101101",
95498=>"001001110",
95499=>"000111111",
95500=>"100010011",
95501=>"001111011",
95502=>"001010010",
95503=>"001101001",
95504=>"000111111",
95505=>"111111110",
95506=>"111001111",
95507=>"000000100",
95508=>"001111111",
95509=>"110101111",
95510=>"100100011",
95511=>"000000000",
95512=>"000000110",
95513=>"010111111",
95514=>"011001011",
95515=>"000001100",
95516=>"001111111",
95517=>"000100111",
95518=>"001011100",
95519=>"001101001",
95520=>"000000000",
95521=>"000111111",
95522=>"111111000",
95523=>"111011000",
95524=>"000111110",
95525=>"110100100",
95526=>"010111001",
95527=>"000000001",
95528=>"010110000",
95529=>"110111111",
95530=>"011000111",
95531=>"001101101",
95532=>"000000001",
95533=>"010111111",
95534=>"110111010",
95535=>"010110111",
95536=>"011010000",
95537=>"010001101",
95538=>"100111100",
95539=>"000000101",
95540=>"010000101",
95541=>"101001110",
95542=>"110100000",
95543=>"000000110",
95544=>"111101101",
95545=>"111001011",
95546=>"010011010",
95547=>"111000000",
95548=>"100110110",
95549=>"111101111",
95550=>"000000000",
95551=>"110111011",
95552=>"111000010",
95553=>"111111000",
95554=>"000000111",
95555=>"011111100",
95556=>"000000000",
95557=>"111111011",
95558=>"110001001",
95559=>"111100111",
95560=>"010110101",
95561=>"111000000",
95562=>"000000001",
95563=>"001000001",
95564=>"111111111",
95565=>"111111011",
95566=>"001100110",
95567=>"000000111",
95568=>"000011001",
95569=>"100111111",
95570=>"000000001",
95571=>"010010001",
95572=>"111110010",
95573=>"000001111",
95574=>"110110011",
95575=>"000111011",
95576=>"101001000",
95577=>"000000001",
95578=>"111100000",
95579=>"100100111",
95580=>"000000111",
95581=>"001000010",
95582=>"011101111",
95583=>"000001001",
95584=>"011010000",
95585=>"001111100",
95586=>"100101101",
95587=>"111000100",
95588=>"110000010",
95589=>"000000011",
95590=>"011010111",
95591=>"001101000",
95592=>"010010001",
95593=>"000011111",
95594=>"010111000",
95595=>"010001001",
95596=>"000110011",
95597=>"110111011",
95598=>"011011010",
95599=>"001111000",
95600=>"111100101",
95601=>"100000101",
95602=>"001000000",
95603=>"111111111",
95604=>"100111100",
95605=>"000000101",
95606=>"111010000",
95607=>"111111000",
95608=>"010000000",
95609=>"010010111",
95610=>"000001000",
95611=>"100110111",
95612=>"100100010",
95613=>"011011100",
95614=>"000000011",
95615=>"001111000",
95616=>"000000010",
95617=>"111111100",
95618=>"000110111",
95619=>"101100111",
95620=>"111111011",
95621=>"001001011",
95622=>"111011101",
95623=>"000001001",
95624=>"100110001",
95625=>"101101001",
95626=>"101110111",
95627=>"101001111",
95628=>"010010000",
95629=>"111000000",
95630=>"001101111",
95631=>"001000000",
95632=>"110111110",
95633=>"111110000",
95634=>"000000000",
95635=>"000000111",
95636=>"000000000",
95637=>"010000011",
95638=>"010010011",
95639=>"011010000",
95640=>"011111111",
95641=>"000000000",
95642=>"111111000",
95643=>"001000000",
95644=>"101000000",
95645=>"010111011",
95646=>"000010111",
95647=>"110010000",
95648=>"000010010",
95649=>"111010000",
95650=>"000010000",
95651=>"111101000",
95652=>"000000000",
95653=>"000110010",
95654=>"110010001",
95655=>"000010011",
95656=>"000000011",
95657=>"100000000",
95658=>"110010110",
95659=>"000111000",
95660=>"110000101",
95661=>"000100000",
95662=>"010010000",
95663=>"000000111",
95664=>"111111111",
95665=>"011111110",
95666=>"000111111",
95667=>"000101000",
95668=>"101010000",
95669=>"011000000",
95670=>"111011011",
95671=>"110111000",
95672=>"001011001",
95673=>"010110110",
95674=>"001000101",
95675=>"000110110",
95676=>"001001111",
95677=>"010111100",
95678=>"001010011",
95679=>"111100010",
95680=>"111101001",
95681=>"011011111",
95682=>"110111010",
95683=>"011011101",
95684=>"011101000",
95685=>"000110001",
95686=>"010000110",
95687=>"111001000",
95688=>"000111111",
95689=>"111000111",
95690=>"111110111",
95691=>"000101111",
95692=>"000111000",
95693=>"010001110",
95694=>"111111111",
95695=>"000100100",
95696=>"001111101",
95697=>"011010100",
95698=>"000000111",
95699=>"000010010",
95700=>"111010111",
95701=>"111111111",
95702=>"111101001",
95703=>"000000000",
95704=>"010000111",
95705=>"100100110",
95706=>"001000011",
95707=>"110011001",
95708=>"001100101",
95709=>"111000001",
95710=>"111000011",
95711=>"111101110",
95712=>"101101100",
95713=>"100000101",
95714=>"001000010",
95715=>"100000110",
95716=>"011000000",
95717=>"011111000",
95718=>"100110110",
95719=>"111001000",
95720=>"101111011",
95721=>"111111111",
95722=>"100100000",
95723=>"110110010",
95724=>"000101001",
95725=>"111110110",
95726=>"000011011",
95727=>"110010000",
95728=>"000000000",
95729=>"000110110",
95730=>"001000111",
95731=>"001000100",
95732=>"000011110",
95733=>"111111111",
95734=>"000100110",
95735=>"001101101",
95736=>"000000011",
95737=>"000010111",
95738=>"100111111",
95739=>"000001101",
95740=>"101000111",
95741=>"011111100",
95742=>"011111100",
95743=>"111010010",
95744=>"111011011",
95745=>"000000001",
95746=>"101100010",
95747=>"101001000",
95748=>"100100001",
95749=>"111001011",
95750=>"101101100",
95751=>"111100001",
95752=>"011000111",
95753=>"000000111",
95754=>"011001100",
95755=>"101011111",
95756=>"000001011",
95757=>"000000000",
95758=>"100100101",
95759=>"011111111",
95760=>"000000010",
95761=>"000000111",
95762=>"111111000",
95763=>"000000111",
95764=>"111110101",
95765=>"111111111",
95766=>"111101101",
95767=>"000010111",
95768=>"000000001",
95769=>"010111111",
95770=>"111000011",
95771=>"000000011",
95772=>"000000010",
95773=>"101011000",
95774=>"111110000",
95775=>"000000101",
95776=>"001010101",
95777=>"111011001",
95778=>"000110110",
95779=>"000010010",
95780=>"000111110",
95781=>"010011001",
95782=>"110010010",
95783=>"000110110",
95784=>"000011001",
95785=>"111111000",
95786=>"000000110",
95787=>"011111111",
95788=>"010000000",
95789=>"111100000",
95790=>"111101101",
95791=>"001101101",
95792=>"101001000",
95793=>"000101111",
95794=>"010000010",
95795=>"010000111",
95796=>"010011011",
95797=>"101000101",
95798=>"000000011",
95799=>"000000000",
95800=>"111101000",
95801=>"000000000",
95802=>"000000000",
95803=>"010000010",
95804=>"010000001",
95805=>"010111001",
95806=>"000000100",
95807=>"000111111",
95808=>"000111111",
95809=>"101000000",
95810=>"010000000",
95811=>"110001110",
95812=>"000000001",
95813=>"000100101",
95814=>"000001001",
95815=>"101111110",
95816=>"001000000",
95817=>"111000000",
95818=>"111111000",
95819=>"000011001",
95820=>"000000111",
95821=>"010000000",
95822=>"001001101",
95823=>"101000010",
95824=>"000000000",
95825=>"100101011",
95826=>"111001101",
95827=>"000000110",
95828=>"110100111",
95829=>"001111111",
95830=>"011011010",
95831=>"101010111",
95832=>"010000100",
95833=>"100000111",
95834=>"011001101",
95835=>"110011000",
95836=>"000111000",
95837=>"001000000",
95838=>"000111010",
95839=>"110100000",
95840=>"000111111",
95841=>"001000000",
95842=>"111000000",
95843=>"111111110",
95844=>"000001011",
95845=>"100111111",
95846=>"110000011",
95847=>"111000000",
95848=>"111111000",
95849=>"111111001",
95850=>"111000010",
95851=>"111000000",
95852=>"111000000",
95853=>"101000001",
95854=>"101001111",
95855=>"000000001",
95856=>"111111001",
95857=>"111101000",
95858=>"000000110",
95859=>"000000000",
95860=>"111100001",
95861=>"111000100",
95862=>"001000000",
95863=>"000110000",
95864=>"000001000",
95865=>"111111111",
95866=>"111111111",
95867=>"111110010",
95868=>"010001011",
95869=>"000100000",
95870=>"001011011",
95871=>"000001111",
95872=>"111111010",
95873=>"100111000",
95874=>"000010000",
95875=>"110111101",
95876=>"111111011",
95877=>"100110001",
95878=>"110100100",
95879=>"000010111",
95880=>"110111101",
95881=>"111111111",
95882=>"101000111",
95883=>"110010110",
95884=>"000110000",
95885=>"000000111",
95886=>"100000111",
95887=>"000000011",
95888=>"011001011",
95889=>"100000010",
95890=>"000010000",
95891=>"000010111",
95892=>"000010111",
95893=>"000000111",
95894=>"000011110",
95895=>"000100000",
95896=>"000001011",
95897=>"000000010",
95898=>"000010010",
95899=>"000100111",
95900=>"111100000",
95901=>"010110101",
95902=>"110111010",
95903=>"111101111",
95904=>"110101011",
95905=>"111001010",
95906=>"111010000",
95907=>"001001011",
95908=>"111101101",
95909=>"000110110",
95910=>"011010101",
95911=>"000000000",
95912=>"001000111",
95913=>"000001111",
95914=>"001101001",
95915=>"111101011",
95916=>"101111110",
95917=>"101000100",
95918=>"000001101",
95919=>"111111111",
95920=>"101110100",
95921=>"000000111",
95922=>"001100000",
95923=>"011011011",
95924=>"010000000",
95925=>"000000000",
95926=>"000111111",
95927=>"111010101",
95928=>"010100000",
95929=>"000110111",
95930=>"010000000",
95931=>"111010111",
95932=>"000111111",
95933=>"011111111",
95934=>"110111011",
95935=>"111000000",
95936=>"011111111",
95937=>"000000000",
95938=>"011100010",
95939=>"100111110",
95940=>"111111111",
95941=>"001111100",
95942=>"100010011",
95943=>"000111111",
95944=>"110111111",
95945=>"010110000",
95946=>"111111001",
95947=>"010111111",
95948=>"000000000",
95949=>"010100111",
95950=>"011101111",
95951=>"010111110",
95952=>"001000100",
95953=>"000001001",
95954=>"000000101",
95955=>"011100111",
95956=>"000010111",
95957=>"000000000",
95958=>"111000000",
95959=>"111100010",
95960=>"111001000",
95961=>"000010111",
95962=>"010111100",
95963=>"000010010",
95964=>"111011111",
95965=>"000001101",
95966=>"010000000",
95967=>"101000111",
95968=>"010000000",
95969=>"111000111",
95970=>"101011101",
95971=>"010111111",
95972=>"110000000",
95973=>"000111001",
95974=>"000000111",
95975=>"110011010",
95976=>"000000110",
95977=>"000000000",
95978=>"110100000",
95979=>"000111101",
95980=>"111110111",
95981=>"000011111",
95982=>"000010000",
95983=>"101000111",
95984=>"000000111",
95985=>"100101101",
95986=>"111011000",
95987=>"000001001",
95988=>"111100110",
95989=>"111110111",
95990=>"100000110",
95991=>"111111111",
95992=>"001111010",
95993=>"110111101",
95994=>"111010010",
95995=>"000011111",
95996=>"011111111",
95997=>"111110000",
95998=>"000111011",
95999=>"111111110",
96000=>"000100111",
96001=>"011011011",
96002=>"000100000",
96003=>"000000001",
96004=>"000010110",
96005=>"011111111",
96006=>"100111111",
96007=>"100011001",
96008=>"000000111",
96009=>"000011111",
96010=>"011110100",
96011=>"000010111",
96012=>"111110000",
96013=>"000011011",
96014=>"100101001",
96015=>"111001001",
96016=>"010000100",
96017=>"111010000",
96018=>"000000100",
96019=>"111111111",
96020=>"100101000",
96021=>"000000111",
96022=>"111100110",
96023=>"111111011",
96024=>"111011000",
96025=>"111000101",
96026=>"000000010",
96027=>"110100100",
96028=>"011011000",
96029=>"001001101",
96030=>"000111011",
96031=>"101000011",
96032=>"000111111",
96033=>"111000110",
96034=>"101000111",
96035=>"000010011",
96036=>"111110110",
96037=>"110111110",
96038=>"000010111",
96039=>"001000100",
96040=>"000000111",
96041=>"010000111",
96042=>"101000000",
96043=>"111000000",
96044=>"011000100",
96045=>"101000000",
96046=>"111111100",
96047=>"000000101",
96048=>"000110111",
96049=>"011001000",
96050=>"111111111",
96051=>"111111101",
96052=>"111111100",
96053=>"111100111",
96054=>"000110110",
96055=>"101000000",
96056=>"011000001",
96057=>"111111000",
96058=>"100000000",
96059=>"111110100",
96060=>"111011010",
96061=>"110100010",
96062=>"100001101",
96063=>"001010110",
96064=>"001101100",
96065=>"111111111",
96066=>"010000000",
96067=>"001011011",
96068=>"000000000",
96069=>"100000000",
96070=>"000111100",
96071=>"001011001",
96072=>"011101011",
96073=>"100111111",
96074=>"111101101",
96075=>"010100000",
96076=>"000011111",
96077=>"001001011",
96078=>"000000100",
96079=>"111101101",
96080=>"101101111",
96081=>"011000000",
96082=>"000011011",
96083=>"100100111",
96084=>"001000000",
96085=>"110011100",
96086=>"001011011",
96087=>"111111011",
96088=>"000000110",
96089=>"000000000",
96090=>"110110001",
96091=>"010100111",
96092=>"010000000",
96093=>"111100100",
96094=>"111101000",
96095=>"000110010",
96096=>"000010010",
96097=>"010001110",
96098=>"110110000",
96099=>"011001000",
96100=>"111101001",
96101=>"111111100",
96102=>"111100110",
96103=>"001001010",
96104=>"000101101",
96105=>"011001101",
96106=>"111111111",
96107=>"000011111",
96108=>"111011111",
96109=>"111101000",
96110=>"000000000",
96111=>"001001000",
96112=>"000001110",
96113=>"000000000",
96114=>"011011101",
96115=>"111101110",
96116=>"000000001",
96117=>"000000100",
96118=>"001000000",
96119=>"100000111",
96120=>"000111101",
96121=>"111010000",
96122=>"001101111",
96123=>"000000000",
96124=>"010000000",
96125=>"000001111",
96126=>"100001000",
96127=>"100011011",
96128=>"000010010",
96129=>"000010011",
96130=>"111010110",
96131=>"111000000",
96132=>"000001111",
96133=>"101101111",
96134=>"111111111",
96135=>"000100100",
96136=>"010110111",
96137=>"100100101",
96138=>"111100100",
96139=>"000000000",
96140=>"000000011",
96141=>"000000000",
96142=>"111111000",
96143=>"000000001",
96144=>"101111000",
96145=>"100000111",
96146=>"010011111",
96147=>"000000011",
96148=>"000000101",
96149=>"011010000",
96150=>"111011000",
96151=>"000100011",
96152=>"010011101",
96153=>"000000000",
96154=>"000010011",
96155=>"111111101",
96156=>"111111001",
96157=>"101100110",
96158=>"111011101",
96159=>"100110111",
96160=>"010011011",
96161=>"111000000",
96162=>"000001010",
96163=>"101000000",
96164=>"010111111",
96165=>"000001111",
96166=>"000000111",
96167=>"111111111",
96168=>"111100000",
96169=>"000001000",
96170=>"000010110",
96171=>"010110111",
96172=>"000000111",
96173=>"101000000",
96174=>"011111110",
96175=>"111101101",
96176=>"000111101",
96177=>"001001101",
96178=>"111011000",
96179=>"001000000",
96180=>"110110100",
96181=>"111111011",
96182=>"000110110",
96183=>"100100111",
96184=>"001100000",
96185=>"000000100",
96186=>"111111011",
96187=>"111011011",
96188=>"110110101",
96189=>"000111111",
96190=>"000000011",
96191=>"000000011",
96192=>"111101100",
96193=>"110000000",
96194=>"111111111",
96195=>"010000100",
96196=>"001000100",
96197=>"011000000",
96198=>"000011111",
96199=>"010000000",
96200=>"100111000",
96201=>"111000100",
96202=>"111011111",
96203=>"011011110",
96204=>"100100110",
96205=>"011000000",
96206=>"000000000",
96207=>"000110100",
96208=>"100010010",
96209=>"000010110",
96210=>"101101111",
96211=>"111100000",
96212=>"000000100",
96213=>"011001111",
96214=>"111011011",
96215=>"111000100",
96216=>"101100100",
96217=>"011011111",
96218=>"011100000",
96219=>"000000101",
96220=>"111000001",
96221=>"010011011",
96222=>"100101100",
96223=>"000011111",
96224=>"101100100",
96225=>"100101000",
96226=>"111000000",
96227=>"000000001",
96228=>"000000111",
96229=>"010110010",
96230=>"101011111",
96231=>"100000000",
96232=>"111111101",
96233=>"000000000",
96234=>"110111101",
96235=>"111111111",
96236=>"000000100",
96237=>"001010110",
96238=>"000000000",
96239=>"000000010",
96240=>"000010111",
96241=>"011101110",
96242=>"011010001",
96243=>"111001000",
96244=>"011010010",
96245=>"001101101",
96246=>"100000010",
96247=>"101110100",
96248=>"111111000",
96249=>"110101101",
96250=>"111100010",
96251=>"001001100",
96252=>"111010000",
96253=>"000000100",
96254=>"000110000",
96255=>"111111000",
96256=>"011011100",
96257=>"000100111",
96258=>"111000000",
96259=>"000000010",
96260=>"110110011",
96261=>"000000000",
96262=>"110101111",
96263=>"000000110",
96264=>"001101001",
96265=>"111011110",
96266=>"011111111",
96267=>"011001000",
96268=>"000000000",
96269=>"111111111",
96270=>"110110010",
96271=>"000000001",
96272=>"000111001",
96273=>"010111111",
96274=>"110110000",
96275=>"000011111",
96276=>"111110011",
96277=>"110000111",
96278=>"110111110",
96279=>"110111111",
96280=>"111001111",
96281=>"111001001",
96282=>"000000110",
96283=>"111111110",
96284=>"111111010",
96285=>"101000000",
96286=>"110000000",
96287=>"010110000",
96288=>"110110010",
96289=>"111111100",
96290=>"000101001",
96291=>"000111111",
96292=>"111111010",
96293=>"110010110",
96294=>"000111101",
96295=>"001111111",
96296=>"000001111",
96297=>"000000110",
96298=>"010111001",
96299=>"111111111",
96300=>"110111111",
96301=>"000000001",
96302=>"101000111",
96303=>"000000000",
96304=>"000000000",
96305=>"111111001",
96306=>"000010000",
96307=>"111110000",
96308=>"101111000",
96309=>"000000000",
96310=>"111111011",
96311=>"001000000",
96312=>"111110010",
96313=>"101111111",
96314=>"010000000",
96315=>"110110010",
96316=>"011001001",
96317=>"100111101",
96318=>"000000000",
96319=>"001000110",
96320=>"111111000",
96321=>"000100000",
96322=>"000100111",
96323=>"010000110",
96324=>"110111111",
96325=>"000001011",
96326=>"010011010",
96327=>"000000001",
96328=>"001010001",
96329=>"000000111",
96330=>"001001111",
96331=>"000000000",
96332=>"000000000",
96333=>"010110000",
96334=>"110110110",
96335=>"010000110",
96336=>"001100101",
96337=>"110111110",
96338=>"011011111",
96339=>"011000000",
96340=>"000000010",
96341=>"100000100",
96342=>"110110100",
96343=>"101000111",
96344=>"111111111",
96345=>"000000011",
96346=>"111111111",
96347=>"000000000",
96348=>"001101101",
96349=>"111100110",
96350=>"110111111",
96351=>"111111111",
96352=>"111111111",
96353=>"110011111",
96354=>"111111000",
96355=>"110110001",
96356=>"001011011",
96357=>"001000000",
96358=>"110111100",
96359=>"001000000",
96360=>"011000001",
96361=>"011000000",
96362=>"011111110",
96363=>"000000010",
96364=>"110000111",
96365=>"110111110",
96366=>"011010000",
96367=>"111111110",
96368=>"110100100",
96369=>"110000000",
96370=>"111111100",
96371=>"000110000",
96372=>"111111001",
96373=>"000000001",
96374=>"000101000",
96375=>"101001010",
96376=>"000101101",
96377=>"110111111",
96378=>"011111111",
96379=>"000000000",
96380=>"110111110",
96381=>"000000000",
96382=>"000001111",
96383=>"111001000",
96384=>"000111000",
96385=>"111100000",
96386=>"111000001",
96387=>"000000000",
96388=>"111011110",
96389=>"000001001",
96390=>"111111110",
96391=>"011111000",
96392=>"111010010",
96393=>"000000001",
96394=>"000111011",
96395=>"001000000",
96396=>"110101101",
96397=>"111110111",
96398=>"000000000",
96399=>"000001001",
96400=>"100000000",
96401=>"000101111",
96402=>"000000011",
96403=>"000011001",
96404=>"110010100",
96405=>"111101010",
96406=>"000000000",
96407=>"000100000",
96408=>"110111100",
96409=>"000000000",
96410=>"000000010",
96411=>"000000000",
96412=>"110110110",
96413=>"111000110",
96414=>"111001001",
96415=>"000000000",
96416=>"001001001",
96417=>"111110000",
96418=>"000000000",
96419=>"000000001",
96420=>"011011111",
96421=>"000000000",
96422=>"000100000",
96423=>"000000000",
96424=>"000111111",
96425=>"000000100",
96426=>"111110111",
96427=>"111110111",
96428=>"000001111",
96429=>"101000100",
96430=>"111110110",
96431=>"000011001",
96432=>"000000111",
96433=>"110110100",
96434=>"110100000",
96435=>"111010000",
96436=>"000000000",
96437=>"000000000",
96438=>"001000000",
96439=>"111111111",
96440=>"010100100",
96441=>"100111001",
96442=>"111111111",
96443=>"000001111",
96444=>"000000000",
96445=>"111110100",
96446=>"100000000",
96447=>"000000111",
96448=>"101001000",
96449=>"011000000",
96450=>"001000000",
96451=>"001000001",
96452=>"000001111",
96453=>"110100110",
96454=>"000000111",
96455=>"000110110",
96456=>"011000000",
96457=>"000000000",
96458=>"000000111",
96459=>"000000000",
96460=>"111011000",
96461=>"111111111",
96462=>"001101000",
96463=>"100001001",
96464=>"111110000",
96465=>"110110000",
96466=>"100011000",
96467=>"000000000",
96468=>"001001111",
96469=>"010111011",
96470=>"111111000",
96471=>"000000000",
96472=>"000000001",
96473=>"010111111",
96474=>"100000000",
96475=>"000000000",
96476=>"011111110",
96477=>"111010000",
96478=>"000010000",
96479=>"111101111",
96480=>"000000000",
96481=>"110101101",
96482=>"000111111",
96483=>"000001100",
96484=>"000000001",
96485=>"111111100",
96486=>"111111111",
96487=>"111111011",
96488=>"000111111",
96489=>"010111111",
96490=>"111111111",
96491=>"000010111",
96492=>"011111111",
96493=>"000111111",
96494=>"110110000",
96495=>"111000111",
96496=>"111010001",
96497=>"111011011",
96498=>"110000001",
96499=>"110110100",
96500=>"100100000",
96501=>"110110111",
96502=>"000000000",
96503=>"000000000",
96504=>"011000000",
96505=>"000000000",
96506=>"000000000",
96507=>"111001000",
96508=>"100101101",
96509=>"000010000",
96510=>"100011000",
96511=>"001000000",
96512=>"100000001",
96513=>"111011000",
96514=>"111000000",
96515=>"101111000",
96516=>"111100100",
96517=>"001110001",
96518=>"111111111",
96519=>"111101101",
96520=>"000001110",
96521=>"000101111",
96522=>"110111000",
96523=>"111111000",
96524=>"000100111",
96525=>"110110000",
96526=>"000001000",
96527=>"111111100",
96528=>"000111111",
96529=>"000111111",
96530=>"111001101",
96531=>"001000000",
96532=>"101111111",
96533=>"111000000",
96534=>"111000100",
96535=>"111111000",
96536=>"111000000",
96537=>"111011111",
96538=>"111101001",
96539=>"100111111",
96540=>"100000010",
96541=>"111000000",
96542=>"111000000",
96543=>"001000000",
96544=>"110110000",
96545=>"111101000",
96546=>"011111001",
96547=>"000000101",
96548=>"100111011",
96549=>"111001000",
96550=>"111001000",
96551=>"000001111",
96552=>"111001000",
96553=>"110100000",
96554=>"110000000",
96555=>"110000111",
96556=>"011111001",
96557=>"111101010",
96558=>"111000000",
96559=>"111011111",
96560=>"000100000",
96561=>"101111100",
96562=>"111101000",
96563=>"111011000",
96564=>"001000100",
96565=>"000000100",
96566=>"001110000",
96567=>"111111111",
96568=>"111111111",
96569=>"110110000",
96570=>"011111000",
96571=>"111111000",
96572=>"000010100",
96573=>"111011010",
96574=>"001000100",
96575=>"011011000",
96576=>"010000111",
96577=>"000000101",
96578=>"100001111",
96579=>"100101111",
96580=>"011011011",
96581=>"010000001",
96582=>"111111000",
96583=>"110111111",
96584=>"111011011",
96585=>"000000111",
96586=>"111000111",
96587=>"000110111",
96588=>"000001101",
96589=>"000011110",
96590=>"100110011",
96591=>"111010111",
96592=>"111101000",
96593=>"111010010",
96594=>"000000000",
96595=>"000111011",
96596=>"101101111",
96597=>"011100101",
96598=>"011000000",
96599=>"000101101",
96600=>"101101000",
96601=>"000111110",
96602=>"111101000",
96603=>"000111111",
96604=>"000001111",
96605=>"000000000",
96606=>"111000011",
96607=>"001000001",
96608=>"000000000",
96609=>"001101000",
96610=>"011101111",
96611=>"111101000",
96612=>"000010010",
96613=>"000100011",
96614=>"001001110",
96615=>"000000110",
96616=>"111000000",
96617=>"101001001",
96618=>"000000101",
96619=>"010000000",
96620=>"010000001",
96621=>"000011010",
96622=>"000000111",
96623=>"111111001",
96624=>"110100010",
96625=>"100111111",
96626=>"111011001",
96627=>"000000000",
96628=>"111111111",
96629=>"000100000",
96630=>"111010000",
96631=>"000000010",
96632=>"000001000",
96633=>"000101000",
96634=>"110010111",
96635=>"001000010",
96636=>"111111001",
96637=>"000001000",
96638=>"111111110",
96639=>"000000111",
96640=>"000000011",
96641=>"111100110",
96642=>"000010111",
96643=>"100000000",
96644=>"000000000",
96645=>"000011111",
96646=>"011000000",
96647=>"010011001",
96648=>"000001111",
96649=>"101000111",
96650=>"111100000",
96651=>"000110111",
96652=>"011000111",
96653=>"000111110",
96654=>"000000111",
96655=>"000100111",
96656=>"011110111",
96657=>"111101101",
96658=>"010000000",
96659=>"010000101",
96660=>"001110110",
96661=>"000000010",
96662=>"111110100",
96663=>"001100110",
96664=>"000111111",
96665=>"110000000",
96666=>"111000000",
96667=>"011000000",
96668=>"100001111",
96669=>"010000100",
96670=>"111111111",
96671=>"000100010",
96672=>"001111110",
96673=>"111101000",
96674=>"000000000",
96675=>"100111101",
96676=>"001000000",
96677=>"000100110",
96678=>"000010111",
96679=>"001101000",
96680=>"000011111",
96681=>"000101011",
96682=>"111111111",
96683=>"001000110",
96684=>"111011111",
96685=>"000101111",
96686=>"011111000",
96687=>"000101111",
96688=>"001001011",
96689=>"110110000",
96690=>"001101010",
96691=>"100000001",
96692=>"001100111",
96693=>"011011000",
96694=>"011000000",
96695=>"011010000",
96696=>"000001001",
96697=>"100110110",
96698=>"011000000",
96699=>"111111101",
96700=>"000111101",
96701=>"111111000",
96702=>"000100001",
96703=>"101111110",
96704=>"100001010",
96705=>"000000111",
96706=>"000010100",
96707=>"110110110",
96708=>"000000100",
96709=>"100011001",
96710=>"000000000",
96711=>"000000111",
96712=>"110111111",
96713=>"000000111",
96714=>"100001101",
96715=>"000000001",
96716=>"111100000",
96717=>"111000110",
96718=>"111001000",
96719=>"111111100",
96720=>"111111000",
96721=>"110011001",
96722=>"000010111",
96723=>"000111111",
96724=>"000001111",
96725=>"111101100",
96726=>"111100100",
96727=>"111111111",
96728=>"000011111",
96729=>"000000010",
96730=>"101111001",
96731=>"000011010",
96732=>"110000011",
96733=>"001100010",
96734=>"000111111",
96735=>"101111111",
96736=>"100000000",
96737=>"100000111",
96738=>"001001111",
96739=>"001110110",
96740=>"000000110",
96741=>"000000000",
96742=>"000100000",
96743=>"010011010",
96744=>"000000111",
96745=>"010000011",
96746=>"111110000",
96747=>"010000001",
96748=>"110000111",
96749=>"111111001",
96750=>"000000000",
96751=>"000100110",
96752=>"110100000",
96753=>"101100100",
96754=>"000010100",
96755=>"000111001",
96756=>"001111110",
96757=>"111001000",
96758=>"100000100",
96759=>"000000111",
96760=>"100100111",
96761=>"101111000",
96762=>"110100010",
96763=>"000010111",
96764=>"111010000",
96765=>"000000101",
96766=>"000000000",
96767=>"001000111",
96768=>"111111000",
96769=>"000111011",
96770=>"000110110",
96771=>"000000011",
96772=>"011111110",
96773=>"000000000",
96774=>"111001011",
96775=>"010000001",
96776=>"100111111",
96777=>"111101111",
96778=>"010100100",
96779=>"111000010",
96780=>"101000000",
96781=>"111110000",
96782=>"000001001",
96783=>"000000100",
96784=>"000000001",
96785=>"001001001",
96786=>"010100101",
96787=>"001100000",
96788=>"101000111",
96789=>"010111110",
96790=>"011110000",
96791=>"011111101",
96792=>"100100100",
96793=>"101100111",
96794=>"010000100",
96795=>"000000000",
96796=>"101111111",
96797=>"101111110",
96798=>"000110111",
96799=>"001001011",
96800=>"010111011",
96801=>"000000000",
96802=>"000111111",
96803=>"111011111",
96804=>"000100110",
96805=>"100100010",
96806=>"010111000",
96807=>"101111001",
96808=>"111111111",
96809=>"000000000",
96810=>"111010010",
96811=>"000000000",
96812=>"000100100",
96813=>"010000000",
96814=>"010000000",
96815=>"001000000",
96816=>"110000001",
96817=>"000000000",
96818=>"000110111",
96819=>"100000001",
96820=>"000000010",
96821=>"111111000",
96822=>"000100010",
96823=>"011111111",
96824=>"010111111",
96825=>"000000000",
96826=>"000000101",
96827=>"000000000",
96828=>"011011111",
96829=>"111111011",
96830=>"000000000",
96831=>"101110000",
96832=>"111101101",
96833=>"111100001",
96834=>"000000000",
96835=>"011001100",
96836=>"000000111",
96837=>"101000001",
96838=>"110011011",
96839=>"111110111",
96840=>"000000000",
96841=>"011010010",
96842=>"101000000",
96843=>"011001011",
96844=>"000100111",
96845=>"001111111",
96846=>"100000000",
96847=>"000000000",
96848=>"100100100",
96849=>"000111111",
96850=>"000000101",
96851=>"001000000",
96852=>"111111010",
96853=>"001100100",
96854=>"001001101",
96855=>"000110101",
96856=>"111000110",
96857=>"000000001",
96858=>"011100000",
96859=>"011001100",
96860=>"011111110",
96861=>"001001011",
96862=>"010111011",
96863=>"111111011",
96864=>"000000100",
96865=>"000101001",
96866=>"000000101",
96867=>"100110000",
96868=>"100100111",
96869=>"100000000",
96870=>"100000001",
96871=>"110110111",
96872=>"111111010",
96873=>"000100111",
96874=>"110100100",
96875=>"010000010",
96876=>"101101101",
96877=>"101111000",
96878=>"000000000",
96879=>"000000111",
96880=>"001000011",
96881=>"000000000",
96882=>"000000000",
96883=>"010010011",
96884=>"000000011",
96885=>"000000111",
96886=>"111110111",
96887=>"100100011",
96888=>"000111111",
96889=>"001001111",
96890=>"000000111",
96891=>"101101101",
96892=>"100110111",
96893=>"100100000",
96894=>"011010000",
96895=>"010011111",
96896=>"111101011",
96897=>"111011010",
96898=>"100000101",
96899=>"000001101",
96900=>"100000000",
96901=>"111101001",
96902=>"011001110",
96903=>"000100000",
96904=>"100011011",
96905=>"101000000",
96906=>"011011000",
96907=>"100010000",
96908=>"011111010",
96909=>"011111111",
96910=>"001011011",
96911=>"100000001",
96912=>"001001001",
96913=>"111000010",
96914=>"011011000",
96915=>"000000001",
96916=>"101111111",
96917=>"000000100",
96918=>"111111111",
96919=>"000000000",
96920=>"101010110",
96921=>"001111111",
96922=>"000111010",
96923=>"000000000",
96924=>"101111000",
96925=>"101000000",
96926=>"000000111",
96927=>"111101000",
96928=>"100011101",
96929=>"010011010",
96930=>"000011000",
96931=>"000010000",
96932=>"011101000",
96933=>"111101111",
96934=>"000110000",
96935=>"100111111",
96936=>"111110111",
96937=>"011000100",
96938=>"000000000",
96939=>"000000000",
96940=>"000001000",
96941=>"000000001",
96942=>"111111110",
96943=>"111111110",
96944=>"111110000",
96945=>"111011000",
96946=>"000000100",
96947=>"100100100",
96948=>"001111000",
96949=>"111111010",
96950=>"100100100",
96951=>"000000000",
96952=>"100111111",
96953=>"100110100",
96954=>"000000100",
96955=>"011111111",
96956=>"000000111",
96957=>"001001111",
96958=>"110011111",
96959=>"111111111",
96960=>"000111111",
96961=>"111011010",
96962=>"001110010",
96963=>"000000000",
96964=>"001000000",
96965=>"001100010",
96966=>"111110111",
96967=>"100000011",
96968=>"001111001",
96969=>"111100111",
96970=>"111111111",
96971=>"010111000",
96972=>"001000011",
96973=>"001001011",
96974=>"000000000",
96975=>"000101001",
96976=>"011111110",
96977=>"001001000",
96978=>"011000110",
96979=>"001000111",
96980=>"011011010",
96981=>"100111111",
96982=>"000000100",
96983=>"000001011",
96984=>"011111000",
96985=>"111101101",
96986=>"001101101",
96987=>"001000000",
96988=>"110011110",
96989=>"011010111",
96990=>"010000111",
96991=>"110111111",
96992=>"000000101",
96993=>"100000001",
96994=>"101101000",
96995=>"100000000",
96996=>"010000000",
96997=>"010010011",
96998=>"101000000",
96999=>"111111011",
97000=>"101000000",
97001=>"110111101",
97002=>"110011001",
97003=>"000010101",
97004=>"000000000",
97005=>"101101111",
97006=>"000000000",
97007=>"100000010",
97008=>"101000000",
97009=>"010001000",
97010=>"000000101",
97011=>"000000000",
97012=>"101000101",
97013=>"010111001",
97014=>"000000111",
97015=>"000000000",
97016=>"000100111",
97017=>"000000100",
97018=>"010111110",
97019=>"001101101",
97020=>"010110100",
97021=>"000000000",
97022=>"100100111",
97023=>"110100001",
97024=>"011110000",
97025=>"010000010",
97026=>"000010110",
97027=>"000000001",
97028=>"000011001",
97029=>"010000000",
97030=>"000000101",
97031=>"111000100",
97032=>"111011100",
97033=>"011010010",
97034=>"110111001",
97035=>"000000000",
97036=>"111111111",
97037=>"111111000",
97038=>"100011111",
97039=>"110001111",
97040=>"010000010",
97041=>"111111010",
97042=>"000001101",
97043=>"011010110",
97044=>"010000111",
97045=>"100000000",
97046=>"111000000",
97047=>"100100111",
97048=>"101100101",
97049=>"111111110",
97050=>"011101000",
97051=>"000010000",
97052=>"010000011",
97053=>"100000111",
97054=>"011110010",
97055=>"001111011",
97056=>"000000000",
97057=>"000000010",
97058=>"100000011",
97059=>"000000000",
97060=>"100110110",
97061=>"110101000",
97062=>"000000101",
97063=>"111111011",
97064=>"010100000",
97065=>"011000000",
97066=>"010000010",
97067=>"011000000",
97068=>"111000100",
97069=>"111000110",
97070=>"111101101",
97071=>"110100111",
97072=>"111111011",
97073=>"100100001",
97074=>"100000001",
97075=>"111011010",
97076=>"011011010",
97077=>"001110110",
97078=>"110000001",
97079=>"000000001",
97080=>"000000000",
97081=>"001001111",
97082=>"000000101",
97083=>"000010000",
97084=>"100000001",
97085=>"111101111",
97086=>"000010000",
97087=>"100000100",
97088=>"000111011",
97089=>"111001111",
97090=>"000000000",
97091=>"000000101",
97092=>"111110110",
97093=>"010000101",
97094=>"111111000",
97095=>"000010100",
97096=>"101001101",
97097=>"011111000",
97098=>"101101111",
97099=>"111111111",
97100=>"000001101",
97101=>"011011011",
97102=>"011011100",
97103=>"100000000",
97104=>"000001101",
97105=>"010000010",
97106=>"111000111",
97107=>"001110110",
97108=>"010010000",
97109=>"100100010",
97110=>"000000000",
97111=>"010110000",
97112=>"110111111",
97113=>"111111011",
97114=>"110110110",
97115=>"000100100",
97116=>"001000000",
97117=>"001000001",
97118=>"111111110",
97119=>"000000001",
97120=>"101000101",
97121=>"001000000",
97122=>"000000101",
97123=>"000001000",
97124=>"101001101",
97125=>"001100100",
97126=>"000001011",
97127=>"001101101",
97128=>"000000111",
97129=>"111100000",
97130=>"111001000",
97131=>"111000111",
97132=>"100000000",
97133=>"111111101",
97134=>"111000000",
97135=>"111111111",
97136=>"011110101",
97137=>"000000110",
97138=>"011000010",
97139=>"000111101",
97140=>"101111111",
97141=>"000000111",
97142=>"001110111",
97143=>"110000100",
97144=>"010010010",
97145=>"111000000",
97146=>"000000010",
97147=>"111001101",
97148=>"000110100",
97149=>"100101101",
97150=>"011000000",
97151=>"000001101",
97152=>"011000000",
97153=>"000000010",
97154=>"111000000",
97155=>"111100011",
97156=>"111101111",
97157=>"101101101",
97158=>"011001100",
97159=>"000001101",
97160=>"100101100",
97161=>"111001101",
97162=>"001000000",
97163=>"000011111",
97164=>"000000000",
97165=>"011110110",
97166=>"101101101",
97167=>"000000100",
97168=>"100100110",
97169=>"111000100",
97170=>"111000000",
97171=>"000010010",
97172=>"000010100",
97173=>"010010110",
97174=>"010010010",
97175=>"000000010",
97176=>"010000010",
97177=>"111010010",
97178=>"010011010",
97179=>"001010000",
97180=>"000001001",
97181=>"000111111",
97182=>"000111111",
97183=>"001000001",
97184=>"001101001",
97185=>"000011010",
97186=>"111111101",
97187=>"000000010",
97188=>"000000011",
97189=>"100001001",
97190=>"110010111",
97191=>"010111010",
97192=>"011010110",
97193=>"000000000",
97194=>"110111110",
97195=>"000011010",
97196=>"111000100",
97197=>"010011000",
97198=>"100100101",
97199=>"010100101",
97200=>"111100111",
97201=>"001110111",
97202=>"000000101",
97203=>"000110000",
97204=>"001101101",
97205=>"100111111",
97206=>"111000100",
97207=>"011111110",
97208=>"000000000",
97209=>"000100101",
97210=>"111000010",
97211=>"001010010",
97212=>"011100000",
97213=>"110111111",
97214=>"001100001",
97215=>"011000000",
97216=>"010000010",
97217=>"101101111",
97218=>"000110111",
97219=>"001001000",
97220=>"000000111",
97221=>"110010010",
97222=>"111111000",
97223=>"010111111",
97224=>"000000000",
97225=>"111101011",
97226=>"000000110",
97227=>"101000111",
97228=>"111100000",
97229=>"000010000",
97230=>"001111000",
97231=>"000000011",
97232=>"000010100",
97233=>"101000101",
97234=>"000111110",
97235=>"111111101",
97236=>"000000111",
97237=>"111111101",
97238=>"110010000",
97239=>"100101101",
97240=>"000000001",
97241=>"111000000",
97242=>"100101101",
97243=>"000001111",
97244=>"000000010",
97245=>"010000111",
97246=>"010110111",
97247=>"000000010",
97248=>"010010000",
97249=>"111111111",
97250=>"000001000",
97251=>"010001110",
97252=>"010111010",
97253=>"110000000",
97254=>"001000001",
97255=>"011001000",
97256=>"000000000",
97257=>"111101100",
97258=>"011111110",
97259=>"111111111",
97260=>"111111000",
97261=>"000111011",
97262=>"000010000",
97263=>"000000111",
97264=>"000000010",
97265=>"011011100",
97266=>"111000000",
97267=>"101101101",
97268=>"111101001",
97269=>"101101100",
97270=>"100000000",
97271=>"000000000",
97272=>"000000011",
97273=>"000000111",
97274=>"010000110",
97275=>"000110101",
97276=>"100000010",
97277=>"101100100",
97278=>"110110111",
97279=>"001000000",
97280=>"100100100",
97281=>"101111010",
97282=>"111000000",
97283=>"110111111",
97284=>"000101101",
97285=>"110101000",
97286=>"000111011",
97287=>"000111111",
97288=>"111000000",
97289=>"011000101",
97290=>"000000000",
97291=>"000001110",
97292=>"001101001",
97293=>"110010010",
97294=>"100011001",
97295=>"101000001",
97296=>"100010100",
97297=>"000000000",
97298=>"110000010",
97299=>"101111011",
97300=>"111111000",
97301=>"011111001",
97302=>"000101011",
97303=>"111111111",
97304=>"000000111",
97305=>"010000110",
97306=>"000000000",
97307=>"000101111",
97308=>"111000010",
97309=>"001001010",
97310=>"010100101",
97311=>"000000000",
97312=>"000000000",
97313=>"010001101",
97314=>"010010010",
97315=>"111111111",
97316=>"101100000",
97317=>"001011001",
97318=>"000111010",
97319=>"011011001",
97320=>"000101111",
97321=>"100111000",
97322=>"000000010",
97323=>"010111010",
97324=>"000111101",
97325=>"101100011",
97326=>"110000000",
97327=>"111001000",
97328=>"011011000",
97329=>"100000000",
97330=>"000001111",
97331=>"000111111",
97332=>"001001000",
97333=>"110010100",
97334=>"001001001",
97335=>"110110000",
97336=>"101110000",
97337=>"000111111",
97338=>"000000100",
97339=>"000111111",
97340=>"001011011",
97341=>"111000011",
97342=>"000000101",
97343=>"001001000",
97344=>"111111111",
97345=>"010101010",
97346=>"011110011",
97347=>"111100001",
97348=>"111111111",
97349=>"010010000",
97350=>"000000111",
97351=>"100010010",
97352=>"001101011",
97353=>"001101111",
97354=>"001001001",
97355=>"011000001",
97356=>"111011111",
97357=>"100101101",
97358=>"010000000",
97359=>"101111111",
97360=>"000000000",
97361=>"101111111",
97362=>"111101010",
97363=>"110110100",
97364=>"110100101",
97365=>"100001000",
97366=>"101101001",
97367=>"111001101",
97368=>"001011101",
97369=>"001101001",
97370=>"001101101",
97371=>"111000000",
97372=>"001010000",
97373=>"000001111",
97374=>"111111000",
97375=>"101001000",
97376=>"111110000",
97377=>"000000011",
97378=>"111000000",
97379=>"100111111",
97380=>"000100101",
97381=>"000000101",
97382=>"000101011",
97383=>"000000010",
97384=>"110111001",
97385=>"000100010",
97386=>"001001000",
97387=>"111000011",
97388=>"001010000",
97389=>"010000100",
97390=>"011000000",
97391=>"000101111",
97392=>"001001100",
97393=>"011101111",
97394=>"100100100",
97395=>"011000001",
97396=>"101101010",
97397=>"000000110",
97398=>"010100101",
97399=>"011000000",
97400=>"000010000",
97401=>"000100010",
97402=>"000000101",
97403=>"000000000",
97404=>"000000101",
97405=>"011001001",
97406=>"111101000",
97407=>"111000000",
97408=>"111101101",
97409=>"110011000",
97410=>"101100000",
97411=>"100101110",
97412=>"111011111",
97413=>"101111111",
97414=>"100100110",
97415=>"000001001",
97416=>"100101011",
97417=>"011111111",
97418=>"010100011",
97419=>"001001001",
97420=>"010101111",
97421=>"011011000",
97422=>"001111010",
97423=>"011000111",
97424=>"001101101",
97425=>"110111111",
97426=>"000001111",
97427=>"110111101",
97428=>"111011101",
97429=>"111001000",
97430=>"110001001",
97431=>"001011000",
97432=>"000100000",
97433=>"111111111",
97434=>"111111111",
97435=>"111111000",
97436=>"011111111",
97437=>"110010010",
97438=>"000001111",
97439=>"000000101",
97440=>"000000000",
97441=>"001001111",
97442=>"111111011",
97443=>"111111111",
97444=>"010001100",
97445=>"001001001",
97446=>"000100111",
97447=>"000000000",
97448=>"010000010",
97449=>"111110000",
97450=>"111000000",
97451=>"011000000",
97452=>"010000111",
97453=>"000000000",
97454=>"001011001",
97455=>"001001010",
97456=>"101010010",
97457=>"000100100",
97458=>"001101111",
97459=>"000100101",
97460=>"100101011",
97461=>"000001010",
97462=>"010000101",
97463=>"000101111",
97464=>"100100101",
97465=>"111100111",
97466=>"111111100",
97467=>"101111101",
97468=>"000000000",
97469=>"111010010",
97470=>"111000000",
97471=>"000000000",
97472=>"000101101",
97473=>"000111001",
97474=>"011111111",
97475=>"100100100",
97476=>"011000000",
97477=>"101001011",
97478=>"111011111",
97479=>"111010000",
97480=>"011000000",
97481=>"010001000",
97482=>"010000110",
97483=>"011111100",
97484=>"100111000",
97485=>"000001101",
97486=>"110000000",
97487=>"111001011",
97488=>"001101111",
97489=>"000000000",
97490=>"110110111",
97491=>"110101000",
97492=>"000000000",
97493=>"000101011",
97494=>"000100000",
97495=>"101001000",
97496=>"101111011",
97497=>"000011011",
97498=>"000001001",
97499=>"011000000",
97500=>"001101100",
97501=>"101111011",
97502=>"011010010",
97503=>"001110110",
97504=>"111000000",
97505=>"000000111",
97506=>"101111010",
97507=>"011101100",
97508=>"010000101",
97509=>"000001001",
97510=>"111000000",
97511=>"000101111",
97512=>"011111011",
97513=>"000111111",
97514=>"100000000",
97515=>"000001001",
97516=>"000000000",
97517=>"110101110",
97518=>"100000000",
97519=>"011000000",
97520=>"101000100",
97521=>"010000100",
97522=>"000101000",
97523=>"001111000",
97524=>"001001111",
97525=>"000000001",
97526=>"100000101",
97527=>"000011010",
97528=>"111111000",
97529=>"001111011",
97530=>"000111111",
97531=>"000000111",
97532=>"111111010",
97533=>"000110000",
97534=>"000001001",
97535=>"110111000",
97536=>"000011110",
97537=>"100111001",
97538=>"100000000",
97539=>"100000111",
97540=>"000011010",
97541=>"101001111",
97542=>"000000000",
97543=>"000010000",
97544=>"000000101",
97545=>"000010000",
97546=>"000011000",
97547=>"100000101",
97548=>"101010010",
97549=>"000000000",
97550=>"101011001",
97551=>"111111000",
97552=>"100010010",
97553=>"000000010",
97554=>"101100101",
97555=>"000010011",
97556=>"111111010",
97557=>"101000100",
97558=>"001000100",
97559=>"111111010",
97560=>"000101001",
97561=>"000111101",
97562=>"000000110",
97563=>"000000101",
97564=>"101100111",
97565=>"100001110",
97566=>"011000000",
97567=>"101101111",
97568=>"010000001",
97569=>"001111000",
97570=>"000010000",
97571=>"101001111",
97572=>"011001001",
97573=>"011101111",
97574=>"101000111",
97575=>"000010010",
97576=>"100100111",
97577=>"101100111",
97578=>"010111000",
97579=>"011011000",
97580=>"110111011",
97581=>"000000110",
97582=>"110110110",
97583=>"111001111",
97584=>"100100111",
97585=>"001001100",
97586=>"100000000",
97587=>"101000011",
97588=>"011011011",
97589=>"101111100",
97590=>"011011100",
97591=>"000111000",
97592=>"100000111",
97593=>"111100110",
97594=>"000101111",
97595=>"000000111",
97596=>"111010111",
97597=>"010011110",
97598=>"000000000",
97599=>"101001001",
97600=>"001011111",
97601=>"010110010",
97602=>"100000111",
97603=>"100000110",
97604=>"000000000",
97605=>"000100000",
97606=>"000111000",
97607=>"101000101",
97608=>"000001101",
97609=>"011011010",
97610=>"111100111",
97611=>"011100001",
97612=>"111101111",
97613=>"100111111",
97614=>"000110110",
97615=>"111111111",
97616=>"011010111",
97617=>"010000010",
97618=>"101000100",
97619=>"011001000",
97620=>"011000000",
97621=>"001100100",
97622=>"100110110",
97623=>"000011111",
97624=>"001101101",
97625=>"100001110",
97626=>"110110110",
97627=>"000001000",
97628=>"000000001",
97629=>"000001001",
97630=>"101101101",
97631=>"110110001",
97632=>"011001111",
97633=>"000000010",
97634=>"101100101",
97635=>"011001010",
97636=>"101000110",
97637=>"001001000",
97638=>"011110111",
97639=>"110110111",
97640=>"000100110",
97641=>"000100100",
97642=>"111111111",
97643=>"101111111",
97644=>"000000000",
97645=>"011111001",
97646=>"000000000",
97647=>"011100011",
97648=>"011001000",
97649=>"000000010",
97650=>"111111000",
97651=>"010011111",
97652=>"111111000",
97653=>"000000001",
97654=>"001100111",
97655=>"111011100",
97656=>"001011010",
97657=>"100101010",
97658=>"101010111",
97659=>"111101111",
97660=>"110110010",
97661=>"110100000",
97662=>"010111000",
97663=>"111101100",
97664=>"001011000",
97665=>"000110110",
97666=>"111000111",
97667=>"100101110",
97668=>"111111111",
97669=>"000000001",
97670=>"011111001",
97671=>"001011000",
97672=>"101101000",
97673=>"001010000",
97674=>"000111010",
97675=>"010000000",
97676=>"110100100",
97677=>"000111000",
97678=>"000111001",
97679=>"100000000",
97680=>"100100011",
97681=>"111000011",
97682=>"010011110",
97683=>"011111000",
97684=>"000001000",
97685=>"100000111",
97686=>"111111010",
97687=>"110000000",
97688=>"001111111",
97689=>"000011110",
97690=>"101100111",
97691=>"110100110",
97692=>"000000100",
97693=>"000000111",
97694=>"010011010",
97695=>"001001111",
97696=>"101100101",
97697=>"000101001",
97698=>"111100110",
97699=>"111101000",
97700=>"100000000",
97701=>"100111000",
97702=>"111010000",
97703=>"000100100",
97704=>"001000111",
97705=>"111010010",
97706=>"101100111",
97707=>"000000000",
97708=>"100100011",
97709=>"101000000",
97710=>"010010010",
97711=>"111010000",
97712=>"100000000",
97713=>"010010001",
97714=>"011010000",
97715=>"100010100",
97716=>"000111111",
97717=>"111011000",
97718=>"010010010",
97719=>"010111101",
97720=>"101111111",
97721=>"100011000",
97722=>"000111011",
97723=>"010111011",
97724=>"110010011",
97725=>"011111111",
97726=>"001000110",
97727=>"010010011",
97728=>"000000000",
97729=>"010011000",
97730=>"000111010",
97731=>"100100100",
97732=>"010010000",
97733=>"110100101",
97734=>"000011011",
97735=>"000000001",
97736=>"010100101",
97737=>"110011000",
97738=>"111111111",
97739=>"011000000",
97740=>"000001001",
97741=>"000011000",
97742=>"001001000",
97743=>"111000000",
97744=>"001000000",
97745=>"001001011",
97746=>"110010111",
97747=>"001001000",
97748=>"001000000",
97749=>"110110111",
97750=>"101000100",
97751=>"110000000",
97752=>"010000000",
97753=>"111111111",
97754=>"010010011",
97755=>"111010000",
97756=>"100100100",
97757=>"110000000",
97758=>"100000000",
97759=>"011001000",
97760=>"111000011",
97761=>"111000111",
97762=>"111111000",
97763=>"111110110",
97764=>"000000111",
97765=>"000010111",
97766=>"000000000",
97767=>"011001110",
97768=>"001111111",
97769=>"000110100",
97770=>"011111100",
97771=>"000011010",
97772=>"101101111",
97773=>"111000011",
97774=>"000000000",
97775=>"101100111",
97776=>"100100101",
97777=>"011001001",
97778=>"010000011",
97779=>"100110000",
97780=>"110110000",
97781=>"001101100",
97782=>"000000011",
97783=>"000000000",
97784=>"010010000",
97785=>"010010101",
97786=>"011100001",
97787=>"001011110",
97788=>"001000000",
97789=>"100000100",
97790=>"000000001",
97791=>"110101111",
97792=>"001011011",
97793=>"111110000",
97794=>"001000000",
97795=>"111000000",
97796=>"001111011",
97797=>"101011011",
97798=>"001111100",
97799=>"000111111",
97800=>"000001001",
97801=>"100101101",
97802=>"110100100",
97803=>"000000000",
97804=>"001000000",
97805=>"000011000",
97806=>"100100000",
97807=>"111010011",
97808=>"101000111",
97809=>"000000010",
97810=>"111001000",
97811=>"111110000",
97812=>"111010010",
97813=>"010000000",
97814=>"001001000",
97815=>"000000111",
97816=>"101111110",
97817=>"010100111",
97818=>"000100010",
97819=>"000000000",
97820=>"100110011",
97821=>"110111100",
97822=>"011000000",
97823=>"010001101",
97824=>"000111111",
97825=>"101001100",
97826=>"010001001",
97827=>"000011111",
97828=>"000001111",
97829=>"100000110",
97830=>"100111010",
97831=>"000010110",
97832=>"000010010",
97833=>"111111110",
97834=>"111101101",
97835=>"111100000",
97836=>"111100000",
97837=>"001001001",
97838=>"000000000",
97839=>"001000100",
97840=>"001101111",
97841=>"000000000",
97842=>"111111000",
97843=>"111111110",
97844=>"000000000",
97845=>"111111101",
97846=>"110000000",
97847=>"110101101",
97848=>"101000000",
97849=>"000111000",
97850=>"010011001",
97851=>"010110111",
97852=>"000000000",
97853=>"111111001",
97854=>"000010000",
97855=>"001001011",
97856=>"001000000",
97857=>"111011110",
97858=>"111010111",
97859=>"001001111",
97860=>"111001001",
97861=>"001001100",
97862=>"010010001",
97863=>"000111011",
97864=>"000001100",
97865=>"000001101",
97866=>"000100101",
97867=>"010000000",
97868=>"000001101",
97869=>"000100101",
97870=>"000110100",
97871=>"111000010",
97872=>"111001101",
97873=>"010111111",
97874=>"000011000",
97875=>"001011011",
97876=>"110111000",
97877=>"000000000",
97878=>"100101010",
97879=>"101001111",
97880=>"011010101",
97881=>"011101011",
97882=>"111101100",
97883=>"001110010",
97884=>"000000011",
97885=>"010111001",
97886=>"001000010",
97887=>"100100100",
97888=>"111001101",
97889=>"111100000",
97890=>"001001000",
97891=>"110100100",
97892=>"000110111",
97893=>"010010110",
97894=>"000000001",
97895=>"100111010",
97896=>"001010100",
97897=>"000001000",
97898=>"110111000",
97899=>"100000000",
97900=>"111111000",
97901=>"111111110",
97902=>"011111111",
97903=>"010000000",
97904=>"000010111",
97905=>"011111111",
97906=>"011001001",
97907=>"101101110",
97908=>"100100010",
97909=>"000000000",
97910=>"111000000",
97911=>"000000101",
97912=>"110101111",
97913=>"010000000",
97914=>"111101001",
97915=>"000000011",
97916=>"011001000",
97917=>"100100100",
97918=>"111111111",
97919=>"111110010",
97920=>"110100111",
97921=>"100111000",
97922=>"010000000",
97923=>"111100100",
97924=>"101111110",
97925=>"111110010",
97926=>"011000011",
97927=>"011111011",
97928=>"100101011",
97929=>"000000010",
97930=>"011111111",
97931=>"000000001",
97932=>"000011111",
97933=>"111100101",
97934=>"000011111",
97935=>"110000000",
97936=>"001011001",
97937=>"000000000",
97938=>"001001011",
97939=>"111111000",
97940=>"000000010",
97941=>"000101101",
97942=>"111011000",
97943=>"000000001",
97944=>"010011111",
97945=>"000000000",
97946=>"111111010",
97947=>"111111001",
97948=>"010111000",
97949=>"100111000",
97950=>"001111101",
97951=>"110110000",
97952=>"001011001",
97953=>"110111111",
97954=>"111101101",
97955=>"010000111",
97956=>"000111111",
97957=>"100111011",
97958=>"011011110",
97959=>"110111111",
97960=>"011000110",
97961=>"001000110",
97962=>"101100000",
97963=>"111111111",
97964=>"111010100",
97965=>"101001100",
97966=>"110110100",
97967=>"101010011",
97968=>"001001111",
97969=>"011111001",
97970=>"001111101",
97971=>"000001000",
97972=>"011101111",
97973=>"111111111",
97974=>"000000101",
97975=>"000001000",
97976=>"000000100",
97977=>"010010110",
97978=>"000000010",
97979=>"001000001",
97980=>"111000000",
97981=>"111111111",
97982=>"100100100",
97983=>"111100001",
97984=>"111010011",
97985=>"000000010",
97986=>"110000100",
97987=>"001001000",
97988=>"000000011",
97989=>"100100001",
97990=>"001000000",
97991=>"000000000",
97992=>"111111110",
97993=>"000000010",
97994=>"000110101",
97995=>"100100110",
97996=>"000100111",
97997=>"110100001",
97998=>"111111000",
97999=>"000001111",
98000=>"000000000",
98001=>"001000011",
98002=>"011111110",
98003=>"111100101",
98004=>"011000110",
98005=>"111111100",
98006=>"111111000",
98007=>"010111010",
98008=>"001111111",
98009=>"000000000",
98010=>"100101000",
98011=>"001000110",
98012=>"011000000",
98013=>"100000000",
98014=>"010110000",
98015=>"000000101",
98016=>"010111111",
98017=>"110000000",
98018=>"010010111",
98019=>"011011111",
98020=>"000110000",
98021=>"000000000",
98022=>"000000100",
98023=>"111111011",
98024=>"000101111",
98025=>"111010000",
98026=>"011011011",
98027=>"101011111",
98028=>"000000000",
98029=>"000011011",
98030=>"101111000",
98031=>"001000101",
98032=>"000110011",
98033=>"001001101",
98034=>"010000000",
98035=>"110000000",
98036=>"100110110",
98037=>"011010110",
98038=>"010000010",
98039=>"010000100",
98040=>"000000111",
98041=>"111111011",
98042=>"101111001",
98043=>"110111001",
98044=>"110000000",
98045=>"111101000",
98046=>"000111100",
98047=>"000010100",
98048=>"111101000",
98049=>"110001110",
98050=>"000000111",
98051=>"101001111",
98052=>"111101010",
98053=>"100000000",
98054=>"000000000",
98055=>"000001000",
98056=>"000110000",
98057=>"000010110",
98058=>"000000110",
98059=>"000000000",
98060=>"011000000",
98061=>"111011010",
98062=>"100111010",
98063=>"000000000",
98064=>"001111000",
98065=>"000110110",
98066=>"111111000",
98067=>"000000000",
98068=>"011111000",
98069=>"111111111",
98070=>"100100001",
98071=>"111011111",
98072=>"001000011",
98073=>"110111111",
98074=>"111111010",
98075=>"000000011",
98076=>"101111011",
98077=>"111010110",
98078=>"001111000",
98079=>"011101000",
98080=>"010000000",
98081=>"111110000",
98082=>"001000000",
98083=>"000000000",
98084=>"001001000",
98085=>"001101100",
98086=>"110110100",
98087=>"001001000",
98088=>"000000111",
98089=>"001000101",
98090=>"001110110",
98091=>"000111111",
98092=>"010011011",
98093=>"000110010",
98094=>"111111111",
98095=>"101000101",
98096=>"000011111",
98097=>"000000001",
98098=>"111111000",
98099=>"000010111",
98100=>"000000111",
98101=>"000000000",
98102=>"000111011",
98103=>"001000000",
98104=>"111111000",
98105=>"111101001",
98106=>"000111100",
98107=>"000000001",
98108=>"111111111",
98109=>"101111001",
98110=>"000000000",
98111=>"101110110",
98112=>"111111111",
98113=>"101111110",
98114=>"111000000",
98115=>"011111111",
98116=>"000000000",
98117=>"111100011",
98118=>"011000000",
98119=>"000000101",
98120=>"010111001",
98121=>"111111111",
98122=>"111001001",
98123=>"110110000",
98124=>"111111000",
98125=>"000010110",
98126=>"010001000",
98127=>"111111111",
98128=>"111111111",
98129=>"110110010",
98130=>"001000111",
98131=>"001010000",
98132=>"000000011",
98133=>"110111110",
98134=>"001001000",
98135=>"111111111",
98136=>"000000100",
98137=>"001000001",
98138=>"111001000",
98139=>"011010000",
98140=>"111111000",
98141=>"111101001",
98142=>"001000001",
98143=>"010011011",
98144=>"010110010",
98145=>"010111011",
98146=>"110100110",
98147=>"001100100",
98148=>"111101000",
98149=>"111111001",
98150=>"111111000",
98151=>"000011111",
98152=>"101101000",
98153=>"011000010",
98154=>"010000101",
98155=>"111111000",
98156=>"111111111",
98157=>"000000000",
98158=>"111001111",
98159=>"110010000",
98160=>"110100000",
98161=>"100111111",
98162=>"000111110",
98163=>"000000011",
98164=>"111000000",
98165=>"000000000",
98166=>"110111110",
98167=>"111010000",
98168=>"000000111",
98169=>"111000000",
98170=>"100000000",
98171=>"000000000",
98172=>"111111111",
98173=>"110100000",
98174=>"111111111",
98175=>"011110110",
98176=>"101111010",
98177=>"110100000",
98178=>"011011010",
98179=>"011001000",
98180=>"000000000",
98181=>"101010000",
98182=>"000111000",
98183=>"110110110",
98184=>"111111111",
98185=>"111101000",
98186=>"101011011",
98187=>"101100101",
98188=>"000000000",
98189=>"111111110",
98190=>"001111110",
98191=>"000000011",
98192=>"101111001",
98193=>"111011000",
98194=>"000000000",
98195=>"100110000",
98196=>"110111110",
98197=>"100111111",
98198=>"100001000",
98199=>"010000000",
98200=>"000000010",
98201=>"010111010",
98202=>"100111111",
98203=>"000000000",
98204=>"110100001",
98205=>"000000111",
98206=>"111000000",
98207=>"000000010",
98208=>"111111101",
98209=>"111111111",
98210=>"111111111",
98211=>"001000111",
98212=>"010110011",
98213=>"110110010",
98214=>"000000000",
98215=>"011111111",
98216=>"000000111",
98217=>"110000111",
98218=>"001000101",
98219=>"000000110",
98220=>"111111111",
98221=>"111010110",
98222=>"111101001",
98223=>"000000001",
98224=>"111000000",
98225=>"111001001",
98226=>"011011011",
98227=>"101011000",
98228=>"111011110",
98229=>"111111111",
98230=>"111101001",
98231=>"001110101",
98232=>"011111101",
98233=>"111111111",
98234=>"110100111",
98235=>"010010111",
98236=>"000000000",
98237=>"111111110",
98238=>"011001100",
98239=>"110001111",
98240=>"000011111",
98241=>"111011011",
98242=>"111110101",
98243=>"111011110",
98244=>"011000000",
98245=>"111000100",
98246=>"000000100",
98247=>"011011000",
98248=>"000000100",
98249=>"111001000",
98250=>"101001111",
98251=>"111111011",
98252=>"001111011",
98253=>"011011101",
98254=>"000000110",
98255=>"000011000",
98256=>"000000010",
98257=>"100110000",
98258=>"100000111",
98259=>"001100000",
98260=>"000000001",
98261=>"100000000",
98262=>"000000000",
98263=>"010000000",
98264=>"000000000",
98265=>"100010000",
98266=>"000011010",
98267=>"001000110",
98268=>"001010000",
98269=>"011011011",
98270=>"000000111",
98271=>"101000010",
98272=>"110111111",
98273=>"000000111",
98274=>"000000000",
98275=>"111111000",
98276=>"000000000",
98277=>"000000000",
98278=>"000000000",
98279=>"011111010",
98280=>"101000001",
98281=>"000000000",
98282=>"000001111",
98283=>"111001000",
98284=>"111000000",
98285=>"001000010",
98286=>"000010000",
98287=>"010000000",
98288=>"000000000",
98289=>"111001001",
98290=>"110111111",
98291=>"010100000",
98292=>"100011000",
98293=>"101101111",
98294=>"010110010",
98295=>"000000111",
98296=>"010110000",
98297=>"111000000",
98298=>"000001111",
98299=>"111011000",
98300=>"110010000",
98301=>"101101111",
98302=>"111100000",
98303=>"001111111",
98304=>"000100100",
98305=>"100111110",
98306=>"100100111",
98307=>"000000011",
98308=>"011111100",
98309=>"000001000",
98310=>"100100000",
98311=>"001011011",
98312=>"011011001",
98313=>"000011011",
98314=>"000000000",
98315=>"000100011",
98316=>"001011100",
98317=>"100100111",
98318=>"100001011",
98319=>"110001011",
98320=>"111010000",
98321=>"000000000",
98322=>"110110010",
98323=>"111000000",
98324=>"100100011",
98325=>"000000000",
98326=>"110111111",
98327=>"111011010",
98328=>"001111001",
98329=>"111101100",
98330=>"001011000",
98331=>"000100110",
98332=>"000010001",
98333=>"100110110",
98334=>"100000000",
98335=>"111110100",
98336=>"011011010",
98337=>"011001101",
98338=>"110000000",
98339=>"001011000",
98340=>"001111111",
98341=>"011111110",
98342=>"010011011",
98343=>"000001000",
98344=>"100100111",
98345=>"010100110",
98346=>"110000100",
98347=>"110100111",
98348=>"000001001",
98349=>"100011001",
98350=>"100110011",
98351=>"111011011",
98352=>"011010010",
98353=>"100111011",
98354=>"011011011",
98355=>"110100000",
98356=>"100100110",
98357=>"101111010",
98358=>"110100011",
98359=>"011000011",
98360=>"011110011",
98361=>"000000011",
98362=>"000000000",
98363=>"100110000",
98364=>"011111111",
98365=>"011111100",
98366=>"100000111",
98367=>"001011001",
98368=>"011000000",
98369=>"011010000",
98370=>"011011001",
98371=>"011100100",
98372=>"110101101",
98373=>"100000000",
98374=>"000011010",
98375=>"001011111",
98376=>"010010011",
98377=>"001011010",
98378=>"011100111",
98379=>"000011110",
98380=>"100000000",
98381=>"110110011",
98382=>"111100011",
98383=>"111011011",
98384=>"010000111",
98385=>"110110111",
98386=>"110111011",
98387=>"001000010",
98388=>"100100110",
98389=>"100000000",
98390=>"001001001",
98391=>"110100011",
98392=>"011100111",
98393=>"010011011",
98394=>"111001010",
98395=>"010101111",
98396=>"011011000",
98397=>"001000001",
98398=>"110100110",
98399=>"000100000",
98400=>"011011000",
98401=>"011001011",
98402=>"000111111",
98403=>"011100111",
98404=>"110110111",
98405=>"011111011",
98406=>"010000000",
98407=>"111111011",
98408=>"010011011",
98409=>"001100000",
98410=>"011011011",
98411=>"000110100",
98412=>"001111000",
98413=>"100100111",
98414=>"000010010",
98415=>"001011011",
98416=>"000001010",
98417=>"011011011",
98418=>"000000110",
98419=>"100011000",
98420=>"000001011",
98421=>"010000000",
98422=>"000010011",
98423=>"000100100",
98424=>"101000011",
98425=>"111110110",
98426=>"111100100",
98427=>"100101101",
98428=>"011011011",
98429=>"110110000",
98430=>"000100011",
98431=>"000000110",
98432=>"011000000",
98433=>"110100110",
98434=>"011011010",
98435=>"000100011",
98436=>"011011011",
98437=>"101010000",
98438=>"010001001",
98439=>"111101000",
98440=>"111011000",
98441=>"000000000",
98442=>"100100000",
98443=>"001100000",
98444=>"100100110",
98445=>"000100101",
98446=>"011000000",
98447=>"111000010",
98448=>"101111000",
98449=>"000110100",
98450=>"000001011",
98451=>"011010000",
98452=>"001011001",
98453=>"100100100",
98454=>"011011000",
98455=>"010001001",
98456=>"011011000",
98457=>"000011011",
98458=>"011011101",
98459=>"011011011",
98460=>"001110000",
98461=>"011010111",
98462=>"011011000",
98463=>"101011001",
98464=>"000000000",
98465=>"000100111",
98466=>"010111000",
98467=>"111110111",
98468=>"011111100",
98469=>"001011000",
98470=>"111001000",
98471=>"001011000",
98472=>"100011011",
98473=>"000011011",
98474=>"001000110",
98475=>"001000100",
98476=>"111000100",
98477=>"011001011",
98478=>"010110111",
98479=>"011111011",
98480=>"011011010",
98481=>"101100100",
98482=>"111100111",
98483=>"100110111",
98484=>"010011110",
98485=>"110000100",
98486=>"011010001",
98487=>"111101110",
98488=>"011011011",
98489=>"001011000",
98490=>"001000000",
98491=>"000001010",
98492=>"101010000",
98493=>"110111111",
98494=>"011011010",
98495=>"100100001",
98496=>"100100111",
98497=>"100100110",
98498=>"011010001",
98499=>"100111100",
98500=>"000000000",
98501=>"101110000",
98502=>"111110100",
98503=>"010111111",
98504=>"001001011",
98505=>"100100100",
98506=>"111111111",
98507=>"000100111",
98508=>"000001010",
98509=>"000100011",
98510=>"100000110",
98511=>"011111011",
98512=>"000000011",
98513=>"111011001",
98514=>"011011001",
98515=>"100001011",
98516=>"011011000",
98517=>"111010101",
98518=>"010000011",
98519=>"001011011",
98520=>"111110000",
98521=>"100100000",
98522=>"100110110",
98523=>"100100100",
98524=>"111101011",
98525=>"110100100",
98526=>"110001000",
98527=>"100100110",
98528=>"100000010",
98529=>"100100111",
98530=>"000000010",
98531=>"101111001",
98532=>"111100111",
98533=>"100100100",
98534=>"001000001",
98535=>"001010011",
98536=>"000011001",
98537=>"110111111",
98538=>"010000000",
98539=>"000100111",
98540=>"000100110",
98541=>"000000011",
98542=>"110100100",
98543=>"011010000",
98544=>"101010000",
98545=>"110110111",
98546=>"000000011",
98547=>"100100111",
98548=>"010000011",
98549=>"111001101",
98550=>"000011011",
98551=>"011000110",
98552=>"100100111",
98553=>"010000000",
98554=>"110110111",
98555=>"101111001",
98556=>"011011000",
98557=>"011110110",
98558=>"011011000",
98559=>"011011011",
98560=>"010000000",
98561=>"011011010",
98562=>"000000111",
98563=>"001000010",
98564=>"100001001",
98565=>"000100111",
98566=>"001111011",
98567=>"000011010",
98568=>"010000111",
98569=>"111011101",
98570=>"011001111",
98571=>"001000111",
98572=>"000000111",
98573=>"000001010",
98574=>"101011010",
98575=>"110111000",
98576=>"111011010",
98577=>"000000000",
98578=>"101000000",
98579=>"010000000",
98580=>"011111001",
98581=>"000000100",
98582=>"000000100",
98583=>"100011110",
98584=>"010001111",
98585=>"101111010",
98586=>"000101011",
98587=>"100000110",
98588=>"111111001",
98589=>"000111111",
98590=>"000000010",
98591=>"000100100",
98592=>"111000000",
98593=>"010010011",
98594=>"111100100",
98595=>"111110010",
98596=>"000110000",
98597=>"010110000",
98598=>"011000010",
98599=>"000011011",
98600=>"000000000",
98601=>"000111011",
98602=>"111011010",
98603=>"001100000",
98604=>"011001011",
98605=>"111000010",
98606=>"000001010",
98607=>"100111110",
98608=>"000000000",
98609=>"000000001",
98610=>"000101100",
98611=>"010000000",
98612=>"000000101",
98613=>"101000111",
98614=>"110010010",
98615=>"111010000",
98616=>"011010000",
98617=>"001001000",
98618=>"000100001",
98619=>"000000000",
98620=>"000000000",
98621=>"111101110",
98622=>"001100100",
98623=>"011011101",
98624=>"100101111",
98625=>"111111101",
98626=>"000000101",
98627=>"000000010",
98628=>"101101001",
98629=>"000000100",
98630=>"000000001",
98631=>"010111000",
98632=>"100001001",
98633=>"110111100",
98634=>"110000001",
98635=>"000010001",
98636=>"000000000",
98637=>"110111111",
98638=>"011100110",
98639=>"010110100",
98640=>"010000101",
98641=>"111000011",
98642=>"011011101",
98643=>"000001100",
98644=>"000010010",
98645=>"100110100",
98646=>"100111110",
98647=>"011000111",
98648=>"000001101",
98649=>"000001001",
98650=>"000111001",
98651=>"011011100",
98652=>"011010110",
98653=>"000001000",
98654=>"111111111",
98655=>"000100111",
98656=>"111101111",
98657=>"000101011",
98658=>"101000111",
98659=>"000100100",
98660=>"100010000",
98661=>"100001111",
98662=>"110100110",
98663=>"111000100",
98664=>"101001101",
98665=>"010000111",
98666=>"101011111",
98667=>"110001101",
98668=>"000000000",
98669=>"001010010",
98670=>"000000011",
98671=>"000001000",
98672=>"001100000",
98673=>"000001010",
98674=>"011011011",
98675=>"000000111",
98676=>"111101001",
98677=>"001000101",
98678=>"101001010",
98679=>"111100100",
98680=>"001000011",
98681=>"111111011",
98682=>"111111010",
98683=>"000101111",
98684=>"100110110",
98685=>"000100001",
98686=>"100101101",
98687=>"000100101",
98688=>"010011000",
98689=>"000000000",
98690=>"010000001",
98691=>"101111110",
98692=>"000000111",
98693=>"001101010",
98694=>"010011000",
98695=>"001011011",
98696=>"000100010",
98697=>"000000010",
98698=>"111011111",
98699=>"000000111",
98700=>"101000000",
98701=>"011111111",
98702=>"000000000",
98703=>"001000100",
98704=>"001001101",
98705=>"111111000",
98706=>"011011000",
98707=>"000000111",
98708=>"100011110",
98709=>"000000010",
98710=>"111011010",
98711=>"000111000",
98712=>"110010100",
98713=>"011111111",
98714=>"111100111",
98715=>"011001001",
98716=>"111101101",
98717=>"101101111",
98718=>"010011111",
98719=>"000111111",
98720=>"101011101",
98721=>"111000000",
98722=>"000010000",
98723=>"010000101",
98724=>"000111111",
98725=>"110110000",
98726=>"111110001",
98727=>"011101010",
98728=>"000000010",
98729=>"111000000",
98730=>"101101111",
98731=>"000000000",
98732=>"101111010",
98733=>"100000101",
98734=>"110110000",
98735=>"111111111",
98736=>"000101010",
98737=>"001101111",
98738=>"101101111",
98739=>"100100010",
98740=>"010110001",
98741=>"100100111",
98742=>"001011000",
98743=>"111011101",
98744=>"100100001",
98745=>"000110111",
98746=>"110000000",
98747=>"011011000",
98748=>"010111001",
98749=>"001111111",
98750=>"100100101",
98751=>"000000010",
98752=>"000000100",
98753=>"101001110",
98754=>"101111010",
98755=>"000000011",
98756=>"010011000",
98757=>"110110010",
98758=>"100011011",
98759=>"011111100",
98760=>"000111011",
98761=>"010111000",
98762=>"111111000",
98763=>"000110100",
98764=>"101000001",
98765=>"100011011",
98766=>"101111010",
98767=>"111000000",
98768=>"111101111",
98769=>"011111110",
98770=>"101010010",
98771=>"000000111",
98772=>"001000011",
98773=>"100001000",
98774=>"010101011",
98775=>"000000100",
98776=>"000000010",
98777=>"111101000",
98778=>"011111110",
98779=>"001000001",
98780=>"000000010",
98781=>"111001101",
98782=>"001000001",
98783=>"000001010",
98784=>"101000101",
98785=>"000000011",
98786=>"001100100",
98787=>"111111011",
98788=>"100000100",
98789=>"101101000",
98790=>"110000000",
98791=>"111011000",
98792=>"011101010",
98793=>"111111110",
98794=>"110011011",
98795=>"100000101",
98796=>"000100000",
98797=>"010001010",
98798=>"010000010",
98799=>"010100000",
98800=>"000010000",
98801=>"001011111",
98802=>"111000110",
98803=>"001101101",
98804=>"110001001",
98805=>"111111111",
98806=>"000000011",
98807=>"011101011",
98808=>"010010000",
98809=>"001001100",
98810=>"000111110",
98811=>"000111111",
98812=>"000000000",
98813=>"010011000",
98814=>"000001011",
98815=>"101000100",
98816=>"000000000",
98817=>"010010010",
98818=>"100001001",
98819=>"010011110",
98820=>"100111011",
98821=>"111110100",
98822=>"100111101",
98823=>"000100111",
98824=>"000000100",
98825=>"000001000",
98826=>"000000010",
98827=>"111110100",
98828=>"101110100",
98829=>"101110101",
98830=>"111111111",
98831=>"111111111",
98832=>"001101011",
98833=>"000011010",
98834=>"000010000",
98835=>"111011110",
98836=>"110111111",
98837=>"000000011",
98838=>"000000110",
98839=>"111110010",
98840=>"101001001",
98841=>"101101100",
98842=>"100000110",
98843=>"000011011",
98844=>"110111011",
98845=>"100010000",
98846=>"110110010",
98847=>"000000000",
98848=>"000001011",
98849=>"110110101",
98850=>"100100001",
98851=>"000000000",
98852=>"111110000",
98853=>"011110000",
98854=>"000001010",
98855=>"011110110",
98856=>"000000100",
98857=>"000010110",
98858=>"000100110",
98859=>"100100000",
98860=>"011111100",
98861=>"011000000",
98862=>"111100000",
98863=>"100100001",
98864=>"110100100",
98865=>"000111111",
98866=>"100100101",
98867=>"100100000",
98868=>"000001011",
98869=>"001001011",
98870=>"011110100",
98871=>"111111110",
98872=>"110100100",
98873=>"100011010",
98874=>"100001011",
98875=>"010100000",
98876=>"001001000",
98877=>"001111111",
98878=>"000000001",
98879=>"010100000",
98880=>"011111001",
98881=>"100100100",
98882=>"110111111",
98883=>"000000000",
98884=>"111001000",
98885=>"000000000",
98886=>"001100110",
98887=>"111101100",
98888=>"101101100",
98889=>"010111111",
98890=>"100000000",
98891=>"100000001",
98892=>"100101000",
98893=>"001011011",
98894=>"011010000",
98895=>"000011001",
98896=>"100111000",
98897=>"110010011",
98898=>"011100001",
98899=>"000000000",
98900=>"111111001",
98901=>"001101000",
98902=>"000100100",
98903=>"000011011",
98904=>"111111111",
98905=>"001111111",
98906=>"001011000",
98907=>"000100101",
98908=>"000001111",
98909=>"001001011",
98910=>"111000011",
98911=>"111100111",
98912=>"111110100",
98913=>"011011011",
98914=>"100000011",
98915=>"110011011",
98916=>"000000000",
98917=>"010110100",
98918=>"011101100",
98919=>"111101110",
98920=>"111111100",
98921=>"011111110",
98922=>"011110110",
98923=>"111011111",
98924=>"000100000",
98925=>"000001011",
98926=>"000000001",
98927=>"011011011",
98928=>"011011010",
98929=>"011110010",
98930=>"000000000",
98931=>"000100000",
98932=>"111111111",
98933=>"000010000",
98934=>"000001011",
98935=>"001011010",
98936=>"100000000",
98937=>"111111100",
98938=>"110100100",
98939=>"010000000",
98940=>"000000000",
98941=>"111111100",
98942=>"111110000",
98943=>"101001011",
98944=>"110100110",
98945=>"100110100",
98946=>"000110110",
98947=>"001100001",
98948=>"111100000",
98949=>"001100000",
98950=>"110110010",
98951=>"000011011",
98952=>"001111101",
98953=>"100000001",
98954=>"001100100",
98955=>"101100001",
98956=>"101011000",
98957=>"100100001",
98958=>"101001111",
98959=>"001001001",
98960=>"000010000",
98961=>"001011011",
98962=>"000000000",
98963=>"011001011",
98964=>"011011000",
98965=>"100001011",
98966=>"001011000",
98967=>"100000111",
98968=>"000110100",
98969=>"100000011",
98970=>"111001001",
98971=>"000000011",
98972=>"001011011",
98973=>"110111111",
98974=>"000010001",
98975=>"000001001",
98976=>"000010101",
98977=>"110000011",
98978=>"001000101",
98979=>"111001000",
98980=>"111110100",
98981=>"111101010",
98982=>"001000010",
98983=>"011110100",
98984=>"000000000",
98985=>"001000001",
98986=>"111000001",
98987=>"000000001",
98988=>"001001000",
98989=>"100010000",
98990=>"111111111",
98991=>"001010011",
98992=>"000000110",
98993=>"000000000",
98994=>"110000000",
98995=>"000000000",
98996=>"000111100",
98997=>"011101000",
98998=>"001101101",
98999=>"001100101",
99000=>"000100100",
99001=>"000000110",
99002=>"111101011",
99003=>"010111010",
99004=>"000000100",
99005=>"111110100",
99006=>"000000100",
99007=>"000000001",
99008=>"000001010",
99009=>"000001011",
99010=>"010110111",
99011=>"011111100",
99012=>"001000000",
99013=>"010000001",
99014=>"111111111",
99015=>"100110110",
99016=>"000000101",
99017=>"101001001",
99018=>"111010001",
99019=>"001011000",
99020=>"001011011",
99021=>"111011111",
99022=>"000000001",
99023=>"011110001",
99024=>"000110100",
99025=>"011010000",
99026=>"001001001",
99027=>"111110100",
99028=>"100000001",
99029=>"001011110",
99030=>"110000010",
99031=>"101111110",
99032=>"101110100",
99033=>"001000100",
99034=>"111000000",
99035=>"110001011",
99036=>"111110000",
99037=>"101001010",
99038=>"001010000",
99039=>"011110000",
99040=>"000001001",
99041=>"000001001",
99042=>"111000100",
99043=>"000001001",
99044=>"000000000",
99045=>"000001000",
99046=>"001111100",
99047=>"000000000",
99048=>"000110110",
99049=>"000000000",
99050=>"010111111",
99051=>"000000110",
99052=>"000011110",
99053=>"111001001",
99054=>"000000000",
99055=>"000000100",
99056=>"000100100",
99057=>"000111111",
99058=>"110000110",
99059=>"010000000",
99060=>"111111111",
99061=>"100100000",
99062=>"100001101",
99063=>"011110101",
99064=>"110010010",
99065=>"111111111",
99066=>"100101011",
99067=>"000010100",
99068=>"111111110",
99069=>"000000110",
99070=>"011111111",
99071=>"110110110",
99072=>"100110110",
99073=>"001101101",
99074=>"111010000",
99075=>"000000000",
99076=>"001001000",
99077=>"101111111",
99078=>"111010000",
99079=>"111000011",
99080=>"001001001",
99081=>"101000000",
99082=>"110100110",
99083=>"111111001",
99084=>"111111100",
99085=>"111001000",
99086=>"010000000",
99087=>"110010011",
99088=>"100101011",
99089=>"000000000",
99090=>"000000000",
99091=>"111101101",
99092=>"111110000",
99093=>"111111000",
99094=>"000000001",
99095=>"110110010",
99096=>"111111111",
99097=>"000101111",
99098=>"111111111",
99099=>"111111000",
99100=>"001100000",
99101=>"011000001",
99102=>"001000010",
99103=>"000000000",
99104=>"111111111",
99105=>"111010111",
99106=>"000000000",
99107=>"111111101",
99108=>"001000000",
99109=>"111111111",
99110=>"111010000",
99111=>"000100011",
99112=>"000011000",
99113=>"111101111",
99114=>"000000000",
99115=>"111111111",
99116=>"111111001",
99117=>"111111111",
99118=>"000100111",
99119=>"001000001",
99120=>"100000111",
99121=>"000000000",
99122=>"010010111",
99123=>"010111111",
99124=>"011001000",
99125=>"111101101",
99126=>"100000000",
99127=>"010110110",
99128=>"000000100",
99129=>"111111000",
99130=>"000000000",
99131=>"001000110",
99132=>"111011011",
99133=>"111001001",
99134=>"000000001",
99135=>"001001010",
99136=>"111101111",
99137=>"101101110",
99138=>"000000111",
99139=>"100000101",
99140=>"111101110",
99141=>"000000000",
99142=>"011011011",
99143=>"000101111",
99144=>"101111111",
99145=>"110100111",
99146=>"000000000",
99147=>"111101001",
99148=>"100100010",
99149=>"000000000",
99150=>"000000000",
99151=>"111101111",
99152=>"000000000",
99153=>"111010111",
99154=>"011111111",
99155=>"000000000",
99156=>"000101001",
99157=>"000011000",
99158=>"001001000",
99159=>"010000000",
99160=>"001011001",
99161=>"100000000",
99162=>"011001000",
99163=>"000000101",
99164=>"000000000",
99165=>"000000000",
99166=>"111111110",
99167=>"001000000",
99168=>"101101111",
99169=>"111111111",
99170=>"000000110",
99171=>"000000000",
99172=>"000000000",
99173=>"101000001",
99174=>"111111000",
99175=>"011011000",
99176=>"000000000",
99177=>"111010111",
99178=>"000010001",
99179=>"111111111",
99180=>"111111110",
99181=>"111111111",
99182=>"111110111",
99183=>"000011100",
99184=>"000000000",
99185=>"111010111",
99186=>"001000000",
99187=>"111111111",
99188=>"000000111",
99189=>"000000000",
99190=>"110000000",
99191=>"100000111",
99192=>"111111010",
99193=>"101011000",
99194=>"111111011",
99195=>"001000000",
99196=>"011000000",
99197=>"000000000",
99198=>"111111111",
99199=>"001000000",
99200=>"000000011",
99201=>"111000000",
99202=>"111000000",
99203=>"010000000",
99204=>"000001010",
99205=>"110101101",
99206=>"100100111",
99207=>"100100001",
99208=>"000100001",
99209=>"101101101",
99210=>"000000000",
99211=>"000000100",
99212=>"111111110",
99213=>"101011110",
99214=>"000000100",
99215=>"000000000",
99216=>"000000000",
99217=>"010010111",
99218=>"010000111",
99219=>"110111011",
99220=>"010101100",
99221=>"000000000",
99222=>"111111111",
99223=>"000000001",
99224=>"101101101",
99225=>"111111101",
99226=>"010111100",
99227=>"111001111",
99228=>"010111100",
99229=>"111111101",
99230=>"001000001",
99231=>"100000000",
99232=>"100000000",
99233=>"000011000",
99234=>"101000001",
99235=>"111111010",
99236=>"110101101",
99237=>"001001001",
99238=>"000000001",
99239=>"111111110",
99240=>"110000001",
99241=>"110111100",
99242=>"111111000",
99243=>"000010110",
99244=>"011001000",
99245=>"000000000",
99246=>"101110010",
99247=>"110100111",
99248=>"000001010",
99249=>"111101011",
99250=>"000000000",
99251=>"000000000",
99252=>"000100000",
99253=>"111111011",
99254=>"000010000",
99255=>"110110001",
99256=>"100011110",
99257=>"010101101",
99258=>"000111111",
99259=>"011111001",
99260=>"111111111",
99261=>"111000000",
99262=>"001000100",
99263=>"111110111",
99264=>"101110001",
99265=>"101101101",
99266=>"000001000",
99267=>"000000100",
99268=>"010010000",
99269=>"001011111",
99270=>"111101000",
99271=>"110110110",
99272=>"000100000",
99273=>"000000000",
99274=>"000101000",
99275=>"111101111",
99276=>"011101110",
99277=>"110100000",
99278=>"001000000",
99279=>"000000000",
99280=>"000000000",
99281=>"001001001",
99282=>"101110111",
99283=>"000000011",
99284=>"000001111",
99285=>"111001100",
99286=>"111111110",
99287=>"000000111",
99288=>"111111001",
99289=>"111111111",
99290=>"001001001",
99291=>"000000010",
99292=>"000001001",
99293=>"100000000",
99294=>"110101001",
99295=>"111001111",
99296=>"101011111",
99297=>"010001111",
99298=>"000000000",
99299=>"101011011",
99300=>"000000001",
99301=>"111111000",
99302=>"000100000",
99303=>"101111101",
99304=>"000000001",
99305=>"111110111",
99306=>"001001000",
99307=>"111101110",
99308=>"010000000",
99309=>"000000111",
99310=>"000000000",
99311=>"000000110",
99312=>"111111000",
99313=>"100110111",
99314=>"000101101",
99315=>"001001000",
99316=>"001001001",
99317=>"100001011",
99318=>"000000101",
99319=>"000000101",
99320=>"111000110",
99321=>"000000111",
99322=>"111111111",
99323=>"111110111",
99324=>"001001111",
99325=>"111111000",
99326=>"001000001",
99327=>"010000001",
99328=>"100100110",
99329=>"111111000",
99330=>"000010110",
99331=>"111001000",
99332=>"011010000",
99333=>"001111111",
99334=>"111101000",
99335=>"010010000",
99336=>"101111011",
99337=>"001000001",
99338=>"110111111",
99339=>"111001000",
99340=>"000110111",
99341=>"110101001",
99342=>"001011000",
99343=>"000101110",
99344=>"111111000",
99345=>"111000000",
99346=>"110110111",
99347=>"111001000",
99348=>"000110111",
99349=>"000111111",
99350=>"010100000",
99351=>"111000100",
99352=>"010101111",
99353=>"110011111",
99354=>"111000000",
99355=>"111001000",
99356=>"000011000",
99357=>"000001110",
99358=>"000001011",
99359=>"001001111",
99360=>"110000101",
99361=>"001000000",
99362=>"001000000",
99363=>"111111000",
99364=>"100100110",
99365=>"111100000",
99366=>"000010111",
99367=>"000000000",
99368=>"000111111",
99369=>"111001000",
99370=>"000000000",
99371=>"111000101",
99372=>"011100111",
99373=>"110110010",
99374=>"010111111",
99375=>"011111111",
99376=>"101000000",
99377=>"111000010",
99378=>"000110000",
99379=>"000000000",
99380=>"111000000",
99381=>"111111111",
99382=>"110100000",
99383=>"101001001",
99384=>"110110110",
99385=>"111101111",
99386=>"000000000",
99387=>"110000000",
99388=>"001100000",
99389=>"001000001",
99390=>"001100000",
99391=>"011011000",
99392=>"000111111",
99393=>"101111000",
99394=>"111001000",
99395=>"100110111",
99396=>"000000000",
99397=>"000111100",
99398=>"111111000",
99399=>"001111111",
99400=>"101100000",
99401=>"101101001",
99402=>"000110110",
99403=>"011000000",
99404=>"111000000",
99405=>"011011110",
99406=>"111011011",
99407=>"000001111",
99408=>"001001001",
99409=>"111110101",
99410=>"111001000",
99411=>"000010010",
99412=>"011111000",
99413=>"000100000",
99414=>"011001001",
99415=>"010111110",
99416=>"000000001",
99417=>"100000000",
99418=>"000000000",
99419=>"111001001",
99420=>"000000000",
99421=>"000110011",
99422=>"000111111",
99423=>"011111111",
99424=>"111001000",
99425=>"000010110",
99426=>"111000000",
99427=>"001011101",
99428=>"000000010",
99429=>"001001111",
99430=>"111101111",
99431=>"000000010",
99432=>"000000000",
99433=>"000000000",
99434=>"011111001",
99435=>"001011010",
99436=>"111101000",
99437=>"111111111",
99438=>"000000111",
99439=>"110111000",
99440=>"011110100",
99441=>"000000000",
99442=>"111001001",
99443=>"000110000",
99444=>"110000000",
99445=>"110111000",
99446=>"000000000",
99447=>"111111100",
99448=>"000111010",
99449=>"111001000",
99450=>"000000000",
99451=>"010110110",
99452=>"011001000",
99453=>"000011110",
99454=>"000010110",
99455=>"000010111",
99456=>"111101000",
99457=>"111001001",
99458=>"101000000",
99459=>"000000100",
99460=>"000000000",
99461=>"001000001",
99462=>"111011000",
99463=>"101000001",
99464=>"010011001",
99465=>"111001000",
99466=>"000111111",
99467=>"111111000",
99468=>"111000000",
99469=>"001100000",
99470=>"000011100",
99471=>"111011101",
99472=>"010011011",
99473=>"000001000",
99474=>"111000000",
99475=>"110111000",
99476=>"000000010",
99477=>"101001000",
99478=>"110100110",
99479=>"000000000",
99480=>"111001010",
99481=>"000011000",
99482=>"001001011",
99483=>"000111110",
99484=>"111101000",
99485=>"110011101",
99486=>"101011101",
99487=>"111001010",
99488=>"111000111",
99489=>"010011000",
99490=>"000111111",
99491=>"111001001",
99492=>"111100000",
99493=>"110100010",
99494=>"000000111",
99495=>"111101000",
99496=>"111110000",
99497=>"110000000",
99498=>"000011111",
99499=>"110110000",
99500=>"110010110",
99501=>"000100111",
99502=>"000011011",
99503=>"000111111",
99504=>"000000000",
99505=>"111001000",
99506=>"000110000",
99507=>"001001011",
99508=>"110001001",
99509=>"000100000",
99510=>"110000000",
99511=>"001110011",
99512=>"000001001",
99513=>"000000100",
99514=>"101101011",
99515=>"000000010",
99516=>"010111111",
99517=>"111111000",
99518=>"110100000",
99519=>"101000100",
99520=>"000110111",
99521=>"010001001",
99522=>"100000000",
99523=>"111111111",
99524=>"011111110",
99525=>"000100101",
99526=>"000001000",
99527=>"000000101",
99528=>"011111000",
99529=>"111000101",
99530=>"001000000",
99531=>"111010000",
99532=>"011010000",
99533=>"100100001",
99534=>"101001001",
99535=>"011000000",
99536=>"111100101",
99537=>"111010010",
99538=>"100000000",
99539=>"000000000",
99540=>"001111000",
99541=>"110000011",
99542=>"001111111",
99543=>"110111010",
99544=>"000111111",
99545=>"000000000",
99546=>"111101111",
99547=>"111000000",
99548=>"000000001",
99549=>"111101111",
99550=>"000000001",
99551=>"110101001",
99552=>"000111111",
99553=>"001111111",
99554=>"000000010",
99555=>"010110010",
99556=>"000010110",
99557=>"111000000",
99558=>"111011011",
99559=>"001001111",
99560=>"100001000",
99561=>"110110010",
99562=>"110111110",
99563=>"000000000",
99564=>"000111111",
99565=>"011111111",
99566=>"000010000",
99567=>"111000000",
99568=>"000000000",
99569=>"001011000",
99570=>"000001000",
99571=>"000100100",
99572=>"001011000",
99573=>"000001111",
99574=>"100101011",
99575=>"000000110",
99576=>"101111000",
99577=>"111110000",
99578=>"110110101",
99579=>"001001110",
99580=>"000111011",
99581=>"000001000",
99582=>"111101011",
99583=>"010111011",
99584=>"000100110",
99585=>"011101100",
99586=>"000011100",
99587=>"011111101",
99588=>"110001011",
99589=>"111101101",
99590=>"011100101",
99591=>"000010000",
99592=>"101100000",
99593=>"000111101",
99594=>"001000000",
99595=>"101000100",
99596=>"111111111",
99597=>"100101110",
99598=>"110100100",
99599=>"000000000",
99600=>"101100100",
99601=>"101100000",
99602=>"111111011",
99603=>"111101101",
99604=>"000011000",
99605=>"000100000",
99606=>"000000100",
99607=>"111111111",
99608=>"000000101",
99609=>"100001101",
99610=>"000000000",
99611=>"000111110",
99612=>"010011110",
99613=>"001010011",
99614=>"000111101",
99615=>"111111111",
99616=>"000000000",
99617=>"101100000",
99618=>"011111000",
99619=>"101000000",
99620=>"001111010",
99621=>"100000110",
99622=>"000100000",
99623=>"000000000",
99624=>"100111111",
99625=>"000111011",
99626=>"100010010",
99627=>"110111111",
99628=>"100100100",
99629=>"000000000",
99630=>"010010010",
99631=>"001111100",
99632=>"000111111",
99633=>"100000110",
99634=>"111100101",
99635=>"000000100",
99636=>"100000111",
99637=>"000000000",
99638=>"100100001",
99639=>"000100100",
99640=>"011000111",
99641=>"010000000",
99642=>"001111010",
99643=>"111111111",
99644=>"010111010",
99645=>"111101111",
99646=>"100000111",
99647=>"001001001",
99648=>"111110111",
99649=>"110100111",
99650=>"111101000",
99651=>"000000100",
99652=>"100000100",
99653=>"100111111",
99654=>"111111111",
99655=>"111011011",
99656=>"010110101",
99657=>"000010000",
99658=>"001111100",
99659=>"000111111",
99660=>"110100100",
99661=>"010011001",
99662=>"011110100",
99663=>"001100100",
99664=>"000000000",
99665=>"101111111",
99666=>"011111111",
99667=>"010111111",
99668=>"101000000",
99669=>"000101000",
99670=>"000110100",
99671=>"000011111",
99672=>"000001111",
99673=>"111110110",
99674=>"010000001",
99675=>"110011000",
99676=>"100100101",
99677=>"010010000",
99678=>"000011110",
99679=>"000000000",
99680=>"101101111",
99681=>"111111111",
99682=>"100110000",
99683=>"011000010",
99684=>"111111111",
99685=>"001001001",
99686=>"000000000",
99687=>"000101111",
99688=>"000000100",
99689=>"100000010",
99690=>"111011010",
99691=>"110000000",
99692=>"001111010",
99693=>"111011111",
99694=>"000000000",
99695=>"100000100",
99696=>"001000001",
99697=>"110111100",
99698=>"001000000",
99699=>"111111011",
99700=>"111111010",
99701=>"010000010",
99702=>"100000000",
99703=>"000111000",
99704=>"111000110",
99705=>"111110010",
99706=>"111000100",
99707=>"011000000",
99708=>"011001000",
99709=>"010011010",
99710=>"000011111",
99711=>"111100110",
99712=>"000100100",
99713=>"011011011",
99714=>"100000000",
99715=>"100000000",
99716=>"111000000",
99717=>"101010010",
99718=>"000100100",
99719=>"001000100",
99720=>"110110110",
99721=>"000100000",
99722=>"000000000",
99723=>"111111011",
99724=>"111111111",
99725=>"000000101",
99726=>"011000000",
99727=>"000111000",
99728=>"110011111",
99729=>"101000010",
99730=>"111000000",
99731=>"111111011",
99732=>"001100011",
99733=>"101110100",
99734=>"101101000",
99735=>"110110010",
99736=>"111101011",
99737=>"111000001",
99738=>"000011000",
99739=>"111111111",
99740=>"110100001",
99741=>"111100111",
99742=>"101100111",
99743=>"111111111",
99744=>"001100111",
99745=>"000000000",
99746=>"000000000",
99747=>"000100101",
99748=>"000000010",
99749=>"000000000",
99750=>"110110110",
99751=>"101000000",
99752=>"101001000",
99753=>"010010011",
99754=>"100000000",
99755=>"111011111",
99756=>"010001000",
99757=>"000000000",
99758=>"101000000",
99759=>"101001010",
99760=>"111011111",
99761=>"000010010",
99762=>"111001100",
99763=>"011001000",
99764=>"101001001",
99765=>"001000101",
99766=>"100010000",
99767=>"010010000",
99768=>"110100101",
99769=>"111101101",
99770=>"111011010",
99771=>"011001000",
99772=>"000000011",
99773=>"010011011",
99774=>"110100110",
99775=>"000000110",
99776=>"000000000",
99777=>"000000100",
99778=>"110000000",
99779=>"001011001",
99780=>"000000010",
99781=>"000011100",
99782=>"011111000",
99783=>"110011000",
99784=>"010110101",
99785=>"111111111",
99786=>"111000100",
99787=>"000000000",
99788=>"111101110",
99789=>"111110101",
99790=>"111100010",
99791=>"111111111",
99792=>"111010000",
99793=>"011011011",
99794=>"100110111",
99795=>"000101001",
99796=>"101000000",
99797=>"000010011",
99798=>"111111011",
99799=>"111111101",
99800=>"001101100",
99801=>"100000000",
99802=>"010001001",
99803=>"111111111",
99804=>"000001000",
99805=>"111110101",
99806=>"111111111",
99807=>"101111111",
99808=>"000000100",
99809=>"000010000",
99810=>"100000011",
99811=>"001001000",
99812=>"000010000",
99813=>"000000000",
99814=>"111111111",
99815=>"000010010",
99816=>"111111110",
99817=>"000000101",
99818=>"000001001",
99819=>"111010111",
99820=>"000000000",
99821=>"110000110",
99822=>"111111111",
99823=>"110000000",
99824=>"110000111",
99825=>"000011111",
99826=>"111111111",
99827=>"110011011",
99828=>"001011111",
99829=>"000000000",
99830=>"111011001",
99831=>"111001111",
99832=>"100000000",
99833=>"001000000",
99834=>"000100111",
99835=>"110000000",
99836=>"011111001",
99837=>"111000011",
99838=>"100100101",
99839=>"111111011",
99840=>"000101110",
99841=>"111111111",
99842=>"011000101",
99843=>"100101100",
99844=>"001001010",
99845=>"000001001",
99846=>"110011000",
99847=>"000000011",
99848=>"000000001",
99849=>"011000000",
99850=>"000000001",
99851=>"000010000",
99852=>"000000000",
99853=>"000010111",
99854=>"111010000",
99855=>"001001000",
99856=>"111001000",
99857=>"111010000",
99858=>"011101111",
99859=>"111111000",
99860=>"111111111",
99861=>"100110000",
99862=>"100111111",
99863=>"010110000",
99864=>"101001101",
99865=>"111010111",
99866=>"000000011",
99867=>"011110111",
99868=>"111111101",
99869=>"000100101",
99870=>"000111111",
99871=>"000000111",
99872=>"111000000",
99873=>"111011111",
99874=>"010011111",
99875=>"000000111",
99876=>"101101000",
99877=>"001001111",
99878=>"010110101",
99879=>"111101001",
99880=>"110000000",
99881=>"110000000",
99882=>"100101111",
99883=>"010111010",
99884=>"011101111",
99885=>"110110011",
99886=>"000101111",
99887=>"100000010",
99888=>"110000000",
99889=>"001001000",
99890=>"111010100",
99891=>"000100000",
99892=>"000000111",
99893=>"000001110",
99894=>"001000100",
99895=>"111000000",
99896=>"011000000",
99897=>"000001101",
99898=>"000101111",
99899=>"000010001",
99900=>"001001001",
99901=>"010111110",
99902=>"000001101",
99903=>"101111110",
99904=>"111001000",
99905=>"000000111",
99906=>"001101000",
99907=>"010100000",
99908=>"111000001",
99909=>"000000000",
99910=>"000000111",
99911=>"000000110",
99912=>"001001111",
99913=>"101101011",
99914=>"000001111",
99915=>"000000000",
99916=>"010000000",
99917=>"010011001",
99918=>"100110000",
99919=>"010010101",
99920=>"101110110",
99921=>"000010111",
99922=>"010011011",
99923=>"100100000",
99924=>"111111101",
99925=>"101111100",
99926=>"001110101",
99927=>"000010011",
99928=>"010111111",
99929=>"001101111",
99930=>"000111111",
99931=>"110000000",
99932=>"111000101",
99933=>"000001111",
99934=>"111010111",
99935=>"000000100",
99936=>"110010000",
99937=>"010000010",
99938=>"010000001",
99939=>"001101111",
99940=>"101101101",
99941=>"101000100",
99942=>"111001000",
99943=>"101110110",
99944=>"000000101",
99945=>"000001111",
99946=>"111000010",
99947=>"010000110",
99948=>"001111100",
99949=>"110010111",
99950=>"111001111",
99951=>"001001100",
99952=>"100000000",
99953=>"000000000",
99954=>"110000000",
99955=>"000011000",
99956=>"000000000",
99957=>"000000111",
99958=>"000001111",
99959=>"010011000",
99960=>"010101101",
99961=>"100100111",
99962=>"111000000",
99963=>"100100010",
99964=>"111011001",
99965=>"000001000",
99966=>"010000000",
99967=>"000000001",
99968=>"111000000",
99969=>"011111111",
99970=>"011010011",
99971=>"111101110",
99972=>"010111001",
99973=>"111100111",
99974=>"100100111",
99975=>"100001001",
99976=>"101101000",
99977=>"111010110",
99978=>"000110001",
99979=>"000001010",
99980=>"110110111",
99981=>"110000000",
99982=>"011000000",
99983=>"101000000",
99984=>"100001001",
99985=>"110011000",
99986=>"000000000",
99987=>"000001001",
99988=>"110110000",
99989=>"111000001",
99990=>"001111111",
99991=>"001000100",
99992=>"111010001",
99993=>"000111101",
99994=>"000010000",
99995=>"010000111",
99996=>"000011111",
99997=>"111010010",
99998=>"101000000",
99999=>"000001111",
100000=>"100100011",
100001=>"000000011",
100002=>"101001111",
100003=>"011011111",
100004=>"111111110",
100005=>"011010000",
100006=>"011011010",
100007=>"000001000",
100008=>"111110000",
100009=>"110110010",
100010=>"111101000",
100011=>"010001001",
100012=>"000111011",
100013=>"000001101",
100014=>"011011001",
100015=>"111000000",
100016=>"011111111",
100017=>"110100111",
100018=>"000101111",
100019=>"110110111",
100020=>"110011000",
100021=>"000000101",
100022=>"011000100",
100023=>"100001001",
100024=>"100100100",
100025=>"001000000",
100026=>"111111010",
100027=>"000001110",
100028=>"000110111",
100029=>"111000001",
100030=>"001011110",
100031=>"010000101",
100032=>"111111000",
100033=>"111000000",
100034=>"110111111",
100035=>"000001001",
100036=>"000000000",
100037=>"100100110",
100038=>"111111101",
100039=>"000010010",
100040=>"010000000",
100041=>"111101101",
100042=>"101101111",
100043=>"101000110",
100044=>"101000000",
100045=>"111100100",
100046=>"000000000",
100047=>"000000000",
100048=>"010111000",
100049=>"100101111",
100050=>"101000110",
100051=>"101001000",
100052=>"111001101",
100053=>"101101101",
100054=>"000010111",
100055=>"111011010",
100056=>"111111000",
100057=>"011111000",
100058=>"101101111",
100059=>"111000000",
100060=>"111110110",
100061=>"010010111",
100062=>"101010000",
100063=>"000000101",
100064=>"000000000",
100065=>"000000101",
100066=>"110111111",
100067=>"111001101",
100068=>"000000000",
100069=>"010110110",
100070=>"011000000",
100071=>"100101101",
100072=>"000000011",
100073=>"000011101",
100074=>"000000100",
100075=>"101111010",
100076=>"000000000",
100077=>"000000101",
100078=>"000000100",
100079=>"000000110",
100080=>"000000010",
100081=>"001001010",
100082=>"010001010",
100083=>"000001110",
100084=>"001101111",
100085=>"001111110",
100086=>"000000000",
100087=>"001001101",
100088=>"011000000",
100089=>"001000010",
100090=>"000110110",
100091=>"000000010",
100092=>"100001111",
100093=>"010110000",
100094=>"111001100",
100095=>"101101110",
100096=>"010010000",
100097=>"101101111",
100098=>"101001011",
100099=>"000111011",
100100=>"110111000",
100101=>"000100000",
100102=>"111110010",
100103=>"001010000",
100104=>"110110000",
100105=>"000000111",
100106=>"000000110",
100107=>"111101000",
100108=>"001101111",
100109=>"110110111",
100110=>"111001011",
100111=>"101111001",
100112=>"000010111",
100113=>"000111111",
100114=>"000001111",
100115=>"101011000",
100116=>"101101111",
100117=>"101001100",
100118=>"110111011",
100119=>"000000000",
100120=>"101000111",
100121=>"000000000",
100122=>"111010101",
100123=>"010100100",
100124=>"000010111",
100125=>"111001001",
100126=>"100010011",
100127=>"010011000",
100128=>"101000000",
100129=>"110101111",
100130=>"000001000",
100131=>"010100000",
100132=>"100000000",
100133=>"111011001",
100134=>"101100110",
100135=>"000000011",
100136=>"000001001",
100137=>"011101000",
100138=>"000000100",
100139=>"000101111",
100140=>"000000000",
100141=>"000000111",
100142=>"010001000",
100143=>"110111111",
100144=>"010111100",
100145=>"110100100",
100146=>"000000000",
100147=>"011110100",
100148=>"101001111",
100149=>"010110111",
100150=>"011001001",
100151=>"101111111",
100152=>"000011111",
100153=>"000111000",
100154=>"010010000",
100155=>"000010000",
100156=>"100001001",
100157=>"000111101",
100158=>"010000011",
100159=>"100110010",
100160=>"111001101",
100161=>"000010001",
100162=>"111110111",
100163=>"100111100",
100164=>"110010000",
100165=>"111100100",
100166=>"110111000",
100167=>"101100000",
100168=>"001110111",
100169=>"000010110",
100170=>"101000101",
100171=>"001010101",
100172=>"000000000",
100173=>"011011000",
100174=>"111111000",
100175=>"111110001",
100176=>"111001000",
100177=>"110000110",
100178=>"111011000",
100179=>"111011110",
100180=>"100000111",
100181=>"100110111",
100182=>"010100000",
100183=>"101101111",
100184=>"110000001",
100185=>"001111110",
100186=>"011111110",
100187=>"011111000",
100188=>"000010010",
100189=>"010011001",
100190=>"101000111",
100191=>"011111111",
100192=>"100000010",
100193=>"000000101",
100194=>"000001111",
100195=>"100111011",
100196=>"011011100",
100197=>"011101000",
100198=>"000000110",
100199=>"011111001",
100200=>"101111000",
100201=>"000010111",
100202=>"101110111",
100203=>"000001000",
100204=>"010000000",
100205=>"010000000",
100206=>"000010110",
100207=>"000100000",
100208=>"110000100",
100209=>"011001000",
100210=>"110100110",
100211=>"101011111",
100212=>"100001111",
100213=>"000000100",
100214=>"101100000",
100215=>"111000000",
100216=>"000110111",
100217=>"000010010",
100218=>"111111111",
100219=>"000000000",
100220=>"100010001",
100221=>"010110101",
100222=>"111111011",
100223=>"011000000",
100224=>"111000000",
100225=>"111100111",
100226=>"010000010",
100227=>"010110000",
100228=>"100000111",
100229=>"010000000",
100230=>"010010010",
100231=>"100110001",
100232=>"011011001",
100233=>"010001001",
100234=>"010000101",
100235=>"101001110",
100236=>"111000110",
100237=>"001011010",
100238=>"000000011",
100239=>"101000000",
100240=>"100011111",
100241=>"000111111",
100242=>"000010111",
100243=>"001000000",
100244=>"101000010",
100245=>"101101111",
100246=>"001010101",
100247=>"010100000",
100248=>"111111111",
100249=>"110110110",
100250=>"111010110",
100251=>"000000101",
100252=>"000000000",
100253=>"100101101",
100254=>"000000000",
100255=>"000001111",
100256=>"100010011",
100257=>"000111010",
100258=>"011000000",
100259=>"110111111",
100260=>"101000000",
100261=>"010110000",
100262=>"011100111",
100263=>"111000100",
100264=>"000101111",
100265=>"000000000",
100266=>"111101011",
100267=>"111101110",
100268=>"111101110",
100269=>"110101011",
100270=>"011011000",
100271=>"101011111",
100272=>"101000111",
100273=>"000110110",
100274=>"000010110",
100275=>"111110110",
100276=>"101110110",
100277=>"101010000",
100278=>"111100000",
100279=>"010000100",
100280=>"010010000",
100281=>"011010110",
100282=>"010010010",
100283=>"001001000",
100284=>"011000100",
100285=>"111000110",
100286=>"100011011",
100287=>"001000011",
100288=>"010011011",
100289=>"000000110",
100290=>"111010000",
100291=>"011101100",
100292=>"000000000",
100293=>"110000001",
100294=>"000111111",
100295=>"111000111",
100296=>"010011100",
100297=>"101101100",
100298=>"001101000",
100299=>"000010011",
100300=>"110010011",
100301=>"001110000",
100302=>"111100000",
100303=>"000110111",
100304=>"111000101",
100305=>"010110011",
100306=>"101001100",
100307=>"010011000",
100308=>"111001010",
100309=>"011011000",
100310=>"010000001",
100311=>"000000000",
100312=>"000000000",
100313=>"110111110",
100314=>"111010110",
100315=>"101101110",
100316=>"011111101",
100317=>"011011000",
100318=>"101001001",
100319=>"110101111",
100320=>"001101111",
100321=>"000101111",
100322=>"010001001",
100323=>"011100100",
100324=>"011001001",
100325=>"001101000",
100326=>"000000000",
100327=>"100110000",
100328=>"111111001",
100329=>"111000111",
100330=>"000011011",
100331=>"100100100",
100332=>"001000111",
100333=>"111111001",
100334=>"111100111",
100335=>"000000000",
100336=>"111000000",
100337=>"011000100",
100338=>"000010111",
100339=>"010011001",
100340=>"001001000",
100341=>"101101101",
100342=>"111000010",
100343=>"011111101",
100344=>"000011000",
100345=>"101000000",
100346=>"011011111",
100347=>"101000001",
100348=>"010010100",
100349=>"100101100",
100350=>"111111000",
100351=>"111111111",
100352=>"110110110",
100353=>"111111111",
100354=>"101000010",
100355=>"001101111",
100356=>"001000000",
100357=>"001101111",
100358=>"010000100",
100359=>"000000110",
100360=>"001001000",
100361=>"110000100",
100362=>"011111011",
100363=>"011100010",
100364=>"101101100",
100365=>"111000000",
100366=>"111001000",
100367=>"000000000",
100368=>"100000101",
100369=>"111111111",
100370=>"111001001",
100371=>"010111111",
100372=>"001000000",
100373=>"010000000",
100374=>"111111111",
100375=>"111011111",
100376=>"011110010",
100377=>"000000000",
100378=>"000000100",
100379=>"000000101",
100380=>"100001111",
100381=>"010111011",
100382=>"010111011",
100383=>"111111000",
100384=>"000001000",
100385=>"111111111",
100386=>"111001111",
100387=>"111011111",
100388=>"001001001",
100389=>"100010001",
100390=>"010111010",
100391=>"010100111",
100392=>"010111111",
100393=>"000000000",
100394=>"111111000",
100395=>"111111001",
100396=>"110111111",
100397=>"000010000",
100398=>"100101111",
100399=>"100100111",
100400=>"111100111",
100401=>"000000000",
100402=>"111111111",
100403=>"000111000",
100404=>"111111111",
100405=>"111101000",
100406=>"011111010",
100407=>"010111100",
100408=>"000000111",
100409=>"101101001",
100410=>"110100000",
100411=>"000000001",
100412=>"000000000",
100413=>"111111111",
100414=>"111100101",
100415=>"101101101",
100416=>"000000000",
100417=>"010010011",
100418=>"000000000",
100419=>"000111011",
100420=>"111101001",
100421=>"100000101",
100422=>"000000100",
100423=>"000111111",
100424=>"100000000",
100425=>"111111111",
100426=>"100100101",
100427=>"100000100",
100428=>"000000000",
100429=>"100100100",
100430=>"000000000",
100431=>"011010101",
100432=>"110111110",
100433=>"111111111",
100434=>"011100000",
100435=>"100101001",
100436=>"010111011",
100437=>"011111111",
100438=>"100100111",
100439=>"111111111",
100440=>"010010111",
100441=>"000000000",
100442=>"000001001",
100443=>"000000000",
100444=>"101000010",
100445=>"011011011",
100446=>"000001000",
100447=>"011111110",
100448=>"101000100",
100449=>"111111011",
100450=>"000000000",
100451=>"000110000",
100452=>"101001000",
100453=>"101101000",
100454=>"111101100",
100455=>"010000000",
100456=>"000101000",
100457=>"000101111",
100458=>"111101101",
100459=>"000000000",
100460=>"111000011",
100461=>"110111000",
100462=>"000000100",
100463=>"100001110",
100464=>"101000000",
100465=>"000000000",
100466=>"111111010",
100467=>"010010000",
100468=>"111101000",
100469=>"100000111",
100470=>"000111000",
100471=>"010000000",
100472=>"000000000",
100473=>"101001101",
100474=>"111101000",
100475=>"000000000",
100476=>"111111101",
100477=>"000001111",
100478=>"000010000",
100479=>"101000110",
100480=>"000000101",
100481=>"101100001",
100482=>"000100101",
100483=>"000001101",
100484=>"101001101",
100485=>"000000000",
100486=>"000000010",
100487=>"100001000",
100488=>"111100100",
100489=>"110000010",
100490=>"001010000",
100491=>"000000101",
100492=>"111011000",
100493=>"000100101",
100494=>"000000000",
100495=>"101000000",
100496=>"000101001",
100497=>"010010110",
100498=>"000000000",
100499=>"110010100",
100500=>"101011000",
100501=>"001000100",
100502=>"011111110",
100503=>"111100000",
100504=>"000110101",
100505=>"010011011",
100506=>"101000000",
100507=>"100101100",
100508=>"101101101",
100509=>"000000000",
100510=>"000000111",
100511=>"101101101",
100512=>"000001001",
100513=>"110111011",
100514=>"011010011",
100515=>"001000111",
100516=>"000110001",
100517=>"000100000",
100518=>"000000000",
100519=>"111111000",
100520=>"110010110",
100521=>"011111111",
100522=>"100000101",
100523=>"100000101",
100524=>"101111111",
100525=>"001000100",
100526=>"011011111",
100527=>"001010000",
100528=>"000000110",
100529=>"011111011",
100530=>"111101101",
100531=>"111000000",
100532=>"011011001",
100533=>"011000001",
100534=>"101000101",
100535=>"001001001",
100536=>"000000000",
100537=>"101011000",
100538=>"000000111",
100539=>"111111111",
100540=>"100110111",
100541=>"111001001",
100542=>"110100101",
100543=>"111011111",
100544=>"000111010",
100545=>"010000011",
100546=>"101111100",
100547=>"000000001",
100548=>"000000101",
100549=>"010110111",
100550=>"000000101",
100551=>"110011010",
100552=>"011111101",
100553=>"001111011",
100554=>"111111000",
100555=>"111000000",
100556=>"000000000",
100557=>"111111001",
100558=>"100000101",
100559=>"000101001",
100560=>"101111000",
100561=>"011111101",
100562=>"110000000",
100563=>"000000100",
100564=>"101100100",
100565=>"111111111",
100566=>"010010000",
100567=>"101001101",
100568=>"000010000",
100569=>"111101000",
100570=>"001001101",
100571=>"000100100",
100572=>"011111111",
100573=>"011011011",
100574=>"000000000",
100575=>"000001000",
100576=>"111100100",
100577=>"100100101",
100578=>"000010111",
100579=>"011011000",
100580=>"000000010",
100581=>"111111111",
100582=>"001000000",
100583=>"101011010",
100584=>"111101001",
100585=>"000111111",
100586=>"110111111",
100587=>"000000000",
100588=>"000000000",
100589=>"000000101",
100590=>"100000001",
100591=>"000000101",
100592=>"001001101",
100593=>"111011111",
100594=>"100000000",
100595=>"010111100",
100596=>"001011000",
100597=>"010111111",
100598=>"000100000",
100599=>"001101011",
100600=>"101100000",
100601=>"111111001",
100602=>"110011011",
100603=>"000111101",
100604=>"111000000",
100605=>"000101000",
100606=>"100000000",
100607=>"000000000",
100608=>"110111001",
100609=>"000000001",
100610=>"101110111",
100611=>"000000011",
100612=>"000000100",
100613=>"000110110",
100614=>"000111110",
100615=>"111101010",
100616=>"000100001",
100617=>"110110000",
100618=>"011111110",
100619=>"000110111",
100620=>"001001001",
100621=>"111111000",
100622=>"000111111",
100623=>"110000111",
100624=>"110000110",
100625=>"000010111",
100626=>"000001000",
100627=>"111000010",
100628=>"000000100",
100629=>"111001001",
100630=>"101001000",
100631=>"110000111",
100632=>"111000001",
100633=>"111111111",
100634=>"000001100",
100635=>"110110000",
100636=>"111111001",
100637=>"111000001",
100638=>"111110110",
100639=>"001001001",
100640=>"000110110",
100641=>"100000101",
100642=>"110100000",
100643=>"000111111",
100644=>"100101101",
100645=>"100110000",
100646=>"001000001",
100647=>"000100110",
100648=>"000100110",
100649=>"111000001",
100650=>"000001000",
100651=>"001100000",
100652=>"000011111",
100653=>"111011100",
100654=>"111111100",
100655=>"000000001",
100656=>"111111000",
100657=>"000011011",
100658=>"111000001",
100659=>"111111111",
100660=>"000110000",
100661=>"001001001",
100662=>"001001011",
100663=>"001001001",
100664=>"011001110",
100665=>"001101000",
100666=>"001001000",
100667=>"011001001",
100668=>"001001000",
100669=>"000001000",
100670=>"000110010",
100671=>"001111011",
100672=>"110000000",
100673=>"111110000",
100674=>"000100111",
100675=>"010011000",
100676=>"111001000",
100677=>"111110110",
100678=>"111111011",
100679=>"110010001",
100680=>"111001000",
100681=>"110111000",
100682=>"000110011",
100683=>"111010001",
100684=>"000111110",
100685=>"011011011",
100686=>"100011101",
100687=>"111111111",
100688=>"000000010",
100689=>"110010010",
100690=>"111110000",
100691=>"011111100",
100692=>"001000001",
100693=>"011000001",
100694=>"111111101",
100695=>"110110110",
100696=>"110000001",
100697=>"000001011",
100698=>"000001001",
100699=>"011001111",
100700=>"000000000",
100701=>"110110000",
100702=>"111001001",
100703=>"000110110",
100704=>"000000100",
100705=>"000111111",
100706=>"100110110",
100707=>"000000001",
100708=>"000100100",
100709=>"010001001",
100710=>"000110000",
100711=>"110110000",
100712=>"110110000",
100713=>"111000011",
100714=>"001000110",
100715=>"110100111",
100716=>"111011001",
100717=>"000111110",
100718=>"110111000",
100719=>"110110101",
100720=>"000111001",
100721=>"111011011",
100722=>"011000000",
100723=>"001000000",
100724=>"111111000",
100725=>"100000000",
100726=>"000101110",
100727=>"101000001",
100728=>"011011001",
100729=>"111000000",
100730=>"111101101",
100731=>"110011001",
100732=>"110100100",
100733=>"010110011",
100734=>"000000000",
100735=>"000110010",
100736=>"000100010",
100737=>"110000000",
100738=>"110001000",
100739=>"110110110",
100740=>"011100000",
100741=>"111110111",
100742=>"111011000",
100743=>"000000011",
100744=>"010111011",
100745=>"111111000",
100746=>"001110101",
100747=>"010000101",
100748=>"000001011",
100749=>"000000010",
100750=>"111001011",
100751=>"101000000",
100752=>"110001011",
100753=>"110100000",
100754=>"110110010",
100755=>"101000100",
100756=>"010110111",
100757=>"110100110",
100758=>"000100110",
100759=>"110100100",
100760=>"110110111",
100761=>"111111110",
100762=>"111010010",
100763=>"000000001",
100764=>"110011110",
100765=>"000111101",
100766=>"100100111",
100767=>"000110110",
100768=>"100101111",
100769=>"001001001",
100770=>"010001111",
100771=>"101000001",
100772=>"111111000",
100773=>"000011011",
100774=>"001010111",
100775=>"101001001",
100776=>"111001000",
100777=>"111001110",
100778=>"011001010",
100779=>"110110000",
100780=>"100000111",
100781=>"111101100",
100782=>"001010011",
100783=>"001011111",
100784=>"100001111",
100785=>"010011000",
100786=>"000110010",
100787=>"000000110",
100788=>"100110110",
100789=>"100000010",
100790=>"011100001",
100791=>"101011111",
100792=>"010110000",
100793=>"010100100",
100794=>"110111000",
100795=>"000110110",
100796=>"000110100",
100797=>"110011110",
100798=>"110110001",
100799=>"110001000",
100800=>"000111111",
100801=>"011011000",
100802=>"100000111",
100803=>"000111000",
100804=>"110010001",
100805=>"100101011",
100806=>"110111011",
100807=>"000010000",
100808=>"110000110",
100809=>"110001001",
100810=>"000001001",
100811=>"111111001",
100812=>"000010000",
100813=>"001011010",
100814=>"010110011",
100815=>"000001011",
100816=>"000110110",
100817=>"011111011",
100818=>"000101111",
100819=>"110111000",
100820=>"100001001",
100821=>"001011001",
100822=>"000010000",
100823=>"111010000",
100824=>"011001111",
100825=>"001001001",
100826=>"110110011",
100827=>"110110110",
100828=>"001001001",
100829=>"100000011",
100830=>"111001111",
100831=>"110110011",
100832=>"000000000",
100833=>"000000000",
100834=>"010001111",
100835=>"111100100",
100836=>"001000000",
100837=>"000001000",
100838=>"011110100",
100839=>"111011001",
100840=>"100000110",
100841=>"001111110",
100842=>"100111110",
100843=>"111111010",
100844=>"110001001",
100845=>"001001001",
100846=>"000000000",
100847=>"000000010",
100848=>"111001001",
100849=>"010001100",
100850=>"000000110",
100851=>"111111011",
100852=>"100100111",
100853=>"011011011",
100854=>"000001110",
100855=>"111101101",
100856=>"111000000",
100857=>"000000111",
100858=>"111101111",
100859=>"000010111",
100860=>"010010000",
100861=>"111001000",
100862=>"000111101",
100863=>"111001001",
100864=>"111011000",
100865=>"010001000",
100866=>"110000111",
100867=>"101001000",
100868=>"011100001",
100869=>"101101100",
100870=>"111101011",
100871=>"000000100",
100872=>"100000000",
100873=>"000000000",
100874=>"001000111",
100875=>"000000000",
100876=>"000001111",
100877=>"110101111",
100878=>"111101101",
100879=>"000010001",
100880=>"100100000",
100881=>"100000001",
100882=>"100110111",
100883=>"010000000",
100884=>"001110000",
100885=>"111101101",
100886=>"011111011",
100887=>"111000110",
100888=>"101100010",
100889=>"111111111",
100890=>"000001001",
100891=>"010111111",
100892=>"111111000",
100893=>"111001000",
100894=>"110000000",
100895=>"000111100",
100896=>"111111000",
100897=>"000000010",
100898=>"001101111",
100899=>"000101100",
100900=>"000000000",
100901=>"111110000",
100902=>"111011000",
100903=>"000011111",
100904=>"010010000",
100905=>"001101100",
100906=>"101000111",
100907=>"011101111",
100908=>"110011110",
100909=>"001010010",
100910=>"011011010",
100911=>"001101011",
100912=>"000010011",
100913=>"000000001",
100914=>"000101011",
100915=>"010000101",
100916=>"111000000",
100917=>"111111111",
100918=>"110000010",
100919=>"000111000",
100920=>"111100101",
100921=>"000000111",
100922=>"111000101",
100923=>"111010110",
100924=>"110110110",
100925=>"111111111",
100926=>"000100000",
100927=>"110111110",
100928=>"011000111",
100929=>"111111000",
100930=>"000000000",
100931=>"111101011",
100932=>"111000110",
100933=>"101101001",
100934=>"000011101",
100935=>"100000001",
100936=>"110001001",
100937=>"101111010",
100938=>"101101110",
100939=>"011101000",
100940=>"011111000",
100941=>"100000100",
100942=>"010000000",
100943=>"110010010",
100944=>"010001000",
100945=>"110111111",
100946=>"100000101",
100947=>"011101001",
100948=>"011111011",
100949=>"010111001",
100950=>"000100000",
100951=>"111001001",
100952=>"001001000",
100953=>"001000000",
100954=>"100100000",
100955=>"001100000",
100956=>"000000101",
100957=>"010001111",
100958=>"010010011",
100959=>"111110001",
100960=>"001000000",
100961=>"001111010",
100962=>"101001111",
100963=>"011100000",
100964=>"100000001",
100965=>"011111011",
100966=>"010010000",
100967=>"000111001",
100968=>"101111011",
100969=>"111000000",
100970=>"000100000",
100971=>"010010011",
100972=>"000000111",
100973=>"101000101",
100974=>"101101011",
100975=>"110110010",
100976=>"100000000",
100977=>"010011001",
100978=>"011000110",
100979=>"101101101",
100980=>"000000000",
100981=>"000000111",
100982=>"111001101",
100983=>"000101101",
100984=>"010111000",
100985=>"000111010",
100986=>"111110011",
100987=>"101000111",
100988=>"100110111",
100989=>"111100000",
100990=>"111111111",
100991=>"111101100",
100992=>"000000000",
100993=>"000100000",
100994=>"011010001",
100995=>"100011111",
100996=>"101001001",
100997=>"000111110",
100998=>"111111000",
100999=>"000011110",
101000=>"001001001",
101001=>"111111000",
101002=>"101000111",
101003=>"000100111",
101004=>"001011000",
101005=>"101111110",
101006=>"010010001",
101007=>"101001100",
101008=>"111111110",
101009=>"011101000",
101010=>"000110000",
101011=>"001011010",
101012=>"000111111",
101013=>"000000000",
101014=>"010010010",
101015=>"110000101",
101016=>"000000000",
101017=>"110111010",
101018=>"000010010",
101019=>"000000100",
101020=>"000100000",
101021=>"101001000",
101022=>"000000000",
101023=>"011000111",
101024=>"000100000",
101025=>"010111001",
101026=>"111100000",
101027=>"010000000",
101028=>"100100101",
101029=>"000100000",
101030=>"100001000",
101031=>"000011000",
101032=>"000000010",
101033=>"001000000",
101034=>"000101111",
101035=>"000000001",
101036=>"010110111",
101037=>"000000001",
101038=>"111000000",
101039=>"101001101",
101040=>"000101001",
101041=>"110000100",
101042=>"000000100",
101043=>"111001001",
101044=>"011111011",
101045=>"101111000",
101046=>"001001100",
101047=>"010010000",
101048=>"001011000",
101049=>"000110111",
101050=>"110111000",
101051=>"010010011",
101052=>"111011000",
101053=>"111011111",
101054=>"111110110",
101055=>"101111011",
101056=>"111011011",
101057=>"000001000",
101058=>"111111000",
101059=>"110001000",
101060=>"111111000",
101061=>"000000010",
101062=>"000000101",
101063=>"000101111",
101064=>"111000000",
101065=>"111111111",
101066=>"111101000",
101067=>"001100101",
101068=>"011011000",
101069=>"001011111",
101070=>"000001010",
101071=>"010110101",
101072=>"111010111",
101073=>"110000101",
101074=>"000010010",
101075=>"010010010",
101076=>"000110111",
101077=>"111011000",
101078=>"101000111",
101079=>"111010000",
101080=>"010000000",
101081=>"101000101",
101082=>"000001011",
101083=>"101000100",
101084=>"010111100",
101085=>"101000001",
101086=>"000101000",
101087=>"110010000",
101088=>"010111100",
101089=>"100100001",
101090=>"110100110",
101091=>"111001001",
101092=>"000010000",
101093=>"111011000",
101094=>"101100000",
101095=>"000000101",
101096=>"001001000",
101097=>"111111010",
101098=>"100000000",
101099=>"111000011",
101100=>"111000000",
101101=>"000000000",
101102=>"000001000",
101103=>"100001001",
101104=>"000001111",
101105=>"100001100",
101106=>"000000010",
101107=>"110100100",
101108=>"110101011",
101109=>"101001100",
101110=>"000000000",
101111=>"000101010",
101112=>"000111111",
101113=>"001101110",
101114=>"111100100",
101115=>"101111110",
101116=>"000001110",
101117=>"001111000",
101118=>"100000010",
101119=>"111000000",
101120=>"101000000",
101121=>"000000001",
101122=>"000000100",
101123=>"010000000",
101124=>"000000010",
101125=>"010000000",
101126=>"010010010",
101127=>"010011111",
101128=>"111000000",
101129=>"111101100",
101130=>"000001001",
101131=>"011001101",
101132=>"101000000",
101133=>"000111000",
101134=>"000011010",
101135=>"000100000",
101136=>"000100000",
101137=>"111111111",
101138=>"111010101",
101139=>"000111111",
101140=>"000001100",
101141=>"111111111",
101142=>"000000001",
101143=>"010111111",
101144=>"111111000",
101145=>"101000001",
101146=>"111000000",
101147=>"000000000",
101148=>"111000111",
101149=>"111111011",
101150=>"110111001",
101151=>"111111101",
101152=>"000000111",
101153=>"000101111",
101154=>"110111111",
101155=>"001100000",
101156=>"111101100",
101157=>"100111000",
101158=>"111000000",
101159=>"000001000",
101160=>"011111111",
101161=>"101100000",
101162=>"010000010",
101163=>"111110000",
101164=>"110110110",
101165=>"100101001",
101166=>"111111111",
101167=>"000101101",
101168=>"000000000",
101169=>"000100000",
101170=>"000101111",
101171=>"010111111",
101172=>"101000000",
101173=>"011100111",
101174=>"001011000",
101175=>"000000000",
101176=>"100000101",
101177=>"010111111",
101178=>"000110111",
101179=>"000000000",
101180=>"011111110",
101181=>"111000101",
101182=>"001100000",
101183=>"111001001",
101184=>"111111111",
101185=>"010000000",
101186=>"000100000",
101187=>"111101101",
101188=>"101011111",
101189=>"101111000",
101190=>"111111000",
101191=>"000000111",
101192=>"000000001",
101193=>"100000001",
101194=>"000000100",
101195=>"111100100",
101196=>"110111111",
101197=>"011001111",
101198=>"000000101",
101199=>"111100000",
101200=>"000000101",
101201=>"111111111",
101202=>"111011111",
101203=>"110100100",
101204=>"001000001",
101205=>"100111001",
101206=>"000100000",
101207=>"100111111",
101208=>"000001001",
101209=>"000111001",
101210=>"001011011",
101211=>"000011111",
101212=>"000000000",
101213=>"010011110",
101214=>"100000000",
101215=>"100001101",
101216=>"111000000",
101217=>"001101100",
101218=>"101000000",
101219=>"000010111",
101220=>"111101001",
101221=>"000001111",
101222=>"100001101",
101223=>"111110111",
101224=>"111111111",
101225=>"000000111",
101226=>"000110111",
101227=>"000000011",
101228=>"000111111",
101229=>"010010010",
101230=>"000000100",
101231=>"000000110",
101232=>"001001000",
101233=>"000000000",
101234=>"000111001",
101235=>"000111010",
101236=>"100111011",
101237=>"111000011",
101238=>"110111110",
101239=>"111111111",
101240=>"001001100",
101241=>"000000000",
101242=>"000000001",
101243=>"000101111",
101244=>"001001000",
101245=>"110011001",
101246=>"111001100",
101247=>"101000000",
101248=>"000000101",
101249=>"011010000",
101250=>"000110111",
101251=>"000110010",
101252=>"011111111",
101253=>"000111111",
101254=>"101110000",
101255=>"101101001",
101256=>"100010010",
101257=>"000100000",
101258=>"000000000",
101259=>"000000111",
101260=>"000000111",
101261=>"111101100",
101262=>"110011000",
101263=>"111000001",
101264=>"010100110",
101265=>"010001000",
101266=>"000000000",
101267=>"000000000",
101268=>"111011001",
101269=>"101101101",
101270=>"101111000",
101271=>"111111000",
101272=>"111000001",
101273=>"001111111",
101274=>"000111101",
101275=>"101000000",
101276=>"010111000",
101277=>"110111111",
101278=>"010111110",
101279=>"010010010",
101280=>"011101101",
101281=>"111111111",
101282=>"000000011",
101283=>"000000011",
101284=>"100111111",
101285=>"000111110",
101286=>"110100010",
101287=>"000100111",
101288=>"110100000",
101289=>"111001100",
101290=>"000000111",
101291=>"000000000",
101292=>"111110110",
101293=>"101000000",
101294=>"000000001",
101295=>"001000000",
101296=>"000000101",
101297=>"000110110",
101298=>"000011010",
101299=>"000000101",
101300=>"110000000",
101301=>"100110101",
101302=>"010000111",
101303=>"110111111",
101304=>"111111001",
101305=>"111110111",
101306=>"110010101",
101307=>"010101100",
101308=>"010000011",
101309=>"010010111",
101310=>"110111110",
101311=>"000000001",
101312=>"000000111",
101313=>"111000100",
101314=>"011111000",
101315=>"111001000",
101316=>"000000010",
101317=>"011101001",
101318=>"110111111",
101319=>"111111010",
101320=>"010010010",
101321=>"000000000",
101322=>"110111101",
101323=>"000000000",
101324=>"110111000",
101325=>"100000100",
101326=>"001011000",
101327=>"100011100",
101328=>"111010111",
101329=>"011001000",
101330=>"000000000",
101331=>"000100000",
101332=>"101000111",
101333=>"000011011",
101334=>"110111010",
101335=>"110110111",
101336=>"000000001",
101337=>"000000101",
101338=>"100011011",
101339=>"000110010",
101340=>"001110000",
101341=>"101100100",
101342=>"111010111",
101343=>"111101111",
101344=>"111000000",
101345=>"111101000",
101346=>"010011000",
101347=>"001011010",
101348=>"100000000",
101349=>"000000101",
101350=>"111000111",
101351=>"000000100",
101352=>"101100101",
101353=>"000000000",
101354=>"001000000",
101355=>"000111111",
101356=>"100100001",
101357=>"011000111",
101358=>"111101111",
101359=>"111000101",
101360=>"011000100",
101361=>"011110000",
101362=>"011000000",
101363=>"011011001",
101364=>"000101101",
101365=>"000000001",
101366=>"110000100",
101367=>"100110000",
101368=>"111111111",
101369=>"001111111",
101370=>"111100100",
101371=>"111001000",
101372=>"010010100",
101373=>"000000000",
101374=>"010110111",
101375=>"010111000",
101376=>"011111110",
101377=>"010000000",
101378=>"001000101",
101379=>"000000000",
101380=>"001111011",
101381=>"000000000",
101382=>"011111010",
101383=>"000000000",
101384=>"000000100",
101385=>"010000000",
101386=>"000011000",
101387=>"111001101",
101388=>"000000000",
101389=>"000000101",
101390=>"000001000",
101391=>"000000101",
101392=>"100100100",
101393=>"111010010",
101394=>"110110111",
101395=>"111000000",
101396=>"111111111",
101397=>"111111000",
101398=>"011101111",
101399=>"011000011",
101400=>"000000011",
101401=>"111101101",
101402=>"000000000",
101403=>"010011000",
101404=>"000100100",
101405=>"111000000",
101406=>"110111111",
101407=>"000000000",
101408=>"000011111",
101409=>"101001000",
101410=>"000011111",
101411=>"011111010",
101412=>"011000000",
101413=>"011100000",
101414=>"111001000",
101415=>"101111111",
101416=>"111100000",
101417=>"001111111",
101418=>"010110000",
101419=>"000010110",
101420=>"000011010",
101421=>"100000000",
101422=>"111000111",
101423=>"000000000",
101424=>"000000010",
101425=>"011111001",
101426=>"000000000",
101427=>"100000001",
101428=>"010011010",
101429=>"000000000",
101430=>"001011011",
101431=>"000001000",
101432=>"000000000",
101433=>"000000001",
101434=>"000000000",
101435=>"000000000",
101436=>"000000000",
101437=>"101100111",
101438=>"100000100",
101439=>"010011000",
101440=>"111111111",
101441=>"011011011",
101442=>"010111110",
101443=>"110110100",
101444=>"011011000",
101445=>"000000111",
101446=>"000011011",
101447=>"111111000",
101448=>"000000000",
101449=>"100110000",
101450=>"111111001",
101451=>"111001000",
101452=>"111110111",
101453=>"110111111",
101454=>"011111111",
101455=>"111101111",
101456=>"010001000",
101457=>"111011101",
101458=>"000000000",
101459=>"001100000",
101460=>"010011000",
101461=>"110111111",
101462=>"000000000",
101463=>"111100001",
101464=>"000010000",
101465=>"000010000",
101466=>"000100000",
101467=>"110000000",
101468=>"110000000",
101469=>"000000000",
101470=>"111111111",
101471=>"000011011",
101472=>"000010000",
101473=>"000000000",
101474=>"000010111",
101475=>"000001000",
101476=>"100101100",
101477=>"100000100",
101478=>"000000110",
101479=>"000000000",
101480=>"001111000",
101481=>"000100111",
101482=>"111001000",
101483=>"111111101",
101484=>"000000000",
101485=>"000100000",
101486=>"000000000",
101487=>"000000010",
101488=>"000011011",
101489=>"000000010",
101490=>"000110110",
101491=>"101110110",
101492=>"101111111",
101493=>"101000000",
101494=>"011111011",
101495=>"100101111",
101496=>"000000000",
101497=>"010111111",
101498=>"100000000",
101499=>"000100000",
101500=>"000100111",
101501=>"100100000",
101502=>"111111110",
101503=>"100000100",
101504=>"001111101",
101505=>"100000000",
101506=>"010001010",
101507=>"101111111",
101508=>"110000000",
101509=>"000000110",
101510=>"110000010",
101511=>"010100000",
101512=>"010111100",
101513=>"100000000",
101514=>"100000111",
101515=>"111111101",
101516=>"000000000",
101517=>"010000000",
101518=>"110111011",
101519=>"000000000",
101520=>"001001000",
101521=>"110111010",
101522=>"000001111",
101523=>"111101000",
101524=>"111001000",
101525=>"000000111",
101526=>"111001111",
101527=>"001011111",
101528=>"000001000",
101529=>"111111111",
101530=>"101100000",
101531=>"000000000",
101532=>"001010111",
101533=>"010000011",
101534=>"000011010",
101535=>"100000010",
101536=>"001111001",
101537=>"110011111",
101538=>"000101000",
101539=>"000111101",
101540=>"000111110",
101541=>"000000000",
101542=>"110111111",
101543=>"110111000",
101544=>"110110111",
101545=>"000000001",
101546=>"000000000",
101547=>"011011010",
101548=>"101100111",
101549=>"111111111",
101550=>"000011011",
101551=>"111101111",
101552=>"110100101",
101553=>"000001000",
101554=>"000000001",
101555=>"000000110",
101556=>"100100000",
101557=>"000011011",
101558=>"100010111",
101559=>"101001011",
101560=>"010000000",
101561=>"010100000",
101562=>"110001000",
101563=>"010010000",
101564=>"111101001",
101565=>"111111111",
101566=>"000110101",
101567=>"000000000",
101568=>"000000000",
101569=>"000010000",
101570=>"001000000",
101571=>"011011000",
101572=>"111001111",
101573=>"111000000",
101574=>"000001111",
101575=>"001000001",
101576=>"001000111",
101577=>"000111011",
101578=>"111111111",
101579=>"000000000",
101580=>"111000000",
101581=>"010011111",
101582=>"000011010",
101583=>"000011111",
101584=>"100101111",
101585=>"110111111",
101586=>"111000001",
101587=>"000000011",
101588=>"101111100",
101589=>"100111000",
101590=>"000000001",
101591=>"000000000",
101592=>"000000000",
101593=>"111000000",
101594=>"110111110",
101595=>"010100100",
101596=>"100111110",
101597=>"011000100",
101598=>"010000111",
101599=>"000000001",
101600=>"010111000",
101601=>"100000000",
101602=>"111111111",
101603=>"011101000",
101604=>"101001000",
101605=>"000111000",
101606=>"000011111",
101607=>"100110110",
101608=>"111100000",
101609=>"000010110",
101610=>"100110010",
101611=>"001111011",
101612=>"000000000",
101613=>"000011111",
101614=>"000010010",
101615=>"100000000",
101616=>"100000000",
101617=>"011111000",
101618=>"101100100",
101619=>"100001000",
101620=>"001111011",
101621=>"000001000",
101622=>"000000000",
101623=>"111101101",
101624=>"000111000",
101625=>"110000000",
101626=>"111111111",
101627=>"000000000",
101628=>"010010000",
101629=>"000001000",
101630=>"011010000",
101631=>"000001011",
101632=>"000000110",
101633=>"000110110",
101634=>"001011101",
101635=>"100111110",
101636=>"111110100",
101637=>"111011001",
101638=>"101000000",
101639=>"110000001",
101640=>"100101111",
101641=>"011011000",
101642=>"010011111",
101643=>"010011110",
101644=>"100100100",
101645=>"001011000",
101646=>"011000000",
101647=>"100000101",
101648=>"011000000",
101649=>"001011001",
101650=>"101101010",
101651=>"010010011",
101652=>"000100011",
101653=>"100110110",
101654=>"000100100",
101655=>"011011011",
101656=>"001010010",
101657=>"010000011",
101658=>"100110111",
101659=>"001011111",
101660=>"011011011",
101661=>"011011000",
101662=>"101001111",
101663=>"100000100",
101664=>"000011001",
101665=>"111110111",
101666=>"000000011",
101667=>"101011001",
101668=>"110110110",
101669=>"111100111",
101670=>"010011000",
101671=>"111111100",
101672=>"011100110",
101673=>"100000001",
101674=>"100100000",
101675=>"011000011",
101676=>"000100110",
101677=>"110110110",
101678=>"100000100",
101679=>"001100100",
101680=>"111000100",
101681=>"000010000",
101682=>"101100111",
101683=>"011000011",
101684=>"001011111",
101685=>"111110010",
101686=>"011001000",
101687=>"100000100",
101688=>"100110111",
101689=>"110000100",
101690=>"001001000",
101691=>"001001111",
101692=>"000000100",
101693=>"001001000",
101694=>"000000100",
101695=>"100111011",
101696=>"011010110",
101697=>"111010011",
101698=>"111011001",
101699=>"001011111",
101700=>"110100110",
101701=>"111011000",
101702=>"101110010",
101703=>"011101000",
101704=>"100100111",
101705=>"110101100",
101706=>"000010000",
101707=>"110100110",
101708=>"001011001",
101709=>"010100110",
101710=>"000100100",
101711=>"111100110",
101712=>"001011000",
101713=>"101101111",
101714=>"101100110",
101715=>"010010110",
101716=>"101000001",
101717=>"111100100",
101718=>"000000000",
101719=>"001011000",
101720=>"100100100",
101721=>"100100001",
101722=>"100101101",
101723=>"110110110",
101724=>"100101100",
101725=>"000010000",
101726=>"110100111",
101727=>"111001000",
101728=>"100110011",
101729=>"010100100",
101730=>"000001101",
101731=>"110110110",
101732=>"011101111",
101733=>"110100111",
101734=>"100110100",
101735=>"011001000",
101736=>"100000101",
101737=>"111101100",
101738=>"110011011",
101739=>"110010110",
101740=>"110110110",
101741=>"011011011",
101742=>"100100100",
101743=>"100100111",
101744=>"110100000",
101745=>"100110110",
101746=>"001011111",
101747=>"000000000",
101748=>"111111011",
101749=>"000001001",
101750=>"110110001",
101751=>"100011011",
101752=>"010011010",
101753=>"110000011",
101754=>"010100110",
101755=>"000100001",
101756=>"110110100",
101757=>"101001000",
101758=>"001001000",
101759=>"011011000",
101760=>"110010001",
101761=>"010010011",
101762=>"011011110",
101763=>"100101101",
101764=>"000000011",
101765=>"110010110",
101766=>"000000000",
101767=>"010000000",
101768=>"101000100",
101769=>"101100010",
101770=>"000000000",
101771=>"110011011",
101772=>"110010000",
101773=>"011001011",
101774=>"110100111",
101775=>"000100101",
101776=>"000100000",
101777=>"000000111",
101778=>"011011001",
101779=>"110010010",
101780=>"010100110",
101781=>"001001001",
101782=>"000100100",
101783=>"010010000",
101784=>"111111110",
101785=>"100000011",
101786=>"011011001",
101787=>"011011100",
101788=>"110100100",
101789=>"011111111",
101790=>"111011110",
101791=>"000001000",
101792=>"110100010",
101793=>"011000011",
101794=>"000100000",
101795=>"010110010",
101796=>"011111100",
101797=>"100000011",
101798=>"101111111",
101799=>"000000000",
101800=>"001011011",
101801=>"000100111",
101802=>"011011111",
101803=>"001011011",
101804=>"101100011",
101805=>"000000101",
101806=>"110110100",
101807=>"100100000",
101808=>"110110000",
101809=>"100110000",
101810=>"111011111",
101811=>"001111111",
101812=>"111111101",
101813=>"110011111",
101814=>"111100000",
101815=>"100100011",
101816=>"100101110",
101817=>"110110111",
101818=>"100110000",
101819=>"110011011",
101820=>"110111011",
101821=>"111011010",
101822=>"010011001",
101823=>"000000000",
101824=>"100100110",
101825=>"011011010",
101826=>"111011011",
101827=>"001100100",
101828=>"100100100",
101829=>"100000100",
101830=>"111010110",
101831=>"111000101",
101832=>"000111001",
101833=>"111110010",
101834=>"111010000",
101835=>"100110111",
101836=>"110011001",
101837=>"001001101",
101838=>"011011011",
101839=>"000011011",
101840=>"001001000",
101841=>"000000100",
101842=>"111100110",
101843=>"111110110",
101844=>"100110111",
101845=>"011101100",
101846=>"100100100",
101847=>"100011111",
101848=>"100100110",
101849=>"000100010",
101850=>"011111111",
101851=>"011011001",
101852=>"100000110",
101853=>"000110111",
101854=>"110110010",
101855=>"100000100",
101856=>"100100110",
101857=>"000000111",
101858=>"000001001",
101859=>"100110111",
101860=>"000000011",
101861=>"111100000",
101862=>"110000100",
101863=>"000000110",
101864=>"111011111",
101865=>"011011010",
101866=>"111111001",
101867=>"100101000",
101868=>"100100011",
101869=>"011111111",
101870=>"011011011",
101871=>"000010011",
101872=>"011010000",
101873=>"000100110",
101874=>"100111101",
101875=>"100100100",
101876=>"111110001",
101877=>"001011001",
101878=>"000000010",
101879=>"010000110",
101880=>"110010111",
101881=>"100000011",
101882=>"110100111",
101883=>"110110000",
101884=>"011110110",
101885=>"110110110",
101886=>"000000010",
101887=>"000100111",
101888=>"010011111",
101889=>"101001011",
101890=>"101101001",
101891=>"111110010",
101892=>"110111011",
101893=>"110000000",
101894=>"111000111",
101895=>"000000000",
101896=>"000111001",
101897=>"001001111",
101898=>"101101111",
101899=>"100101011",
101900=>"000111110",
101901=>"010110110",
101902=>"100000100",
101903=>"111000001",
101904=>"101101000",
101905=>"001001111",
101906=>"100100000",
101907=>"001011010",
101908=>"111101100",
101909=>"000000110",
101910=>"100111111",
101911=>"111000010",
101912=>"100000000",
101913=>"000001111",
101914=>"100001000",
101915=>"101001101",
101916=>"111000000",
101917=>"011101100",
101918=>"111110001",
101919=>"101111000",
101920=>"000000100",
101921=>"110011111",
101922=>"000011100",
101923=>"000010100",
101924=>"010111111",
101925=>"110000111",
101926=>"000000000",
101927=>"100001110",
101928=>"000010010",
101929=>"100111110",
101930=>"000000100",
101931=>"000010010",
101932=>"000011111",
101933=>"000000111",
101934=>"010011111",
101935=>"110010010",
101936=>"101101101",
101937=>"100111110",
101938=>"010010111",
101939=>"101000001",
101940=>"101101111",
101941=>"110110111",
101942=>"100000011",
101943=>"101001001",
101944=>"110000000",
101945=>"101000000",
101946=>"010101011",
101947=>"010001111",
101948=>"000000100",
101949=>"010111010",
101950=>"011001100",
101951=>"111011100",
101952=>"000110110",
101953=>"100010110",
101954=>"110111111",
101955=>"100000010",
101956=>"000110000",
101957=>"001000000",
101958=>"010101101",
101959=>"111101001",
101960=>"010001011",
101961=>"111101111",
101962=>"101000001",
101963=>"101101101",
101964=>"111000000",
101965=>"110110110",
101966=>"001011011",
101967=>"110111111",
101968=>"001000000",
101969=>"010010000",
101970=>"001000111",
101971=>"010000001",
101972=>"111101111",
101973=>"110111110",
101974=>"010011101",
101975=>"111001111",
101976=>"111000101",
101977=>"000001011",
101978=>"000100100",
101979=>"100010000",
101980=>"010000000",
101981=>"100001010",
101982=>"111001111",
101983=>"001000101",
101984=>"010010010",
101985=>"000000111",
101986=>"011000111",
101987=>"000000111",
101988=>"101001111",
101989=>"101100111",
101990=>"111110100",
101991=>"111010111",
101992=>"011000101",
101993=>"111000000",
101994=>"010111111",
101995=>"110111000",
101996=>"100111110",
101997=>"001000010",
101998=>"000101011",
101999=>"011000111",
102000=>"001000111",
102001=>"000000100",
102002=>"000000100",
102003=>"000010000",
102004=>"111010011",
102005=>"100101111",
102006=>"111000010",
102007=>"111000000",
102008=>"110111111",
102009=>"010011111",
102010=>"001001100",
102011=>"101001010",
102012=>"000100000",
102013=>"011101110",
102014=>"111110110",
102015=>"001101101",
102016=>"110110000",
102017=>"001111000",
102018=>"011000000",
102019=>"000010110",
102020=>"101001101",
102021=>"100111000",
102022=>"111001010",
102023=>"000000011",
102024=>"101100111",
102025=>"001000011",
102026=>"111001001",
102027=>"110010000",
102028=>"000000000",
102029=>"000000111",
102030=>"001001000",
102031=>"110000000",
102032=>"011111110",
102033=>"011111011",
102034=>"000000010",
102035=>"001100101",
102036=>"000101000",
102037=>"000000000",
102038=>"001001101",
102039=>"000010011",
102040=>"000111101",
102041=>"100010011",
102042=>"001101001",
102043=>"010001111",
102044=>"111100110",
102045=>"011101111",
102046=>"010010000",
102047=>"000100110",
102048=>"000111110",
102049=>"101000000",
102050=>"000110100",
102051=>"010101100",
102052=>"110010111",
102053=>"000110100",
102054=>"000110000",
102055=>"010111000",
102056=>"001000111",
102057=>"000001111",
102058=>"111101000",
102059=>"111000000",
102060=>"000000100",
102061=>"111000000",
102062=>"111100100",
102063=>"000100010",
102064=>"110010011",
102065=>"001000110",
102066=>"101101101",
102067=>"000000000",
102068=>"100011001",
102069=>"111011101",
102070=>"000011011",
102071=>"110110101",
102072=>"011010101",
102073=>"000101101",
102074=>"010000101",
102075=>"111111000",
102076=>"110000000",
102077=>"000100111",
102078=>"001001000",
102079=>"000000000",
102080=>"101000000",
102081=>"111001101",
102082=>"001000110",
102083=>"011010110",
102084=>"000110000",
102085=>"001010011",
102086=>"010100000",
102087=>"000010111",
102088=>"000010100",
102089=>"000110010",
102090=>"110111111",
102091=>"000000111",
102092=>"111100100",
102093=>"001001000",
102094=>"011000001",
102095=>"000010111",
102096=>"000000010",
102097=>"000110110",
102098=>"001101111",
102099=>"000111111",
102100=>"111100000",
102101=>"100001101",
102102=>"111001010",
102103=>"000011000",
102104=>"000000000",
102105=>"000110010",
102106=>"000110110",
102107=>"111000000",
102108=>"001111111",
102109=>"100000011",
102110=>"010000101",
102111=>"001000000",
102112=>"100111111",
102113=>"101000001",
102114=>"111101001",
102115=>"001100000",
102116=>"100101001",
102117=>"100001011",
102118=>"000010011",
102119=>"001001010",
102120=>"010010111",
102121=>"100001101",
102122=>"101111110",
102123=>"100110000",
102124=>"000110110",
102125=>"000110110",
102126=>"000000000",
102127=>"000101000",
102128=>"001011111",
102129=>"100011111",
102130=>"000001101",
102131=>"010100101",
102132=>"110110100",
102133=>"111100111",
102134=>"000000111",
102135=>"001001111",
102136=>"000000000",
102137=>"101110110",
102138=>"100100000",
102139=>"101111111",
102140=>"111110001",
102141=>"000101011",
102142=>"111111101",
102143=>"000000000",
102144=>"110111000",
102145=>"100000110",
102146=>"001000101",
102147=>"111101101",
102148=>"111011001",
102149=>"000001111",
102150=>"010111110",
102151=>"110000010",
102152=>"111000101",
102153=>"010110000",
102154=>"111111011",
102155=>"111111111",
102156=>"101001001",
102157=>"111011111",
102158=>"011111111",
102159=>"000001110",
102160=>"111111001",
102161=>"000111010",
102162=>"100101101",
102163=>"000000011",
102164=>"000011011",
102165=>"011111000",
102166=>"000000000",
102167=>"111101000",
102168=>"010111001",
102169=>"101001111",
102170=>"011010111",
102171=>"010111110",
102172=>"000011101",
102173=>"010000010",
102174=>"111101101",
102175=>"001000000",
102176=>"001000001",
102177=>"001000100",
102178=>"111000010",
102179=>"000100101",
102180=>"001001101",
102181=>"100011111",
102182=>"110110110",
102183=>"001111111",
102184=>"011110011",
102185=>"010000011",
102186=>"111111011",
102187=>"010001100",
102188=>"011001000",
102189=>"001000001",
102190=>"000000000",
102191=>"111001111",
102192=>"000000010",
102193=>"111011001",
102194=>"000001000",
102195=>"001001001",
102196=>"111110111",
102197=>"111110011",
102198=>"010000000",
102199=>"010000110",
102200=>"111001111",
102201=>"000000000",
102202=>"001001000",
102203=>"000000001",
102204=>"110110110",
102205=>"111111111",
102206=>"000010010",
102207=>"111111011",
102208=>"011010000",
102209=>"111111000",
102210=>"101101111",
102211=>"111110111",
102212=>"001000111",
102213=>"010101000",
102214=>"000010001",
102215=>"111000100",
102216=>"001001011",
102217=>"110110000",
102218=>"000001111",
102219=>"101001001",
102220=>"000000000",
102221=>"100101110",
102222=>"011001110",
102223=>"001101001",
102224=>"110110110",
102225=>"000010100",
102226=>"110111111",
102227=>"111001001",
102228=>"000010010",
102229=>"100101100",
102230=>"111101110",
102231=>"110111001",
102232=>"100101110",
102233=>"110100101",
102234=>"110100000",
102235=>"101101111",
102236=>"000000110",
102237=>"001000000",
102238=>"001001000",
102239=>"011111111",
102240=>"000011111",
102241=>"110110110",
102242=>"010000000",
102243=>"100000000",
102244=>"111101100",
102245=>"001011001",
102246=>"010110111",
102247=>"010000001",
102248=>"010111111",
102249=>"010111111",
102250=>"001000000",
102251=>"101110111",
102252=>"010011111",
102253=>"110111010",
102254=>"111000000",
102255=>"000000101",
102256=>"010110100",
102257=>"111111110",
102258=>"000110000",
102259=>"101111111",
102260=>"111111010",
102261=>"000100011",
102262=>"111110110",
102263=>"110110110",
102264=>"101000000",
102265=>"111101000",
102266=>"000000011",
102267=>"111101001",
102268=>"010100110",
102269=>"011001000",
102270=>"111110111",
102271=>"110110110",
102272=>"001111110",
102273=>"111010000",
102274=>"111110111",
102275=>"111011100",
102276=>"110111111",
102277=>"000000001",
102278=>"001111111",
102279=>"100111101",
102280=>"011001011",
102281=>"110110110",
102282=>"010111010",
102283=>"001000000",
102284=>"001000000",
102285=>"110000000",
102286=>"111111111",
102287=>"001000001",
102288=>"001100100",
102289=>"000101000",
102290=>"101101111",
102291=>"100000000",
102292=>"101111111",
102293=>"110110101",
102294=>"111001000",
102295=>"110001001",
102296=>"010110010",
102297=>"101100111",
102298=>"001000000",
102299=>"000000100",
102300=>"000000000",
102301=>"101100101",
102302=>"111001111",
102303=>"110110000",
102304=>"100000000",
102305=>"000010000",
102306=>"010000011",
102307=>"111100000",
102308=>"011011101",
102309=>"000011110",
102310=>"011111010",
102311=>"000010110",
102312=>"000101111",
102313=>"110101111",
102314=>"101000000",
102315=>"110000000",
102316=>"001000101",
102317=>"111010000",
102318=>"001001011",
102319=>"000000000",
102320=>"000000000",
102321=>"001011011",
102322=>"000010000",
102323=>"111101000",
102324=>"010111001",
102325=>"100000000",
102326=>"100100100",
102327=>"101111111",
102328=>"111110011",
102329=>"101111111",
102330=>"111111110",
102331=>"111000011",
102332=>"000110111",
102333=>"011111111",
102334=>"101001111",
102335=>"000000000",
102336=>"001000000",
102337=>"111000000",
102338=>"111111010",
102339=>"111101100",
102340=>"010111110",
102341=>"001001011",
102342=>"000000111",
102343=>"100000000",
102344=>"101100000",
102345=>"101110110",
102346=>"100000111",
102347=>"101000000",
102348=>"110010010",
102349=>"110010110",
102350=>"000010000",
102351=>"000111111",
102352=>"001010000",
102353=>"010111110",
102354=>"110100111",
102355=>"100100110",
102356=>"101000001",
102357=>"000000000",
102358=>"110110000",
102359=>"110100000",
102360=>"000000000",
102361=>"000110111",
102362=>"011001010",
102363=>"101111001",
102364=>"000000010",
102365=>"001011001",
102366=>"001000001",
102367=>"111100000",
102368=>"010010010",
102369=>"010111111",
102370=>"111110000",
102371=>"101111111",
102372=>"011000000",
102373=>"000000000",
102374=>"110000111",
102375=>"010000000",
102376=>"111110111",
102377=>"000000111",
102378=>"110110110",
102379=>"110110010",
102380=>"110111110",
102381=>"111101001",
102382=>"001001000",
102383=>"110110110",
102384=>"000110110",
102385=>"111001001",
102386=>"111111101",
102387=>"111111010",
102388=>"010100100",
102389=>"000001000",
102390=>"110111111",
102391=>"110111100",
102392=>"000000000",
102393=>"111111010",
102394=>"000111110",
102395=>"000111111",
102396=>"000111111",
102397=>"010010100",
102398=>"001100110",
102399=>"000000000",
102400=>"010110110",
102401=>"010011111",
102402=>"000000000",
102403=>"000000010",
102404=>"010110111",
102405=>"000000011",
102406=>"111111111",
102407=>"111111010",
102408=>"000000000",
102409=>"001001101",
102410=>"000000001",
102411=>"001100100",
102412=>"000000000",
102413=>"000000001",
102414=>"010110100",
102415=>"111111111",
102416=>"000000000",
102417=>"001111101",
102418=>"111111110",
102419=>"111100111",
102420=>"100000011",
102421=>"001001111",
102422=>"111100100",
102423=>"010111000",
102424=>"111001111",
102425=>"111110000",
102426=>"011000000",
102427=>"111101000",
102428=>"111111001",
102429=>"000111101",
102430=>"101100011",
102431=>"001111100",
102432=>"000000000",
102433=>"011000000",
102434=>"111001101",
102435=>"000000000",
102436=>"010111011",
102437=>"111111101",
102438=>"110111010",
102439=>"111000000",
102440=>"000010000",
102441=>"100111000",
102442=>"110111000",
102443=>"100000000",
102444=>"011111011",
102445=>"010101101",
102446=>"000111110",
102447=>"110000000",
102448=>"111111101",
102449=>"101100001",
102450=>"101000000",
102451=>"001011110",
102452=>"001100111",
102453=>"011111111",
102454=>"111010000",
102455=>"100000110",
102456=>"000000111",
102457=>"111111111",
102458=>"111101000",
102459=>"111011001",
102460=>"111110001",
102461=>"111111111",
102462=>"111101101",
102463=>"000001000",
102464=>"101101100",
102465=>"100111110",
102466=>"001101010",
102467=>"000000111",
102468=>"111110101",
102469=>"101101101",
102470=>"111000100",
102471=>"000011111",
102472=>"000010000",
102473=>"111000010",
102474=>"111111111",
102475=>"110100000",
102476=>"000000000",
102477=>"111111111",
102478=>"111001011",
102479=>"110001101",
102480=>"000110111",
102481=>"111111111",
102482=>"111010111",
102483=>"011111110",
102484=>"111111111",
102485=>"001001000",
102486=>"101111110",
102487=>"101101101",
102488=>"001000000",
102489=>"111111110",
102490=>"100001001",
102491=>"000110100",
102492=>"111111000",
102493=>"101101100",
102494=>"111101111",
102495=>"001000111",
102496=>"000000000",
102497=>"000000000",
102498=>"111001111",
102499=>"111111110",
102500=>"111111111",
102501=>"000100100",
102502=>"110111111",
102503=>"100111101",
102504=>"101101111",
102505=>"010000000",
102506=>"001111000",
102507=>"110110111",
102508=>"000000000",
102509=>"000100000",
102510=>"000111111",
102511=>"101011000",
102512=>"010111111",
102513=>"111111010",
102514=>"111101100",
102515=>"001000000",
102516=>"111110111",
102517=>"100100100",
102518=>"000000110",
102519=>"010000101",
102520=>"000010010",
102521=>"111111000",
102522=>"011111111",
102523=>"000000000",
102524=>"111011111",
102525=>"101101011",
102526=>"001000111",
102527=>"101001111",
102528=>"110111111",
102529=>"000000000",
102530=>"010010100",
102531=>"001000111",
102532=>"111111111",
102533=>"000111111",
102534=>"100110111",
102535=>"000010000",
102536=>"100110111",
102537=>"001011011",
102538=>"100101100",
102539=>"000101110",
102540=>"000000101",
102541=>"101100110",
102542=>"100000001",
102543=>"001000000",
102544=>"110011001",
102545=>"000100101",
102546=>"111111001",
102547=>"000000111",
102548=>"111111101",
102549=>"000101111",
102550=>"110111010",
102551=>"111110110",
102552=>"111110000",
102553=>"000010101",
102554=>"000010000",
102555=>"000000001",
102556=>"110100100",
102557=>"000100000",
102558=>"010111010",
102559=>"001111111",
102560=>"000000000",
102561=>"111011111",
102562=>"000000001",
102563=>"110000000",
102564=>"011111110",
102565=>"011111101",
102566=>"101001001",
102567=>"000010000",
102568=>"000111111",
102569=>"001000000",
102570=>"011001111",
102571=>"011101011",
102572=>"000000101",
102573=>"101101111",
102574=>"111011011",
102575=>"000000100",
102576=>"000000111",
102577=>"000000000",
102578=>"000101000",
102579=>"001000000",
102580=>"111000001",
102581=>"011101111",
102582=>"000110100",
102583=>"111110111",
102584=>"010110100",
102585=>"101101101",
102586=>"110110100",
102587=>"111101101",
102588=>"111110110",
102589=>"000000000",
102590=>"000000000",
102591=>"000001111",
102592=>"000000110",
102593=>"111111101",
102594=>"010011000",
102595=>"001001001",
102596=>"111111000",
102597=>"111111111",
102598=>"010111000",
102599=>"110111110",
102600=>"111111001",
102601=>"100100000",
102602=>"111010111",
102603=>"000001001",
102604=>"110110111",
102605=>"111111111",
102606=>"111101111",
102607=>"001000001",
102608=>"000111111",
102609=>"001001001",
102610=>"111100111",
102611=>"111111011",
102612=>"010111111",
102613=>"011001101",
102614=>"000000000",
102615=>"110111011",
102616=>"110110010",
102617=>"010011010",
102618=>"000000001",
102619=>"000000000",
102620=>"111101001",
102621=>"000000000",
102622=>"111011000",
102623=>"111011111",
102624=>"000001111",
102625=>"000001111",
102626=>"001000100",
102627=>"000000000",
102628=>"000100000",
102629=>"010100011",
102630=>"101000000",
102631=>"011011110",
102632=>"000000000",
102633=>"001001110",
102634=>"000000100",
102635=>"101001111",
102636=>"000000000",
102637=>"011110001",
102638=>"000111110",
102639=>"110101111",
102640=>"001100101",
102641=>"000010111",
102642=>"111111000",
102643=>"111111001",
102644=>"111111001",
102645=>"000000001",
102646=>"010011111",
102647=>"101000111",
102648=>"110111000",
102649=>"001101100",
102650=>"011111111",
102651=>"001111111",
102652=>"111111010",
102653=>"001000000",
102654=>"000111000",
102655=>"111111110",
102656=>"010000101",
102657=>"010000000",
102658=>"101100100",
102659=>"100000000",
102660=>"011001011",
102661=>"001001110",
102662=>"111000111",
102663=>"000111111",
102664=>"000011011",
102665=>"000010011",
102666=>"000000001",
102667=>"100000000",
102668=>"000000100",
102669=>"010000000",
102670=>"000111111",
102671=>"100100111",
102672=>"100011000",
102673=>"000000000",
102674=>"000100011",
102675=>"100100000",
102676=>"001011010",
102677=>"100000100",
102678=>"111111101",
102679=>"011000011",
102680=>"000000000",
102681=>"111100011",
102682=>"000100111",
102683=>"111011010",
102684=>"100100000",
102685=>"000000111",
102686=>"000011000",
102687=>"000010011",
102688=>"000101111",
102689=>"111011011",
102690=>"010110100",
102691=>"000000000",
102692=>"011011001",
102693=>"001110110",
102694=>"100100100",
102695=>"011100111",
102696=>"100100111",
102697=>"010111111",
102698=>"111011010",
102699=>"110100010",
102700=>"001011000",
102701=>"000001000",
102702=>"000000100",
102703=>"010110011",
102704=>"000111111",
102705=>"000100011",
102706=>"000101111",
102707=>"000101100",
102708=>"001000110",
102709=>"100000100",
102710=>"111110110",
102711=>"011011000",
102712=>"000000000",
102713=>"000000000",
102714=>"111100110",
102715=>"100101000",
102716=>"010001110",
102717=>"111111111",
102718=>"000000100",
102719=>"011011011",
102720=>"100100111",
102721=>"101111001",
102722=>"111011011",
102723=>"011111011",
102724=>"000010000",
102725=>"100100100",
102726=>"011111011",
102727=>"111011011",
102728=>"100011110",
102729=>"011011000",
102730=>"000000000",
102731=>"111001100",
102732=>"000111111",
102733=>"100111111",
102734=>"000110110",
102735=>"000010100",
102736=>"100110000",
102737=>"111011001",
102738=>"011110101",
102739=>"000100001",
102740=>"100100110",
102741=>"100000111",
102742=>"110100110",
102743=>"000000011",
102744=>"000000111",
102745=>"100110000",
102746=>"100110110",
102747=>"010010000",
102748=>"111011000",
102749=>"100001001",
102750=>"011111011",
102751=>"111011110",
102752=>"111000010",
102753=>"101000010",
102754=>"100000000",
102755=>"011000000",
102756=>"000001000",
102757=>"000100111",
102758=>"101000101",
102759=>"111111101",
102760=>"010011111",
102761=>"011000010",
102762=>"011000100",
102763=>"111101111",
102764=>"100100111",
102765=>"111100000",
102766=>"010100110",
102767=>"001000010",
102768=>"000000000",
102769=>"110000000",
102770=>"011011000",
102771=>"011101100",
102772=>"111010000",
102773=>"111100000",
102774=>"011011011",
102775=>"111111011",
102776=>"010000011",
102777=>"011011000",
102778=>"000100101",
102779=>"100101010",
102780=>"000010011",
102781=>"001000010",
102782=>"100111111",
102783=>"000000000",
102784=>"000011010",
102785=>"111110011",
102786=>"111111010",
102787=>"000111000",
102788=>"001111000",
102789=>"000100100",
102790=>"010001001",
102791=>"001001000",
102792=>"000111101",
102793=>"101100001",
102794=>"000100100",
102795=>"111000111",
102796=>"010010000",
102797=>"000000101",
102798=>"111111011",
102799=>"010101100",
102800=>"000110110",
102801=>"000000100",
102802=>"100100111",
102803=>"011000000",
102804=>"001001000",
102805=>"111111100",
102806=>"000000010",
102807=>"000000011",
102808=>"000011111",
102809=>"000101111",
102810=>"110100100",
102811=>"111110111",
102812=>"111111111",
102813=>"000011111",
102814=>"000100010",
102815=>"110100100",
102816=>"000100001",
102817=>"100110000",
102818=>"111011111",
102819=>"000000011",
102820=>"111100001",
102821=>"000000000",
102822=>"100111111",
102823=>"100000000",
102824=>"111100000",
102825=>"000011011",
102826=>"111100100",
102827=>"000000000",
102828=>"111001100",
102829=>"001011111",
102830=>"011110000",
102831=>"000011111",
102832=>"100000111",
102833=>"001110000",
102834=>"111101010",
102835=>"000000011",
102836=>"000111000",
102837=>"011011100",
102838=>"000111111",
102839=>"000100011",
102840=>"000001011",
102841=>"001011001",
102842=>"011111000",
102843=>"010011010",
102844=>"000000000",
102845=>"000111011",
102846=>"111111000",
102847=>"111111000",
102848=>"000000100",
102849=>"010000000",
102850=>"000011111",
102851=>"100100110",
102852=>"011000010",
102853=>"111111000",
102854=>"000011011",
102855=>"111101000",
102856=>"111111000",
102857=>"100110000",
102858=>"000011000",
102859=>"011011011",
102860=>"111111000",
102861=>"100010011",
102862=>"000000110",
102863=>"111111100",
102864=>"000000000",
102865=>"000000000",
102866=>"110100000",
102867=>"111111000",
102868=>"000000000",
102869=>"100111111",
102870=>"111000010",
102871=>"010000000",
102872=>"100100111",
102873=>"000011011",
102874=>"110100000",
102875=>"100100100",
102876=>"111111101",
102877=>"000011001",
102878=>"100111111",
102879=>"010000000",
102880=>"111011011",
102881=>"101100100",
102882=>"111000000",
102883=>"100001000",
102884=>"010101111",
102885=>"011011011",
102886=>"000010100",
102887=>"001111011",
102888=>"000100000",
102889=>"011000001",
102890=>"100000000",
102891=>"000000001",
102892=>"001000000",
102893=>"110100000",
102894=>"111100101",
102895=>"011000000",
102896=>"000100100",
102897=>"001001110",
102898=>"111011100",
102899=>"000000010",
102900=>"111101000",
102901=>"000000000",
102902=>"000000111",
102903=>"111100111",
102904=>"101000110",
102905=>"000111111",
102906=>"011000000",
102907=>"101111010",
102908=>"100000000",
102909=>"000011011",
102910=>"000110110",
102911=>"001011010",
102912=>"000000100",
102913=>"101101111",
102914=>"101000101",
102915=>"000000000",
102916=>"101000000",
102917=>"100000001",
102918=>"111000110",
102919=>"111111111",
102920=>"111101000",
102921=>"101101100",
102922=>"010100111",
102923=>"100000001",
102924=>"101000110",
102925=>"000001000",
102926=>"011000110",
102927=>"000011111",
102928=>"011000000",
102929=>"000101000",
102930=>"111101011",
102931=>"101100000",
102932=>"111111111",
102933=>"000010000",
102934=>"100000010",
102935=>"101111101",
102936=>"000101001",
102937=>"111101101",
102938=>"111001000",
102939=>"000100111",
102940=>"100101000",
102941=>"010011111",
102942=>"000101000",
102943=>"000010000",
102944=>"110111101",
102945=>"000000111",
102946=>"010110111",
102947=>"111000000",
102948=>"100110110",
102949=>"100001111",
102950=>"000010000",
102951=>"111010100",
102952=>"000010000",
102953=>"011111011",
102954=>"101100010",
102955=>"110010000",
102956=>"001111000",
102957=>"111100000",
102958=>"100101111",
102959=>"111001000",
102960=>"000101000",
102961=>"000000000",
102962=>"110110010",
102963=>"000101000",
102964=>"101010111",
102965=>"000010010",
102966=>"101110110",
102967=>"000000010",
102968=>"010111001",
102969=>"000001011",
102970=>"110010010",
102971=>"101110100",
102972=>"110001001",
102973=>"101010100",
102974=>"100000100",
102975=>"011111011",
102976=>"111101111",
102977=>"000111001",
102978=>"011101101",
102979=>"100000101",
102980=>"111101111",
102981=>"000101000",
102982=>"000111111",
102983=>"111111011",
102984=>"010110000",
102985=>"111101111",
102986=>"100100110",
102987=>"000010000",
102988=>"010000001",
102989=>"000000011",
102990=>"100000100",
102991=>"010110100",
102992=>"001101111",
102993=>"111111110",
102994=>"011101101",
102995=>"110011000",
102996=>"101100101",
102997=>"111110111",
102998=>"001011001",
102999=>"101000111",
103000=>"111000101",
103001=>"100001000",
103002=>"011001000",
103003=>"001001100",
103004=>"000000101",
103005=>"011001000",
103006=>"111010000",
103007=>"001000100",
103008=>"111001000",
103009=>"000000000",
103010=>"101000001",
103011=>"110100000",
103012=>"110000011",
103013=>"110100100",
103014=>"010101111",
103015=>"010111000",
103016=>"101111000",
103017=>"100101000",
103018=>"110000010",
103019=>"010100111",
103020=>"010111111",
103021=>"010011001",
103022=>"100100101",
103023=>"000111111",
103024=>"001000111",
103025=>"100100100",
103026=>"101111001",
103027=>"011000100",
103028=>"110010010",
103029=>"111101000",
103030=>"101101010",
103031=>"010000000",
103032=>"110000000",
103033=>"000110010",
103034=>"000111101",
103035=>"000011000",
103036=>"011001010",
103037=>"011110000",
103038=>"010110000",
103039=>"101001111",
103040=>"000000000",
103041=>"001000111",
103042=>"000000101",
103043=>"010010110",
103044=>"101000000",
103045=>"110111000",
103046=>"000100110",
103047=>"000000100",
103048=>"101001111",
103049=>"000101001",
103050=>"011011011",
103051=>"101001000",
103052=>"000000101",
103053=>"101001101",
103054=>"000000000",
103055=>"101000000",
103056=>"001011010",
103057=>"100000100",
103058=>"101000100",
103059=>"000001110",
103060=>"011101000",
103061=>"100100000",
103062=>"111101111",
103063=>"100111011",
103064=>"010010001",
103065=>"101000000",
103066=>"010111111",
103067=>"111111000",
103068=>"111100101",
103069=>"000000101",
103070=>"100111000",
103071=>"101101111",
103072=>"110111110",
103073=>"101111011",
103074=>"110011000",
103075=>"100010111",
103076=>"010110000",
103077=>"000100101",
103078=>"001110000",
103079=>"000101000",
103080=>"000100100",
103081=>"101101111",
103082=>"111101100",
103083=>"101000101",
103084=>"000111111",
103085=>"110000011",
103086=>"011011111",
103087=>"111010100",
103088=>"000000000",
103089=>"000001010",
103090=>"111100110",
103091=>"000000010",
103092=>"010011001",
103093=>"011111110",
103094=>"011011000",
103095=>"000001001",
103096=>"100000110",
103097=>"100001000",
103098=>"000000101",
103099=>"011111101",
103100=>"010000000",
103101=>"111001100",
103102=>"110001000",
103103=>"000000000",
103104=>"010110010",
103105=>"000000010",
103106=>"101011010",
103107=>"110100010",
103108=>"000000000",
103109=>"100110000",
103110=>"000110101",
103111=>"001000010",
103112=>"110101000",
103113=>"000100100",
103114=>"111100100",
103115=>"100000100",
103116=>"001000000",
103117=>"111110010",
103118=>"111000111",
103119=>"000001000",
103120=>"011110111",
103121=>"010111110",
103122=>"100100000",
103123=>"100100101",
103124=>"000000111",
103125=>"110100111",
103126=>"111001101",
103127=>"001001111",
103128=>"010010000",
103129=>"001001111",
103130=>"000010010",
103131=>"110000000",
103132=>"001011010",
103133=>"111011100",
103134=>"010111111",
103135=>"001100111",
103136=>"111000111",
103137=>"100000000",
103138=>"100010000",
103139=>"001000011",
103140=>"000000000",
103141=>"111001000",
103142=>"000101000",
103143=>"110110010",
103144=>"111101111",
103145=>"010000000",
103146=>"011010011",
103147=>"111000000",
103148=>"101001000",
103149=>"000000010",
103150=>"111101110",
103151=>"000000111",
103152=>"000000000",
103153=>"110011000",
103154=>"111110111",
103155=>"100110000",
103156=>"000110001",
103157=>"111011101",
103158=>"000000111",
103159=>"010011011",
103160=>"000010111",
103161=>"110010000",
103162=>"000010010",
103163=>"010011010",
103164=>"000010011",
103165=>"101100101",
103166=>"000001110",
103167=>"000111111",
103168=>"011000000",
103169=>"110110110",
103170=>"000000000",
103171=>"100100100",
103172=>"110010011",
103173=>"001100111",
103174=>"110110000",
103175=>"110101101",
103176=>"011111111",
103177=>"000000100",
103178=>"111111111",
103179=>"011010111",
103180=>"110101111",
103181=>"000000000",
103182=>"001101011",
103183=>"010010000",
103184=>"000110111",
103185=>"011011110",
103186=>"100010000",
103187=>"110110100",
103188=>"111111010",
103189=>"001101110",
103190=>"011100111",
103191=>"111110110",
103192=>"000000100",
103193=>"011000000",
103194=>"011011100",
103195=>"000010000",
103196=>"010001001",
103197=>"111011101",
103198=>"001100000",
103199=>"000111011",
103200=>"111011110",
103201=>"011011011",
103202=>"111111000",
103203=>"101111100",
103204=>"110101111",
103205=>"010100111",
103206=>"000001001",
103207=>"110110110",
103208=>"100011011",
103209=>"010010101",
103210=>"000100000",
103211=>"001001000",
103212=>"000101011",
103213=>"011100101",
103214=>"011000110",
103215=>"111111001",
103216=>"010000001",
103217=>"111011001",
103218=>"111101001",
103219=>"111010000",
103220=>"111111110",
103221=>"110100000",
103222=>"000000001",
103223=>"111101000",
103224=>"110000011",
103225=>"110100111",
103226=>"000100111",
103227=>"011100100",
103228=>"011000000",
103229=>"000011011",
103230=>"000000000",
103231=>"001001011",
103232=>"110111011",
103233=>"000000110",
103234=>"011111111",
103235=>"011110110",
103236=>"000010010",
103237=>"010000000",
103238=>"000000000",
103239=>"011011111",
103240=>"001101110",
103241=>"100100110",
103242=>"100100011",
103243=>"100010010",
103244=>"011000000",
103245=>"011001101",
103246=>"110110100",
103247=>"110011111",
103248=>"100001001",
103249=>"001010101",
103250=>"010000100",
103251=>"001000110",
103252=>"010010000",
103253=>"100111110",
103254=>"000001011",
103255=>"001000100",
103256=>"001111110",
103257=>"100101101",
103258=>"000000000",
103259=>"111001011",
103260=>"011110100",
103261=>"001001011",
103262=>"000110110",
103263=>"101101011",
103264=>"000011011",
103265=>"100000100",
103266=>"100100100",
103267=>"000000011",
103268=>"100100001",
103269=>"000110110",
103270=>"111110111",
103271=>"010001001",
103272=>"110000110",
103273=>"111100110",
103274=>"011010111",
103275=>"110110011",
103276=>"011111011",
103277=>"010011001",
103278=>"101111100",
103279=>"111011011",
103280=>"110110010",
103281=>"111101111",
103282=>"111110110",
103283=>"000001000",
103284=>"111000010",
103285=>"010100100",
103286=>"010000000",
103287=>"111001100",
103288=>"000000100",
103289=>"001010000",
103290=>"110000000",
103291=>"000000000",
103292=>"001001111",
103293=>"110100001",
103294=>"110100010",
103295=>"000001000",
103296=>"111000010",
103297=>"000000000",
103298=>"011011100",
103299=>"011111011",
103300=>"011010000",
103301=>"001010010",
103302=>"000000000",
103303=>"000000000",
103304=>"100101000",
103305=>"010000010",
103306=>"100000111",
103307=>"001000111",
103308=>"000001011",
103309=>"111111011",
103310=>"011111111",
103311=>"000000000",
103312=>"110100100",
103313=>"101011011",
103314=>"000000110",
103315=>"101110111",
103316=>"100001000",
103317=>"001000110",
103318=>"010010010",
103319=>"011111011",
103320=>"011111001",
103321=>"100110001",
103322=>"000010000",
103323=>"000000101",
103324=>"000011011",
103325=>"001011011",
103326=>"011110110",
103327=>"001001011",
103328=>"111100100",
103329=>"010111000",
103330=>"111110101",
103331=>"110000111",
103332=>"011110110",
103333=>"010110110",
103334=>"110000001",
103335=>"001010010",
103336=>"011000000",
103337=>"000110111",
103338=>"011001000",
103339=>"010100000",
103340=>"111111000",
103341=>"111111111",
103342=>"111111111",
103343=>"000100100",
103344=>"000000000",
103345=>"000000000",
103346=>"110111100",
103347=>"000100111",
103348=>"101100001",
103349=>"111100111",
103350=>"101001000",
103351=>"001001000",
103352=>"001010000",
103353=>"001000000",
103354=>"001000000",
103355=>"011111011",
103356=>"100100000",
103357=>"001111011",
103358=>"001001001",
103359=>"100000000",
103360=>"110010000",
103361=>"010000000",
103362=>"111000101",
103363=>"011101001",
103364=>"001100111",
103365=>"110000111",
103366=>"111111111",
103367=>"010001101",
103368=>"000001100",
103369=>"010010010",
103370=>"111001110",
103371=>"000000010",
103372=>"001000000",
103373=>"111111100",
103374=>"100111000",
103375=>"110110011",
103376=>"010010000",
103377=>"011101001",
103378=>"000001011",
103379=>"011111110",
103380=>"111011001",
103381=>"111111111",
103382=>"100000100",
103383=>"010000000",
103384=>"010100100",
103385=>"000000110",
103386=>"110110110",
103387=>"100000000",
103388=>"111001010",
103389=>"000001000",
103390=>"011010010",
103391=>"011010001",
103392=>"000111001",
103393=>"111100000",
103394=>"010110100",
103395=>"001000000",
103396=>"000000000",
103397=>"011001000",
103398=>"111001100",
103399=>"000000000",
103400=>"000001010",
103401=>"011011110",
103402=>"000000000",
103403=>"001011111",
103404=>"100101011",
103405=>"111111100",
103406=>"001011010",
103407=>"001000100",
103408=>"010010000",
103409=>"001111100",
103410=>"001000000",
103411=>"001101011",
103412=>"111111111",
103413=>"100101101",
103414=>"000000000",
103415=>"100110001",
103416=>"000110000",
103417=>"110100100",
103418=>"111111011",
103419=>"110110110",
103420=>"110111101",
103421=>"011011000",
103422=>"101111101",
103423=>"000010000",
103424=>"100100110",
103425=>"111111000",
103426=>"000000100",
103427=>"111010000",
103428=>"000000000",
103429=>"111111111",
103430=>"101000000",
103431=>"111111100",
103432=>"010011011",
103433=>"000000001",
103434=>"100001100",
103435=>"000000000",
103436=>"111111001",
103437=>"000111111",
103438=>"110100000",
103439=>"000000000",
103440=>"101110111",
103441=>"111100100",
103442=>"101000000",
103443=>"000000000",
103444=>"101000000",
103445=>"101101101",
103446=>"011000000",
103447=>"111111111",
103448=>"111010011",
103449=>"000110000",
103450=>"000000000",
103451=>"100111010",
103452=>"001000100",
103453=>"000101000",
103454=>"000100110",
103455=>"000000001",
103456=>"011101100",
103457=>"000010011",
103458=>"111101100",
103459=>"011000000",
103460=>"000100000",
103461=>"000000000",
103462=>"111000101",
103463=>"111001101",
103464=>"101100101",
103465=>"101101111",
103466=>"101000000",
103467=>"010111111",
103468=>"000101101",
103469=>"111110011",
103470=>"011101111",
103471=>"101000100",
103472=>"100100111",
103473=>"101110111",
103474=>"000000100",
103475=>"011101111",
103476=>"101000000",
103477=>"000110100",
103478=>"100100001",
103479=>"000000000",
103480=>"010111111",
103481=>"101101101",
103482=>"101000111",
103483=>"011000111",
103484=>"001000011",
103485=>"100111111",
103486=>"000000010",
103487=>"101010001",
103488=>"111111011",
103489=>"011000000",
103490=>"111001101",
103491=>"000001110",
103492=>"000111111",
103493=>"101100000",
103494=>"100111011",
103495=>"111111111",
103496=>"000111111",
103497=>"000000111",
103498=>"111111000",
103499=>"001000000",
103500=>"000001101",
103501=>"101111000",
103502=>"010111111",
103503=>"000001111",
103504=>"000100101",
103505=>"110111111",
103506=>"100001101",
103507=>"101000000",
103508=>"110000000",
103509=>"010101110",
103510=>"000000000",
103511=>"000000000",
103512=>"100111111",
103513=>"000000000",
103514=>"000110011",
103515=>"111111010",
103516=>"001011011",
103517=>"100110010",
103518=>"011111111",
103519=>"000000000",
103520=>"000001000",
103521=>"111111000",
103522=>"000110101",
103523=>"001111110",
103524=>"000000000",
103525=>"100000000",
103526=>"001100000",
103527=>"000101111",
103528=>"111010001",
103529=>"000000000",
103530=>"001000000",
103531=>"000010111",
103532=>"000000000",
103533=>"000111100",
103534=>"000000000",
103535=>"111111111",
103536=>"100111111",
103537=>"000000000",
103538=>"001001000",
103539=>"100000000",
103540=>"000101111",
103541=>"111110110",
103542=>"000000000",
103543=>"000000000",
103544=>"001010011",
103545=>"111111010",
103546=>"001110110",
103547=>"101000111",
103548=>"011001000",
103549=>"001011011",
103550=>"100111111",
103551=>"000001010",
103552=>"000010000",
103553=>"000000000",
103554=>"000001011",
103555=>"101000010",
103556=>"000000000",
103557=>"101010101",
103558=>"001000010",
103559=>"100000000",
103560=>"000111000",
103561=>"000100101",
103562=>"100000000",
103563=>"101010111",
103564=>"000011111",
103565=>"111111111",
103566=>"011000010",
103567=>"001000000",
103568=>"111010111",
103569=>"000101000",
103570=>"000000000",
103571=>"111011000",
103572=>"010000000",
103573=>"000001000",
103574=>"010111011",
103575=>"000000101",
103576=>"001000100",
103577=>"111011011",
103578=>"001111111",
103579=>"111000000",
103580=>"100000000",
103581=>"111111111",
103582=>"111000011",
103583=>"000000000",
103584=>"000001111",
103585=>"010111111",
103586=>"000011111",
103587=>"100001111",
103588=>"000011010",
103589=>"001100100",
103590=>"111101001",
103591=>"000000000",
103592=>"111010000",
103593=>"111000101",
103594=>"000111011",
103595=>"000010001",
103596=>"110111000",
103597=>"111100111",
103598=>"000011111",
103599=>"101111001",
103600=>"000000000",
103601=>"100110110",
103602=>"111000000",
103603=>"011011011",
103604=>"111111111",
103605=>"100000001",
103606=>"000101001",
103607=>"000111011",
103608=>"100100000",
103609=>"000000000",
103610=>"000001111",
103611=>"000000010",
103612=>"000000000",
103613=>"110111111",
103614=>"001111010",
103615=>"110000100",
103616=>"000000000",
103617=>"000101010",
103618=>"111111100",
103619=>"000001001",
103620=>"001000110",
103621=>"010010110",
103622=>"111111111",
103623=>"001111001",
103624=>"000110011",
103625=>"100000000",
103626=>"000000010",
103627=>"111000000",
103628=>"000000000",
103629=>"010100100",
103630=>"011111011",
103631=>"111111111",
103632=>"000111001",
103633=>"000110110",
103634=>"010111001",
103635=>"101100101",
103636=>"001000000",
103637=>"001011011",
103638=>"000000101",
103639=>"000010101",
103640=>"001000100",
103641=>"110111000",
103642=>"000000011",
103643=>"000010110",
103644=>"010011010",
103645=>"110110111",
103646=>"101000000",
103647=>"000100101",
103648=>"101000000",
103649=>"000011111",
103650=>"111011111",
103651=>"011011001",
103652=>"000000001",
103653=>"000000010",
103654=>"011001101",
103655=>"000111010",
103656=>"111111011",
103657=>"110111111",
103658=>"101100000",
103659=>"000000011",
103660=>"000011010",
103661=>"100100000",
103662=>"000111000",
103663=>"010000000",
103664=>"111100111",
103665=>"010000011",
103666=>"000000110",
103667=>"111011001",
103668=>"000001011",
103669=>"000010111",
103670=>"111010110",
103671=>"111010011",
103672=>"000000000",
103673=>"000011101",
103674=>"100000000",
103675=>"010010000",
103676=>"111111101",
103677=>"011010010",
103678=>"100000000",
103679=>"111001000",
103680=>"110011000",
103681=>"111111111",
103682=>"010111111",
103683=>"111101100",
103684=>"010010111",
103685=>"110111111",
103686=>"000000101",
103687=>"101000000",
103688=>"111000101",
103689=>"101100001",
103690=>"000000000",
103691=>"101101111",
103692=>"111111011",
103693=>"101101101",
103694=>"010000011",
103695=>"010100000",
103696=>"001000100",
103697=>"111101101",
103698=>"010011010",
103699=>"111000100",
103700=>"010111010",
103701=>"001010000",
103702=>"100011011",
103703=>"000000000",
103704=>"010111000",
103705=>"000001010",
103706=>"111101111",
103707=>"111010000",
103708=>"111111010",
103709=>"101110111",
103710=>"011111101",
103711=>"111000101",
103712=>"111111111",
103713=>"001111010",
103714=>"111101110",
103715=>"111111111",
103716=>"001000100",
103717=>"100000110",
103718=>"100101001",
103719=>"111000111",
103720=>"000100100",
103721=>"101101001",
103722=>"000000101",
103723=>"111111111",
103724=>"100000100",
103725=>"000011111",
103726=>"000000010",
103727=>"100001000",
103728=>"001101111",
103729=>"110010110",
103730=>"111101111",
103731=>"111111000",
103732=>"111111000",
103733=>"110001000",
103734=>"111110100",
103735=>"111010000",
103736=>"101101001",
103737=>"011011000",
103738=>"111111111",
103739=>"000000101",
103740=>"111111111",
103741=>"000000000",
103742=>"011111010",
103743=>"000000100",
103744=>"000000000",
103745=>"111101111",
103746=>"001001101",
103747=>"011011001",
103748=>"111101101",
103749=>"000010010",
103750=>"111111111",
103751=>"111111111",
103752=>"010000010",
103753=>"101100101",
103754=>"111111111",
103755=>"110110100",
103756=>"110111101",
103757=>"110000011",
103758=>"001000000",
103759=>"000011011",
103760=>"111101111",
103761=>"000010000",
103762=>"101000000",
103763=>"110100111",
103764=>"111111111",
103765=>"010000000",
103766=>"111100100",
103767=>"111101111",
103768=>"101101100",
103769=>"111000110",
103770=>"111011111",
103771=>"001000111",
103772=>"111000000",
103773=>"111111110",
103774=>"100111000",
103775=>"000110100",
103776=>"101101101",
103777=>"101101100",
103778=>"011111010",
103779=>"011010010",
103780=>"011000011",
103781=>"000000011",
103782=>"101000000",
103783=>"110000001",
103784=>"010010000",
103785=>"111000000",
103786=>"000000000",
103787=>"100101000",
103788=>"111011111",
103789=>"111110010",
103790=>"000011011",
103791=>"101111111",
103792=>"011001001",
103793=>"101001000",
103794=>"001011000",
103795=>"110111111",
103796=>"110100101",
103797=>"011111011",
103798=>"100100100",
103799=>"001100111",
103800=>"111101100",
103801=>"001000000",
103802=>"000000000",
103803=>"011011011",
103804=>"011011001",
103805=>"011011111",
103806=>"011111000",
103807=>"010111110",
103808=>"110111101",
103809=>"000001011",
103810=>"101000101",
103811=>"101000001",
103812=>"010001000",
103813=>"000001000",
103814=>"001001111",
103815=>"000010100",
103816=>"010000110",
103817=>"000001101",
103818=>"110000100",
103819=>"111111111",
103820=>"101111111",
103821=>"000000010",
103822=>"111011011",
103823=>"110111111",
103824=>"010000110",
103825=>"111001001",
103826=>"010111101",
103827=>"001101000",
103828=>"111100001",
103829=>"011001001",
103830=>"001010000",
103831=>"111100100",
103832=>"000001000",
103833=>"111101000",
103834=>"011011010",
103835=>"010111111",
103836=>"101101111",
103837=>"100100000",
103838=>"000101101",
103839=>"011011011",
103840=>"110110110",
103841=>"111111101",
103842=>"001000111",
103843=>"111111010",
103844=>"011001001",
103845=>"001100111",
103846=>"100101101",
103847=>"111000101",
103848=>"000000001",
103849=>"111101101",
103850=>"000011000",
103851=>"111111010",
103852=>"100111111",
103853=>"111001111",
103854=>"011011010",
103855=>"100000101",
103856=>"111011010",
103857=>"110001001",
103858=>"111111111",
103859=>"111111011",
103860=>"101000100",
103861=>"111111111",
103862=>"100000111",
103863=>"100111110",
103864=>"101111111",
103865=>"110000010",
103866=>"111000000",
103867=>"001100000",
103868=>"101100111",
103869=>"000111111",
103870=>"111001111",
103871=>"111101101",
103872=>"111111000",
103873=>"111000111",
103874=>"010101101",
103875=>"011101011",
103876=>"100101111",
103877=>"000110011",
103878=>"111100000",
103879=>"000010000",
103880=>"101100010",
103881=>"000010011",
103882=>"000111011",
103883=>"111110000",
103884=>"111000000",
103885=>"111111100",
103886=>"111101101",
103887=>"011000000",
103888=>"010111010",
103889=>"011001011",
103890=>"000111101",
103891=>"010010000",
103892=>"010011010",
103893=>"111111111",
103894=>"111111100",
103895=>"111101000",
103896=>"000000000",
103897=>"011001001",
103898=>"011011011",
103899=>"010111111",
103900=>"001000111",
103901=>"100100100",
103902=>"101101111",
103903=>"001001001",
103904=>"010011011",
103905=>"010111010",
103906=>"000000010",
103907=>"110001111",
103908=>"111101111",
103909=>"000111101",
103910=>"111111110",
103911=>"111101001",
103912=>"101101000",
103913=>"111111111",
103914=>"000010001",
103915=>"101101111",
103916=>"111111111",
103917=>"111111111",
103918=>"110110111",
103919=>"000010110",
103920=>"010010011",
103921=>"000110110",
103922=>"100101100",
103923=>"011001011",
103924=>"110000101",
103925=>"000110000",
103926=>"101111101",
103927=>"101101000",
103928=>"001111011",
103929=>"101101001",
103930=>"000111000",
103931=>"001101000",
103932=>"000000000",
103933=>"000000111",
103934=>"011001110",
103935=>"010010111",
103936=>"000000000",
103937=>"011000111",
103938=>"000000101",
103939=>"010000000",
103940=>"100110111",
103941=>"100100110",
103942=>"011000100",
103943=>"000000010",
103944=>"000111110",
103945=>"000101101",
103946=>"001001001",
103947=>"111111100",
103948=>"111111101",
103949=>"011101011",
103950=>"100111001",
103951=>"111011000",
103952=>"010000011",
103953=>"010111100",
103954=>"010100100",
103955=>"111100010",
103956=>"110111110",
103957=>"111100100",
103958=>"011100101",
103959=>"000010100",
103960=>"000000011",
103961=>"111111001",
103962=>"011111011",
103963=>"100100001",
103964=>"000000001",
103965=>"000100111",
103966=>"110000000",
103967=>"101111000",
103968=>"101101111",
103969=>"111111000",
103970=>"010011001",
103971=>"000111111",
103972=>"100110100",
103973=>"010010000",
103974=>"010011110",
103975=>"000001111",
103976=>"111011000",
103977=>"111000000",
103978=>"100100000",
103979=>"000010000",
103980=>"110101011",
103981=>"100000010",
103982=>"010010011",
103983=>"110111101",
103984=>"100111111",
103985=>"100110111",
103986=>"000110011",
103987=>"000000000",
103988=>"000000100",
103989=>"000000001",
103990=>"000000000",
103991=>"000000100",
103992=>"010010111",
103993=>"000000000",
103994=>"000000110",
103995=>"000101111",
103996=>"001000111",
103997=>"100111101",
103998=>"000101111",
103999=>"111000110",
104000=>"111111111",
104001=>"000000111",
104002=>"000000110",
104003=>"011001010",
104004=>"011111111",
104005=>"000000000",
104006=>"001001011",
104007=>"110011101",
104008=>"000111111",
104009=>"000111111",
104010=>"000011111",
104011=>"000000011",
104012=>"000100111",
104013=>"111111011",
104014=>"101001001",
104015=>"011011111",
104016=>"001000000",
104017=>"111100000",
104018=>"111011010",
104019=>"111100001",
104020=>"111010000",
104021=>"111100001",
104022=>"001001111",
104023=>"000000101",
104024=>"111110101",
104025=>"000011000",
104026=>"111111000",
104027=>"111011001",
104028=>"010111111",
104029=>"000001001",
104030=>"111011000",
104031=>"000000001",
104032=>"000000000",
104033=>"111100000",
104034=>"000000100",
104035=>"001011011",
104036=>"000100000",
104037=>"000110100",
104038=>"000111100",
104039=>"011001111",
104040=>"011111100",
104041=>"100000000",
104042=>"111100111",
104043=>"000101011",
104044=>"011111111",
104045=>"000010010",
104046=>"101101011",
104047=>"000000000",
104048=>"001011111",
104049=>"000000111",
104050=>"000100000",
104051=>"100000000",
104052=>"010110000",
104053=>"000000000",
104054=>"000001010",
104055=>"010010000",
104056=>"100000101",
104057=>"111111111",
104058=>"101111011",
104059=>"100110100",
104060=>"000100000",
104061=>"000100100",
104062=>"001111111",
104063=>"000000100",
104064=>"011011000",
104065=>"000100000",
104066=>"000111011",
104067=>"100101011",
104068=>"111000000",
104069=>"100100000",
104070=>"010001011",
104071=>"000011000",
104072=>"101001111",
104073=>"100000000",
104074=>"010111101",
104075=>"000001111",
104076=>"011000000",
104077=>"101011000",
104078=>"111011011",
104079=>"000000000",
104080=>"001101011",
104081=>"100111101",
104082=>"101111110",
104083=>"001010111",
104084=>"010110001",
104085=>"000000111",
104086=>"111000001",
104087=>"001001000",
104088=>"100111011",
104089=>"000000000",
104090=>"011011000",
104091=>"000000010",
104092=>"100000100",
104093=>"101111111",
104094=>"011100101",
104095=>"111010110",
104096=>"111100100",
104097=>"000000011",
104098=>"001111111",
104099=>"111111000",
104100=>"110101111",
104101=>"110111010",
104102=>"101000010",
104103=>"000000000",
104104=>"110000010",
104105=>"000010010",
104106=>"001111101",
104107=>"000011111",
104108=>"011011000",
104109=>"001101111",
104110=>"000001011",
104111=>"111011001",
104112=>"111111100",
104113=>"100010000",
104114=>"000100000",
104115=>"000100000",
104116=>"001011000",
104117=>"101110000",
104118=>"011111000",
104119=>"000000000",
104120=>"000001111",
104121=>"101110100",
104122=>"010001000",
104123=>"011011111",
104124=>"000001010",
104125=>"101101111",
104126=>"001001001",
104127=>"111110101",
104128=>"000000001",
104129=>"000000000",
104130=>"000101101",
104131=>"111110000",
104132=>"011000111",
104133=>"110001001",
104134=>"111100101",
104135=>"000100111",
104136=>"000001101",
104137=>"111011010",
104138=>"111010000",
104139=>"000000111",
104140=>"000000111",
104141=>"000000000",
104142=>"000000001",
104143=>"101101001",
104144=>"100101111",
104145=>"101101111",
104146=>"101111011",
104147=>"000010111",
104148=>"101111010",
104149=>"000100000",
104150=>"000000101",
104151=>"011011001",
104152=>"011011000",
104153=>"001000010",
104154=>"101101000",
104155=>"111001000",
104156=>"100000111",
104157=>"111111000",
104158=>"111111000",
104159=>"111000000",
104160=>"010111010",
104161=>"000000101",
104162=>"110000000",
104163=>"111110110",
104164=>"000000001",
104165=>"100000000",
104166=>"111111000",
104167=>"010000101",
104168=>"000000001",
104169=>"000100010",
104170=>"000000010",
104171=>"100000101",
104172=>"010010110",
104173=>"000000100",
104174=>"000000000",
104175=>"000100111",
104176=>"100111111",
104177=>"011000110",
104178=>"111000000",
104179=>"000111111",
104180=>"101100110",
104181=>"100001101",
104182=>"000000011",
104183=>"111001000",
104184=>"000010010",
104185=>"000011100",
104186=>"111010000",
104187=>"101100100",
104188=>"000001111",
104189=>"101010010",
104190=>"111111110",
104191=>"100000110",
104192=>"101101100",
104193=>"000000011",
104194=>"100100110",
104195=>"010010001",
104196=>"101101101",
104197=>"010010111",
104198=>"011011001",
104199=>"000001000",
104200=>"011000000",
104201=>"100100100",
104202=>"100010000",
104203=>"000000110",
104204=>"011010011",
104205=>"111111110",
104206=>"000110101",
104207=>"110111111",
104208=>"000000100",
104209=>"111110100",
104210=>"110110100",
104211=>"111001001",
104212=>"000100000",
104213=>"001101111",
104214=>"110100000",
104215=>"001001011",
104216=>"110100100",
104217=>"011100110",
104218=>"010110100",
104219=>"100100000",
104220=>"000000110",
104221=>"111010111",
104222=>"001111111",
104223=>"000000011",
104224=>"100100000",
104225=>"000000100",
104226=>"111110000",
104227=>"000000001",
104228=>"010110100",
104229=>"001110110",
104230=>"101001011",
104231=>"111111111",
104232=>"010011011",
104233=>"000001100",
104234=>"000001001",
104235=>"000100100",
104236=>"000010111",
104237=>"000000001",
104238=>"001111110",
104239=>"001010111",
104240=>"111111110",
104241=>"001111101",
104242=>"101000111",
104243=>"110110110",
104244=>"000000001",
104245=>"111011111",
104246=>"110110100",
104247=>"001011011",
104248=>"111110100",
104249=>"011000010",
104250=>"010110011",
104251=>"110100000",
104252=>"010010111",
104253=>"011011011",
104254=>"000100000",
104255=>"101001001",
104256=>"110100100",
104257=>"001101001",
104258=>"100011111",
104259=>"100111101",
104260=>"000000001",
104261=>"011000001",
104262=>"100001000",
104263=>"100100001",
104264=>"000001111",
104265=>"010000000",
104266=>"000000111",
104267=>"001001000",
104268=>"001001101",
104269=>"010110101",
104270=>"011011010",
104271=>"111110000",
104272=>"110101000",
104273=>"111110100",
104274=>"000000110",
104275=>"101100000",
104276=>"100101001",
104277=>"000011010",
104278=>"000010000",
104279=>"100000100",
104280=>"110110110",
104281=>"000010101",
104282=>"100010001",
104283=>"001111100",
104284=>"100100100",
104285=>"000100101",
104286=>"001011001",
104287=>"000011110",
104288=>"110110000",
104289=>"100011011",
104290=>"110100100",
104291=>"100000100",
104292=>"001011011",
104293=>"010010001",
104294=>"001000000",
104295=>"001011010",
104296=>"000011011",
104297=>"111110110",
104298=>"111010110",
104299=>"011000100",
104300=>"000101000",
104301=>"110100001",
104302=>"001100110",
104303=>"011000110",
104304=>"000001001",
104305=>"011111011",
104306=>"100100000",
104307=>"000100001",
104308=>"111000100",
104309=>"110100100",
104310=>"000101111",
104311=>"001001011",
104312=>"110100110",
104313=>"001100100",
104314=>"110000110",
104315=>"111011011",
104316=>"010001011",
104317=>"011010110",
104318=>"011011011",
104319=>"101100000",
104320=>"001011101",
104321=>"011110110",
104322=>"100100001",
104323=>"001000100",
104324=>"100100101",
104325=>"111111111",
104326=>"100100000",
104327=>"100010000",
104328=>"011011101",
104329=>"100111010",
104330=>"010110000",
104331=>"111001000",
104332=>"100101001",
104333=>"111100001",
104334=>"001010001",
104335=>"100000000",
104336=>"111011110",
104337=>"011000001",
104338=>"001001000",
104339=>"001111011",
104340=>"001111001",
104341=>"100100100",
104342=>"000000000",
104343=>"000000111",
104344=>"011010010",
104345=>"000110111",
104346=>"110110010",
104347=>"110100000",
104348=>"000001011",
104349=>"110111101",
104350=>"000110111",
104351=>"011011000",
104352=>"000010010",
104353=>"110100110",
104354=>"011011010",
104355=>"111111110",
104356=>"100110010",
104357=>"111101111",
104358=>"011011110",
104359=>"001001001",
104360=>"101100000",
104361=>"110110100",
104362=>"110110100",
104363=>"100100100",
104364=>"100100000",
104365=>"001011011",
104366=>"110010110",
104367=>"110000110",
104368=>"001011010",
104369=>"110100000",
104370=>"000010111",
104371=>"010100111",
104372=>"101111100",
104373=>"000000010",
104374=>"001111110",
104375=>"001111100",
104376=>"000001001",
104377=>"001001000",
104378=>"111011100",
104379=>"110110000",
104380=>"000110111",
104381=>"110110010",
104382=>"001010000",
104383=>"110000100",
104384=>"110110110",
104385=>"111100000",
104386=>"110001011",
104387=>"000101110",
104388=>"000001000",
104389=>"100100000",
104390=>"011111111",
104391=>"110101111",
104392=>"011010011",
104393=>"000101011",
104394=>"111101100",
104395=>"100000000",
104396=>"001001001",
104397=>"100000101",
104398=>"000100100",
104399=>"111110100",
104400=>"100111101",
104401=>"011110110",
104402=>"010001110",
104403=>"111111111",
104404=>"100111000",
104405=>"100000100",
104406=>"100110110",
104407=>"111010110",
104408=>"001011011",
104409=>"111011000",
104410=>"011101000",
104411=>"110100100",
104412=>"100111101",
104413=>"110100100",
104414=>"111110101",
104415=>"111011110",
104416=>"110000010",
104417=>"110110100",
104418=>"111011011",
104419=>"101111011",
104420=>"110100000",
104421=>"001011111",
104422=>"011001011",
104423=>"000001011",
104424=>"111111110",
104425=>"100101100",
104426=>"000000100",
104427=>"111100100",
104428=>"001001011",
104429=>"000011111",
104430=>"001000000",
104431=>"001000100",
104432=>"001011101",
104433=>"010110110",
104434=>"001001110",
104435=>"011111110",
104436=>"001011010",
104437=>"110100000",
104438=>"101100100",
104439=>"000000000",
104440=>"111100111",
104441=>"000111111",
104442=>"011110110",
104443=>"001011111",
104444=>"100011010",
104445=>"000111100",
104446=>"111111011",
104447=>"100000000",
104448=>"001100111",
104449=>"000000000",
104450=>"000000000",
104451=>"101101000",
104452=>"001011111",
104453=>"110000000",
104454=>"100010111",
104455=>"100000000",
104456=>"010011001",
104457=>"111000000",
104458=>"100000111",
104459=>"000000101",
104460=>"000000111",
104461=>"000000000",
104462=>"010101000",
104463=>"100111111",
104464=>"111000000",
104465=>"000000000",
104466=>"000101000",
104467=>"100000000",
104468=>"110000000",
104469=>"111000000",
104470=>"011111111",
104471=>"000110110",
104472=>"101000000",
104473=>"111011111",
104474=>"111111000",
104475=>"000000000",
104476=>"010111111",
104477=>"000001001",
104478=>"000000101",
104479=>"000000001",
104480=>"000011001",
104481=>"010000110",
104482=>"111111111",
104483=>"000010010",
104484=>"111010000",
104485=>"000111111",
104486=>"111001001",
104487=>"000000110",
104488=>"111101001",
104489=>"111111000",
104490=>"111110110",
104491=>"000101000",
104492=>"111111101",
104493=>"110110111",
104494=>"010000101",
104495=>"000000000",
104496=>"111111111",
104497=>"111111110",
104498=>"000010100",
104499=>"000000101",
104500=>"000100000",
104501=>"100010101",
104502=>"011100111",
104503=>"000000111",
104504=>"000111101",
104505=>"000000101",
104506=>"000100110",
104507=>"100111000",
104508=>"011010011",
104509=>"001000010",
104510=>"000000000",
104511=>"111011011",
104512=>"100000101",
104513=>"000011111",
104514=>"111000000",
104515=>"111111001",
104516=>"010000000",
104517=>"001000101",
104518=>"000000111",
104519=>"011000001",
104520=>"000100111",
104521=>"000000101",
104522=>"000000000",
104523=>"111010000",
104524=>"000001111",
104525=>"111111110",
104526=>"101110000",
104527=>"000101100",
104528=>"111000000",
104529=>"011000110",
104530=>"010001001",
104531=>"001100000",
104532=>"001000010",
104533=>"001000111",
104534=>"001000111",
104535=>"001101110",
104536=>"111111001",
104537=>"000010100",
104538=>"111110000",
104539=>"110110001",
104540=>"000001010",
104541=>"001111000",
104542=>"111011010",
104543=>"111100110",
104544=>"111111000",
104545=>"101000000",
104546=>"111000101",
104547=>"001001101",
104548=>"110111001",
104549=>"000011011",
104550=>"111100110",
104551=>"110101111",
104552=>"010111111",
104553=>"000011111",
104554=>"000001000",
104555=>"010000111",
104556=>"011111001",
104557=>"111111000",
104558=>"000000000",
104559=>"000101111",
104560=>"110100000",
104561=>"000010010",
104562=>"100100110",
104563=>"111101000",
104564=>"000000001",
104565=>"010000000",
104566=>"111111001",
104567=>"111001000",
104568=>"010100010",
104569=>"110000101",
104570=>"111010111",
104571=>"101101001",
104572=>"001001000",
104573=>"100101001",
104574=>"101111010",
104575=>"111111011",
104576=>"000111000",
104577=>"000000010",
104578=>"000000011",
104579=>"001000110",
104580=>"101000011",
104581=>"001111011",
104582=>"100111111",
104583=>"111000010",
104584=>"011001000",
104585=>"110000000",
104586=>"111010000",
104587=>"001000000",
104588=>"111001000",
104589=>"101110111",
104590=>"000000110",
104591=>"001000000",
104592=>"110100100",
104593=>"110111001",
104594=>"001111111",
104595=>"001000101",
104596=>"000000010",
104597=>"111001000",
104598=>"110110010",
104599=>"011111000",
104600=>"001111111",
104601=>"000100011",
104602=>"000000111",
104603=>"111000000",
104604=>"100000101",
104605=>"011001001",
104606=>"101111111",
104607=>"000001111",
104608=>"111100110",
104609=>"010000011",
104610=>"110000000",
104611=>"111000000",
104612=>"010000001",
104613=>"011111100",
104614=>"111010101",
104615=>"010011000",
104616=>"110000001",
104617=>"100111111",
104618=>"011110100",
104619=>"101000000",
104620=>"101111010",
104621=>"111000000",
104622=>"000110001",
104623=>"111001000",
104624=>"001111101",
104625=>"101110110",
104626=>"010010010",
104627=>"000001001",
104628=>"111111011",
104629=>"111111000",
104630=>"100000011",
104631=>"010110010",
104632=>"010010011",
104633=>"000000110",
104634=>"110000000",
104635=>"010111111",
104636=>"100110000",
104637=>"111101001",
104638=>"001000000",
104639=>"000000010",
104640=>"000001111",
104641=>"001101111",
104642=>"110111001",
104643=>"011000111",
104644=>"000010110",
104645=>"000001111",
104646=>"100111100",
104647=>"000000101",
104648=>"011011111",
104649=>"000001000",
104650=>"001000011",
104651=>"111000000",
104652=>"110000011",
104653=>"000000000",
104654=>"011101001",
104655=>"001000111",
104656=>"000000000",
104657=>"110110001",
104658=>"110000111",
104659=>"110111110",
104660=>"101000110",
104661=>"101001011",
104662=>"000000101",
104663=>"111010000",
104664=>"000111111",
104665=>"111000101",
104666=>"111001001",
104667=>"000000000",
104668=>"000110110",
104669=>"111111101",
104670=>"111111111",
104671=>"000111100",
104672=>"000000111",
104673=>"101000111",
104674=>"000111111",
104675=>"111011110",
104676=>"001001111",
104677=>"111000011",
104678=>"111111101",
104679=>"010110111",
104680=>"111100001",
104681=>"000000010",
104682=>"001000100",
104683=>"000001000",
104684=>"111000000",
104685=>"000011011",
104686=>"011000000",
104687=>"010101111",
104688=>"000000001",
104689=>"110000001",
104690=>"010000001",
104691=>"100000010",
104692=>"000001110",
104693=>"111111000",
104694=>"000000010",
104695=>"100000000",
104696=>"000000111",
104697=>"111111110",
104698=>"001000110",
104699=>"000001101",
104700=>"000010111",
104701=>"101001011",
104702=>"110111011",
104703=>"000000010",
104704=>"111000101",
104705=>"101111000",
104706=>"000000111",
104707=>"101101001",
104708=>"011000100",
104709=>"111100100",
104710=>"000101111",
104711=>"111011110",
104712=>"000000000",
104713=>"011110000",
104714=>"011010000",
104715=>"101010000",
104716=>"001001111",
104717=>"100000111",
104718=>"001001000",
104719=>"101000001",
104720=>"000010110",
104721=>"000000000",
104722=>"000000010",
104723=>"000010000",
104724=>"110010100",
104725=>"100101111",
104726=>"100100000",
104727=>"101111000",
104728=>"000010011",
104729=>"100010010",
104730=>"111011001",
104731=>"010011100",
104732=>"111111000",
104733=>"110110010",
104734=>"010001000",
104735=>"000001101",
104736=>"111001101",
104737=>"101010101",
104738=>"110000101",
104739=>"100111110",
104740=>"000100100",
104741=>"000100100",
104742=>"010000010",
104743=>"011111000",
104744=>"111010110",
104745=>"110110001",
104746=>"101111110",
104747=>"010110010",
104748=>"011011100",
104749=>"111010010",
104750=>"101111000",
104751=>"100110111",
104752=>"111010000",
104753=>"000001100",
104754=>"000010000",
104755=>"010010000",
104756=>"101000101",
104757=>"110000100",
104758=>"001001000",
104759=>"100010000",
104760=>"010100000",
104761=>"000000000",
104762=>"000101000",
104763=>"101111111",
104764=>"011101101",
104765=>"101100111",
104766=>"010000001",
104767=>"100100100",
104768=>"111111011",
104769=>"111000111",
104770=>"100111111",
104771=>"111110101",
104772=>"101101011",
104773=>"000000111",
104774=>"001000000",
104775=>"000111000",
104776=>"110110001",
104777=>"010100100",
104778=>"110100111",
104779=>"100101101",
104780=>"011000000",
104781=>"000101110",
104782=>"000110001",
104783=>"111111010",
104784=>"000001111",
104785=>"100101111",
104786=>"111010110",
104787=>"111100000",
104788=>"111111100",
104789=>"000000111",
104790=>"000001001",
104791=>"011111111",
104792=>"000010111",
104793=>"010111100",
104794=>"000100100",
104795=>"000110001",
104796=>"001011111",
104797=>"000001000",
104798=>"100101100",
104799=>"101001000",
104800=>"000000000",
104801=>"010001001",
104802=>"000000111",
104803=>"111111001",
104804=>"110001000",
104805=>"000001000",
104806=>"001000000",
104807=>"101100100",
104808=>"011000000",
104809=>"111101011",
104810=>"010010010",
104811=>"011101111",
104812=>"111011011",
104813=>"101000100",
104814=>"111111111",
104815=>"110010010",
104816=>"001100000",
104817=>"000010011",
104818=>"000110100",
104819=>"000000101",
104820=>"101111011",
104821=>"000001000",
104822=>"110011000",
104823=>"010100101",
104824=>"100100000",
104825=>"111101101",
104826=>"011011101",
104827=>"000001011",
104828=>"110110001",
104829=>"111100000",
104830=>"111110101",
104831=>"111000111",
104832=>"011000000",
104833=>"000001001",
104834=>"000001001",
104835=>"101101101",
104836=>"000010111",
104837=>"101100110",
104838=>"101001001",
104839=>"100011110",
104840=>"000101000",
104841=>"000000000",
104842=>"100100100",
104843=>"001111111",
104844=>"111000100",
104845=>"000001011",
104846=>"111111101",
104847=>"000001000",
104848=>"111110000",
104849=>"101000111",
104850=>"100000001",
104851=>"111000110",
104852=>"111011000",
104853=>"000010010",
104854=>"011111110",
104855=>"001001000",
104856=>"010010000",
104857=>"111110101",
104858=>"010000110",
104859=>"111001010",
104860=>"100100010",
104861=>"001000000",
104862=>"111010010",
104863=>"111011000",
104864=>"100000101",
104865=>"110010101",
104866=>"010111101",
104867=>"101000000",
104868=>"011111110",
104869=>"000000111",
104870=>"000100111",
104871=>"000111010",
104872=>"001010010",
104873=>"100111000",
104874=>"111000111",
104875=>"000001000",
104876=>"011111111",
104877=>"000100101",
104878=>"011100101",
104879=>"010110111",
104880=>"101000111",
104881=>"001011001",
104882=>"101101000",
104883=>"100100001",
104884=>"110000111",
104885=>"001101000",
104886=>"000100100",
104887=>"010111001",
104888=>"000001101",
104889=>"111110001",
104890=>"001000010",
104891=>"010010000",
104892=>"000100111",
104893=>"110000000",
104894=>"001000101",
104895=>"010010111",
104896=>"000101100",
104897=>"000000001",
104898=>"100100000",
104899=>"100000100",
104900=>"000100101",
104901=>"111110111",
104902=>"111011101",
104903=>"100101100",
104904=>"000000011",
104905=>"111101101",
104906=>"111101011",
104907=>"001000000",
104908=>"000000000",
104909=>"011001100",
104910=>"010111111",
104911=>"111110111",
104912=>"000101111",
104913=>"101110101",
104914=>"100010010",
104915=>"100100101",
104916=>"011011111",
104917=>"000110001",
104918=>"011011101",
104919=>"001011010",
104920=>"101001011",
104921=>"010011000",
104922=>"011111100",
104923=>"111000111",
104924=>"011001100",
104925=>"111101111",
104926=>"000010000",
104927=>"001110110",
104928=>"001101111",
104929=>"010000101",
104930=>"111001111",
104931=>"100100000",
104932=>"010000000",
104933=>"111101000",
104934=>"000011000",
104935=>"110110111",
104936=>"100000011",
104937=>"001011111",
104938=>"110000111",
104939=>"010110100",
104940=>"000000110",
104941=>"000100111",
104942=>"000000000",
104943=>"011000000",
104944=>"000000000",
104945=>"111111111",
104946=>"111011101",
104947=>"011001000",
104948=>"101001100",
104949=>"001111110",
104950=>"000001011",
104951=>"111011000",
104952=>"010010000",
104953=>"011001000",
104954=>"101001111",
104955=>"110111001",
104956=>"000000000",
104957=>"111110000",
104958=>"010001001",
104959=>"011001001",
104960=>"111011100",
104961=>"000100111",
104962=>"101000000",
104963=>"000000000",
104964=>"000101011",
104965=>"110000101",
104966=>"111101111",
104967=>"011010111",
104968=>"111101011",
104969=>"000000000",
104970=>"000000001",
104971=>"111111000",
104972=>"000000000",
104973=>"111100000",
104974=>"110100111",
104975=>"010000111",
104976=>"011000111",
104977=>"010000111",
104978=>"000111111",
104979=>"010000000",
104980=>"110010110",
104981=>"101000000",
104982=>"000000010",
104983=>"000100010",
104984=>"111000001",
104985=>"110111101",
104986=>"110101111",
104987=>"000011011",
104988=>"111111101",
104989=>"000101111",
104990=>"101100000",
104991=>"000000111",
104992=>"001111100",
104993=>"110010111",
104994=>"000000100",
104995=>"000000110",
104996=>"000000100",
104997=>"011001100",
104998=>"011001101",
104999=>"011111000",
105000=>"111000111",
105001=>"111000000",
105002=>"010110010",
105003=>"010111111",
105004=>"011000101",
105005=>"001101101",
105006=>"001000000",
105007=>"010000011",
105008=>"111101011",
105009=>"100100110",
105010=>"110010010",
105011=>"000111110",
105012=>"000000000",
105013=>"111111001",
105014=>"100100011",
105015=>"000010010",
105016=>"111110010",
105017=>"000010000",
105018=>"010010100",
105019=>"001100111",
105020=>"110011011",
105021=>"111111110",
105022=>"110100100",
105023=>"111001001",
105024=>"111101000",
105025=>"001000000",
105026=>"000000010",
105027=>"101100111",
105028=>"010111010",
105029=>"000010010",
105030=>"010100101",
105031=>"111000111",
105032=>"100000011",
105033=>"111000001",
105034=>"000001000",
105035=>"111000000",
105036=>"100110100",
105037=>"100111011",
105038=>"000011011",
105039=>"100111000",
105040=>"000000000",
105041=>"111011100",
105042=>"111111000",
105043=>"011011001",
105044=>"101000010",
105045=>"100100100",
105046=>"000000011",
105047=>"111000101",
105048=>"111101001",
105049=>"000001001",
105050=>"100110111",
105051=>"011110010",
105052=>"000111000",
105053=>"010000001",
105054=>"011010011",
105055=>"001000101",
105056=>"111110111",
105057=>"000000001",
105058=>"111000000",
105059=>"000010000",
105060=>"000101010",
105061=>"011111100",
105062=>"100000000",
105063=>"010011101",
105064=>"101010110",
105065=>"010000000",
105066=>"110100000",
105067=>"000001110",
105068=>"000000100",
105069=>"000111010",
105070=>"000000001",
105071=>"101001101",
105072=>"010000001",
105073=>"000000000",
105074=>"001001111",
105075=>"010000000",
105076=>"111000011",
105077=>"001000101",
105078=>"000111010",
105079=>"111000001",
105080=>"001000001",
105081=>"000111111",
105082=>"000100010",
105083=>"000000000",
105084=>"100011011",
105085=>"110100100",
105086=>"000000000",
105087=>"101101111",
105088=>"010011000",
105089=>"111000000",
105090=>"111101000",
105091=>"000000000",
105092=>"010000000",
105093=>"110110000",
105094=>"100101001",
105095=>"001100110",
105096=>"000000100",
105097=>"100111011",
105098=>"011111010",
105099=>"000000100",
105100=>"111101101",
105101=>"010111100",
105102=>"000010110",
105103=>"000000101",
105104=>"000100011",
105105=>"111100101",
105106=>"110110000",
105107=>"110111111",
105108=>"000010101",
105109=>"000000000",
105110=>"000000111",
105111=>"100100110",
105112=>"000010011",
105113=>"001001001",
105114=>"000111000",
105115=>"000000000",
105116=>"000100101",
105117=>"111011001",
105118=>"111111101",
105119=>"000000000",
105120=>"000000111",
105121=>"001000000",
105122=>"000100011",
105123=>"001000000",
105124=>"100111111",
105125=>"110110110",
105126=>"001101111",
105127=>"000110111",
105128=>"111010000",
105129=>"000010110",
105130=>"101000101",
105131=>"110000010",
105132=>"001111111",
105133=>"111001000",
105134=>"000001011",
105135=>"001111000",
105136=>"111000001",
105137=>"100101111",
105138=>"111011000",
105139=>"000000000",
105140=>"000111111",
105141=>"100101111",
105142=>"000011111",
105143=>"010111111",
105144=>"011110100",
105145=>"000111011",
105146=>"010000100",
105147=>"100010010",
105148=>"111000111",
105149=>"111111111",
105150=>"011101111",
105151=>"000000000",
105152=>"000000000",
105153=>"111101000",
105154=>"100101111",
105155=>"001001111",
105156=>"000011011",
105157=>"100101111",
105158=>"000000011",
105159=>"011000000",
105160=>"000000101",
105161=>"000000110",
105162=>"010111111",
105163=>"000101111",
105164=>"000000100",
105165=>"000110110",
105166=>"000000000",
105167=>"010111111",
105168=>"111111000",
105169=>"110000110",
105170=>"010111101",
105171=>"101111111",
105172=>"110011010",
105173=>"001101101",
105174=>"001000110",
105175=>"111100111",
105176=>"010111010",
105177=>"000011010",
105178=>"011001010",
105179=>"001000100",
105180=>"001000011",
105181=>"111111100",
105182=>"000010000",
105183=>"101100011",
105184=>"000000011",
105185=>"111000000",
105186=>"111101100",
105187=>"111001011",
105188=>"110000000",
105189=>"010001101",
105190=>"000101000",
105191=>"000101110",
105192=>"111110000",
105193=>"111111100",
105194=>"000000100",
105195=>"000000111",
105196=>"000011111",
105197=>"111111000",
105198=>"100000000",
105199=>"000000111",
105200=>"111111010",
105201=>"001001101",
105202=>"000111101",
105203=>"110110111",
105204=>"110100100",
105205=>"000001000",
105206=>"000110000",
105207=>"000000001",
105208=>"010010010",
105209=>"101000000",
105210=>"111111000",
105211=>"000111111",
105212=>"110010010",
105213=>"011111111",
105214=>"011110111",
105215=>"001110101",
105216=>"000001101",
105217=>"111100100",
105218=>"111000000",
105219=>"001000000",
105220=>"001010001",
105221=>"111011010",
105222=>"010000000",
105223=>"100100110",
105224=>"100010111",
105225=>"000000100",
105226=>"100100110",
105227=>"000001100",
105228=>"100111111",
105229=>"111000000",
105230=>"100011000",
105231=>"010000000",
105232=>"001010111",
105233=>"111011001",
105234=>"010001000",
105235=>"011111101",
105236=>"001000011",
105237=>"100001111",
105238=>"001011011",
105239=>"101111010",
105240=>"111101101",
105241=>"100001100",
105242=>"110111111",
105243=>"111000100",
105244=>"010111100",
105245=>"000000000",
105246=>"011101011",
105247=>"000000010",
105248=>"110000000",
105249=>"111100101",
105250=>"000000000",
105251=>"000011011",
105252=>"000100100",
105253=>"100100001",
105254=>"000000110",
105255=>"000010111",
105256=>"111001111",
105257=>"111111101",
105258=>"000000001",
105259=>"000111001",
105260=>"100110110",
105261=>"000000111",
105262=>"000100101",
105263=>"010000000",
105264=>"000000010",
105265=>"111001001",
105266=>"000101110",
105267=>"111000000",
105268=>"000101000",
105269=>"110000001",
105270=>"000110101",
105271=>"111001000",
105272=>"100000000",
105273=>"111101001",
105274=>"010111010",
105275=>"010010111",
105276=>"101111111",
105277=>"111011010",
105278=>"100000100",
105279=>"110010010",
105280=>"111100010",
105281=>"100111010",
105282=>"100100000",
105283=>"010110011",
105284=>"011110111",
105285=>"111001000",
105286=>"000010011",
105287=>"010011000",
105288=>"100011011",
105289=>"010010101",
105290=>"111101101",
105291=>"111101101",
105292=>"111101000",
105293=>"001000000",
105294=>"100100000",
105295=>"001001011",
105296=>"101101101",
105297=>"011000001",
105298=>"011010111",
105299=>"000011001",
105300=>"000000000",
105301=>"011110110",
105302=>"000011011",
105303=>"000010111",
105304=>"100100100",
105305=>"000011001",
105306=>"110110110",
105307=>"000011011",
105308=>"100000101",
105309=>"110001001",
105310=>"111100101",
105311=>"000011111",
105312=>"000010000",
105313=>"000001111",
105314=>"000100100",
105315=>"101001101",
105316=>"111101001",
105317=>"011011010",
105318=>"000010111",
105319=>"111000000",
105320=>"111110001",
105321=>"111100010",
105322=>"101100010",
105323=>"111111111",
105324=>"010001000",
105325=>"000000000",
105326=>"111100000",
105327=>"101101111",
105328=>"100001100",
105329=>"111100110",
105330=>"000001101",
105331=>"000010011",
105332=>"001111010",
105333=>"111000100",
105334=>"111100100",
105335=>"110100100",
105336=>"000000000",
105337=>"010111111",
105338=>"010000100",
105339=>"100001001",
105340=>"010111010",
105341=>"110110100",
105342=>"101000000",
105343=>"010010010",
105344=>"010010010",
105345=>"010110010",
105346=>"000000000",
105347=>"000111111",
105348=>"000000000",
105349=>"000111110",
105350=>"001011011",
105351=>"000001001",
105352=>"111110110",
105353=>"101100100",
105354=>"101001111",
105355=>"010011010",
105356=>"111000000",
105357=>"000000000",
105358=>"111000000",
105359=>"100000000",
105360=>"101100101",
105361=>"010001000",
105362=>"111000000",
105363=>"100000000",
105364=>"000011010",
105365=>"110111111",
105366=>"111101101",
105367=>"001101000",
105368=>"000000000",
105369=>"101100000",
105370=>"000000010",
105371=>"000000000",
105372=>"000110101",
105373=>"111100000",
105374=>"111111000",
105375=>"000010011",
105376=>"011111011",
105377=>"111011110",
105378=>"000111101",
105379=>"011110000",
105380=>"001100101",
105381=>"100110110",
105382=>"000110110",
105383=>"111000000",
105384=>"000111000",
105385=>"100101111",
105386=>"111110100",
105387=>"111000000",
105388=>"011010010",
105389=>"111100000",
105390=>"110110111",
105391=>"000000100",
105392=>"111101000",
105393=>"011000100",
105394=>"101101101",
105395=>"000110110",
105396=>"011011011",
105397=>"000000100",
105398=>"000000100",
105399=>"100000000",
105400=>"100000111",
105401=>"100110010",
105402=>"101110100",
105403=>"111111001",
105404=>"000010111",
105405=>"110000000",
105406=>"001000000",
105407=>"000101011",
105408=>"000000000",
105409=>"101101000",
105410=>"111000000",
105411=>"001110010",
105412=>"000000011",
105413=>"100100000",
105414=>"000110011",
105415=>"000000010",
105416=>"000111111",
105417=>"100010010",
105418=>"101101001",
105419=>"111101101",
105420=>"111100000",
105421=>"111110110",
105422=>"001101000",
105423=>"001000100",
105424=>"111000000",
105425=>"110111011",
105426=>"100100000",
105427=>"000101001",
105428=>"010010000",
105429=>"111001101",
105430=>"000111111",
105431=>"110011000",
105432=>"000011010",
105433=>"101000011",
105434=>"111111010",
105435=>"110010101",
105436=>"000011111",
105437=>"000001111",
105438=>"000000000",
105439=>"111010010",
105440=>"101000000",
105441=>"111100101",
105442=>"100000000",
105443=>"000101110",
105444=>"101100000",
105445=>"000111000",
105446=>"000000011",
105447=>"000010011",
105448=>"000100110",
105449=>"000011111",
105450=>"000001001",
105451=>"101101000",
105452=>"111000000",
105453=>"000100001",
105454=>"000000001",
105455=>"100000000",
105456=>"010011111",
105457=>"001011001",
105458=>"000010000",
105459=>"000110010",
105460=>"101100000",
105461=>"101101100",
105462=>"000000000",
105463=>"001111001",
105464=>"000010111",
105465=>"000111100",
105466=>"010000001",
105467=>"000100001",
105468=>"101100010",
105469=>"000000000",
105470=>"000001011",
105471=>"111000000",
105472=>"011011101",
105473=>"111110010",
105474=>"101000000",
105475=>"110100000",
105476=>"000001001",
105477=>"111111000",
105478=>"010001011",
105479=>"110111101",
105480=>"000110000",
105481=>"111111111",
105482=>"000110111",
105483=>"010111010",
105484=>"111000101",
105485=>"000000000",
105486=>"101011001",
105487=>"000101000",
105488=>"000010110",
105489=>"111000011",
105490=>"000000000",
105491=>"011001111",
105492=>"101011111",
105493=>"101000000",
105494=>"000010001",
105495=>"111000010",
105496=>"000000000",
105497=>"100000000",
105498=>"000010111",
105499=>"000110111",
105500=>"111001110",
105501=>"010010001",
105502=>"111111000",
105503=>"000000000",
105504=>"100111111",
105505=>"010010010",
105506=>"001000000",
105507=>"000111111",
105508=>"001111011",
105509=>"101100100",
105510=>"001101101",
105511=>"111101111",
105512=>"111111111",
105513=>"000010110",
105514=>"001101001",
105515=>"010000000",
105516=>"010000100",
105517=>"000001000",
105518=>"111101111",
105519=>"110110000",
105520=>"111010010",
105521=>"011111011",
105522=>"010000000",
105523=>"100001101",
105524=>"110111111",
105525=>"101110111",
105526=>"110110011",
105527=>"000010000",
105528=>"010000000",
105529=>"111111111",
105530=>"101000000",
105531=>"111100101",
105532=>"100110100",
105533=>"111001000",
105534=>"000000111",
105535=>"000011011",
105536=>"111111111",
105537=>"101111000",
105538=>"111101110",
105539=>"001111011",
105540=>"000101001",
105541=>"000001000",
105542=>"000011110",
105543=>"000000000",
105544=>"000000000",
105545=>"000000000",
105546=>"111101001",
105547=>"111111111",
105548=>"110000000",
105549=>"000011001",
105550=>"001100110",
105551=>"001000000",
105552=>"000000101",
105553=>"111000000",
105554=>"000000101",
105555=>"011001100",
105556=>"011111000",
105557=>"011100111",
105558=>"000100100",
105559=>"000000000",
105560=>"100101000",
105561=>"110100100",
105562=>"000100100",
105563=>"101100101",
105564=>"110111000",
105565=>"001001001",
105566=>"110111111",
105567=>"100110111",
105568=>"000100000",
105569=>"000111111",
105570=>"111101000",
105571=>"000111101",
105572=>"101110101",
105573=>"001001011",
105574=>"000000000",
105575=>"000010000",
105576=>"010111111",
105577=>"000000010",
105578=>"010110000",
105579=>"100000000",
105580=>"111000111",
105581=>"111111111",
105582=>"000000000",
105583=>"101000000",
105584=>"000110100",
105585=>"110100111",
105586=>"011011110",
105587=>"000101111",
105588=>"011111111",
105589=>"111000000",
105590=>"000011111",
105591=>"111001000",
105592=>"100010010",
105593=>"111011000",
105594=>"011001011",
105595=>"100000000",
105596=>"001110110",
105597=>"110100000",
105598=>"111100001",
105599=>"000010111",
105600=>"101001000",
105601=>"111100000",
105602=>"011001001",
105603=>"110010000",
105604=>"010111101",
105605=>"000000000",
105606=>"111001000",
105607=>"000001001",
105608=>"000001001",
105609=>"111001000",
105610=>"000111111",
105611=>"000000000",
105612=>"000110010",
105613=>"100010111",
105614=>"101101100",
105615=>"101001000",
105616=>"001100101",
105617=>"001100101",
105618=>"111111011",
105619=>"000001010",
105620=>"000011111",
105621=>"111010010",
105622=>"100111010",
105623=>"010011001",
105624=>"111111110",
105625=>"000000001",
105626=>"111001000",
105627=>"100000110",
105628=>"001001110",
105629=>"101111101",
105630=>"101000010",
105631=>"000000000",
105632=>"011000000",
105633=>"011010010",
105634=>"111000000",
105635=>"000000000",
105636=>"001101111",
105637=>"111001100",
105638=>"010000101",
105639=>"000010110",
105640=>"111111000",
105641=>"000000000",
105642=>"011011101",
105643=>"000100000",
105644=>"000010100",
105645=>"000111001",
105646=>"110110101",
105647=>"111101001",
105648=>"000111000",
105649=>"000000000",
105650=>"001111000",
105651=>"000100100",
105652=>"001100001",
105653=>"111000101",
105654=>"000001000",
105655=>"000010110",
105656=>"000001011",
105657=>"000100110",
105658=>"000000000",
105659=>"110000010",
105660=>"010111000",
105661=>"111110110",
105662=>"100100111",
105663=>"000000000",
105664=>"000000000",
105665=>"111000000",
105666=>"111000000",
105667=>"001011101",
105668=>"001001000",
105669=>"100001000",
105670=>"000000011",
105671=>"010111000",
105672=>"000110011",
105673=>"000000001",
105674=>"000000000",
105675=>"111010000",
105676=>"000000010",
105677=>"000011011",
105678=>"000010010",
105679=>"100101011",
105680=>"000010010",
105681=>"000110100",
105682=>"000000010",
105683=>"100011010",
105684=>"101000000",
105685=>"000110000",
105686=>"000110110",
105687=>"111100000",
105688=>"111000000",
105689=>"000000101",
105690=>"100000000",
105691=>"011000000",
105692=>"100001110",
105693=>"000000000",
105694=>"111000000",
105695=>"000010110",
105696=>"000000000",
105697=>"101000000",
105698=>"000100100",
105699=>"001111111",
105700=>"000000110",
105701=>"000111111",
105702=>"111001111",
105703=>"111101111",
105704=>"010000000",
105705=>"000010001",
105706=>"011111111",
105707=>"000101110",
105708=>"100000111",
105709=>"000110000",
105710=>"010000000",
105711=>"010001101",
105712=>"111111111",
105713=>"101111100",
105714=>"111000000",
105715=>"000001001",
105716=>"000100011",
105717=>"000001101",
105718=>"000010000",
105719=>"010000000",
105720=>"111000000",
105721=>"001011111",
105722=>"110010000",
105723=>"100111011",
105724=>"001001101",
105725=>"010011111",
105726=>"110110100",
105727=>"111001000",
105728=>"110001001",
105729=>"101111111",
105730=>"101000111",
105731=>"110000000",
105732=>"100010011",
105733=>"000000010",
105734=>"000011111",
105735=>"110011001",
105736=>"000001001",
105737=>"000000000",
105738=>"010010110",
105739=>"000110010",
105740=>"000000010",
105741=>"010000000",
105742=>"001011110",
105743=>"011001000",
105744=>"111111111",
105745=>"111000111",
105746=>"111101000",
105747=>"111011000",
105748=>"000110111",
105749=>"111001001",
105750=>"011000001",
105751=>"111111100",
105752=>"001001101",
105753=>"001010111",
105754=>"000100101",
105755=>"000011111",
105756=>"000100010",
105757=>"000111111",
105758=>"100000110",
105759=>"011101101",
105760=>"001000111",
105761=>"000110111",
105762=>"111111101",
105763=>"111111000",
105764=>"000011011",
105765=>"101000001",
105766=>"111010110",
105767=>"000000000",
105768=>"111111111",
105769=>"111111101",
105770=>"001000000",
105771=>"010010010",
105772=>"000100011",
105773=>"011111111",
105774=>"100000000",
105775=>"001110101",
105776=>"110000111",
105777=>"110001001",
105778=>"000010001",
105779=>"101100110",
105780=>"000000000",
105781=>"110111101",
105782=>"110100001",
105783=>"111111101",
105784=>"010010110",
105785=>"101001101",
105786=>"100111111",
105787=>"111001101",
105788=>"010100011",
105789=>"010000111",
105790=>"000000111",
105791=>"111001100",
105792=>"101101101",
105793=>"100000000",
105794=>"000000000",
105795=>"001100011",
105796=>"000000000",
105797=>"111011101",
105798=>"000010110",
105799=>"011000101",
105800=>"111100001",
105801=>"000111111",
105802=>"111101101",
105803=>"000000000",
105804=>"111101100",
105805=>"000110110",
105806=>"101010000",
105807=>"010110111",
105808=>"000000111",
105809=>"010010110",
105810=>"000000111",
105811=>"000001001",
105812=>"100000010",
105813=>"001110111",
105814=>"001100100",
105815=>"111111111",
105816=>"111001111",
105817=>"001111010",
105818=>"111100000",
105819=>"000000100",
105820=>"010000000",
105821=>"001100101",
105822=>"000101000",
105823=>"000000100",
105824=>"101001000",
105825=>"000010010",
105826=>"000000000",
105827=>"111001001",
105828=>"010100111",
105829=>"000000001",
105830=>"000110111",
105831=>"111001001",
105832=>"010000000",
105833=>"000111111",
105834=>"111111101",
105835=>"011000000",
105836=>"000000000",
105837=>"110111111",
105838=>"111010010",
105839=>"000111111",
105840=>"100100110",
105841=>"000101010",
105842=>"011000000",
105843=>"111000000",
105844=>"111111101",
105845=>"000000001",
105846=>"000110111",
105847=>"101111001",
105848=>"010011101",
105849=>"010111001",
105850=>"000000001",
105851=>"010010111",
105852=>"101100100",
105853=>"011001010",
105854=>"000000111",
105855=>"000000111",
105856=>"110000000",
105857=>"111110110",
105858=>"011110000",
105859=>"001000110",
105860=>"010011000",
105861=>"111101101",
105862=>"111000000",
105863=>"001000000",
105864=>"011001011",
105865=>"100001110",
105866=>"011010111",
105867=>"111010011",
105868=>"010111111",
105869=>"001010111",
105870=>"111111001",
105871=>"000001000",
105872=>"110100100",
105873=>"110001101",
105874=>"011101010",
105875=>"000000000",
105876=>"000000010",
105877=>"101000111",
105878=>"010001000",
105879=>"011111100",
105880=>"101011001",
105881=>"000010010",
105882=>"110000000",
105883=>"000000000",
105884=>"000000111",
105885=>"001001010",
105886=>"110000000",
105887=>"111000000",
105888=>"111111100",
105889=>"100100000",
105890=>"001010011",
105891=>"101011000",
105892=>"000000000",
105893=>"110100000",
105894=>"111111001",
105895=>"001000111",
105896=>"000000000",
105897=>"111111101",
105898=>"001000000",
105899=>"000000010",
105900=>"011111010",
105901=>"000010111",
105902=>"000001000",
105903=>"111000010",
105904=>"111001000",
105905=>"001101001",
105906=>"000000010",
105907=>"000101110",
105908=>"010010010",
105909=>"010000000",
105910=>"111111100",
105911=>"000000000",
105912=>"011001010",
105913=>"101100001",
105914=>"000000111",
105915=>"011000101",
105916=>"010000011",
105917=>"011111111",
105918=>"111100000",
105919=>"000010011",
105920=>"000000000",
105921=>"100000000",
105922=>"001011000",
105923=>"100011011",
105924=>"000000000",
105925=>"000111010",
105926=>"000000000",
105927=>"111000000",
105928=>"001110111",
105929=>"111101000",
105930=>"101011101",
105931=>"111101001",
105932=>"011100100",
105933=>"001001000",
105934=>"010101101",
105935=>"111000000",
105936=>"111011000",
105937=>"111001001",
105938=>"001000101",
105939=>"011111101",
105940=>"000000000",
105941=>"111111111",
105942=>"100010000",
105943=>"111111101",
105944=>"111110100",
105945=>"000101101",
105946=>"100101000",
105947=>"000100000",
105948=>"000001001",
105949=>"111000000",
105950=>"011000000",
105951=>"011000000",
105952=>"000000111",
105953=>"100110111",
105954=>"111011011",
105955=>"110110111",
105956=>"001101100",
105957=>"000011011",
105958=>"000000000",
105959=>"111111000",
105960=>"000000110",
105961=>"010000100",
105962=>"000010111",
105963=>"101000000",
105964=>"000010111",
105965=>"111010000",
105966=>"000000010",
105967=>"111110100",
105968=>"111101100",
105969=>"000110111",
105970=>"111011101",
105971=>"100100100",
105972=>"101110101",
105973=>"001101111",
105974=>"000101000",
105975=>"000000000",
105976=>"000000110",
105977=>"111010000",
105978=>"000110000",
105979=>"101001011",
105980=>"111101100",
105981=>"000111010",
105982=>"001110110",
105983=>"000111111",
105984=>"000100100",
105985=>"010000010",
105986=>"010100100",
105987=>"100110010",
105988=>"011111000",
105989=>"000100111",
105990=>"101000010",
105991=>"111000101",
105992=>"010000000",
105993=>"000000000",
105994=>"100110001",
105995=>"000100000",
105996=>"000000000",
105997=>"001010111",
105998=>"111100001",
105999=>"111101000",
106000=>"101101000",
106001=>"000000000",
106002=>"101101101",
106003=>"110110001",
106004=>"111000010",
106005=>"011111111",
106006=>"101100101",
106007=>"101101101",
106008=>"000001000",
106009=>"001000000",
106010=>"111010000",
106011=>"100000000",
106012=>"001101111",
106013=>"000011111",
106014=>"000000000",
106015=>"111000111",
106016=>"000100101",
106017=>"111011000",
106018=>"100100111",
106019=>"000000100",
106020=>"111101100",
106021=>"000001110",
106022=>"000000111",
106023=>"110101111",
106024=>"111111111",
106025=>"100101101",
106026=>"001101101",
106027=>"000001000",
106028=>"000101100",
106029=>"100110110",
106030=>"010010011",
106031=>"000001000",
106032=>"011111010",
106033=>"111100000",
106034=>"100000110",
106035=>"111111101",
106036=>"000100100",
106037=>"111101001",
106038=>"000000101",
106039=>"010010011",
106040=>"111010001",
106041=>"110110110",
106042=>"100101101",
106043=>"001011101",
106044=>"110111111",
106045=>"111111110",
106046=>"000000000",
106047=>"011011000",
106048=>"000000001",
106049=>"010000100",
106050=>"111111011",
106051=>"110100000",
106052=>"010010111",
106053=>"000000000",
106054=>"010110100",
106055=>"000100010",
106056=>"011011000",
106057=>"010001001",
106058=>"001000010",
106059=>"101111000",
106060=>"111110001",
106061=>"111001001",
106062=>"110111000",
106063=>"011010001",
106064=>"000000111",
106065=>"011000010",
106066=>"010111111",
106067=>"100100100",
106068=>"010000000",
106069=>"100011010",
106070=>"101101100",
106071=>"001000110",
106072=>"000000110",
106073=>"001001000",
106074=>"100000000",
106075=>"110100011",
106076=>"000110010",
106077=>"011111101",
106078=>"010010010",
106079=>"011010100",
106080=>"000000000",
106081=>"001000010",
106082=>"000101000",
106083=>"001001000",
106084=>"110111110",
106085=>"111001011",
106086=>"010001100",
106087=>"010000100",
106088=>"111011111",
106089=>"101000101",
106090=>"011011000",
106091=>"110001101",
106092=>"101000011",
106093=>"101111111",
106094=>"000100000",
106095=>"010100000",
106096=>"111001001",
106097=>"111100000",
106098=>"000000110",
106099=>"001101111",
106100=>"001011111",
106101=>"000101111",
106102=>"000001000",
106103=>"000010100",
106104=>"000000001",
106105=>"001101101",
106106=>"011111101",
106107=>"111111000",
106108=>"000100100",
106109=>"000001101",
106110=>"000100001",
106111=>"010010000",
106112=>"000000000",
106113=>"111000000",
106114=>"000001111",
106115=>"111111111",
106116=>"111111011",
106117=>"101000111",
106118=>"100100101",
106119=>"000100000",
106120=>"010000000",
106121=>"110111111",
106122=>"111111000",
106123=>"001000000",
106124=>"010000010",
106125=>"100100000",
106126=>"110001001",
106127=>"001101101",
106128=>"101101101",
106129=>"101001001",
106130=>"111101001",
106131=>"001000000",
106132=>"111111111",
106133=>"000000000",
106134=>"010111111",
106135=>"011011100",
106136=>"011101000",
106137=>"010101111",
106138=>"000011110",
106139=>"000011000",
106140=>"111010010",
106141=>"001000101",
106142=>"111101010",
106143=>"111101000",
106144=>"011111111",
106145=>"011001111",
106146=>"111101101",
106147=>"111000000",
106148=>"100110110",
106149=>"000000001",
106150=>"000001000",
106151=>"011011001",
106152=>"110111011",
106153=>"010000010",
106154=>"101101101",
106155=>"000000000",
106156=>"111110111",
106157=>"010000100",
106158=>"100001111",
106159=>"110111010",
106160=>"111110000",
106161=>"010000011",
106162=>"101111111",
106163=>"110001000",
106164=>"111101001",
106165=>"000111100",
106166=>"000000100",
106167=>"000001001",
106168=>"111111011",
106169=>"011011110",
106170=>"000101001",
106171=>"001110010",
106172=>"000101101",
106173=>"101100000",
106174=>"011110000",
106175=>"100000010",
106176=>"111000000",
106177=>"001101000",
106178=>"110111111",
106179=>"111100001",
106180=>"000000000",
106181=>"001011110",
106182=>"111011000",
106183=>"100000001",
106184=>"011011010",
106185=>"010010011",
106186=>"001000101",
106187=>"000000001",
106188=>"010110111",
106189=>"110000001",
106190=>"000000000",
106191=>"000101001",
106192=>"010010111",
106193=>"100110011",
106194=>"100010000",
106195=>"011111011",
106196=>"000001000",
106197=>"101001110",
106198=>"001000111",
106199=>"100111010",
106200=>"001000000",
106201=>"110010011",
106202=>"110100101",
106203=>"101000000",
106204=>"101101000",
106205=>"010100010",
106206=>"000101100",
106207=>"010110010",
106208=>"010010000",
106209=>"000111000",
106210=>"111101000",
106211=>"110011011",
106212=>"100101001",
106213=>"111001111",
106214=>"110110101",
106215=>"011000110",
106216=>"111111101",
106217=>"110000000",
106218=>"001010111",
106219=>"000001100",
106220=>"000000000",
106221=>"111001000",
106222=>"110100000",
106223=>"111111100",
106224=>"000000101",
106225=>"000100001",
106226=>"000010010",
106227=>"001001000",
106228=>"100001001",
106229=>"101011010",
106230=>"000000000",
106231=>"010000000",
106232=>"001000000",
106233=>"111001111",
106234=>"111100100",
106235=>"100000110",
106236=>"000011001",
106237=>"011100000",
106238=>"110110000",
106239=>"000101111",
106240=>"111101111",
106241=>"100000000",
106242=>"000110010",
106243=>"000000000",
106244=>"001101000",
106245=>"000100111",
106246=>"001010000",
106247=>"111000001",
106248=>"000000000",
106249=>"011111000",
106250=>"000111111",
106251=>"001001001",
106252=>"111001000",
106253=>"100000000",
106254=>"001011110",
106255=>"010000111",
106256=>"000011101",
106257=>"000000110",
106258=>"000000000",
106259=>"110000111",
106260=>"110101101",
106261=>"111001111",
106262=>"111100000",
106263=>"000011000",
106264=>"000010101",
106265=>"001000001",
106266=>"100000101",
106267=>"111111010",
106268=>"100000110",
106269=>"010011010",
106270=>"000100010",
106271=>"000000000",
106272=>"111111111",
106273=>"000000001",
106274=>"011000001",
106275=>"100000001",
106276=>"011110110",
106277=>"100100111",
106278=>"001001000",
106279=>"001111111",
106280=>"111011101",
106281=>"111101000",
106282=>"000000000",
106283=>"001000100",
106284=>"000000000",
106285=>"111000110",
106286=>"011011000",
106287=>"001110000",
106288=>"000000001",
106289=>"011111011",
106290=>"000101101",
106291=>"000111000",
106292=>"000111111",
106293=>"110111111",
106294=>"111111111",
106295=>"000000000",
106296=>"010000101",
106297=>"000000000",
106298=>"000010111",
106299=>"100010001",
106300=>"111100000",
106301=>"000011011",
106302=>"110010010",
106303=>"000000000",
106304=>"111111110",
106305=>"000000011",
106306=>"000100000",
106307=>"000001111",
106308=>"000000001",
106309=>"101101101",
106310=>"110000110",
106311=>"110111110",
106312=>"000000000",
106313=>"011010000",
106314=>"000000000",
106315=>"000000111",
106316=>"100110111",
106317=>"100110011",
106318=>"100111111",
106319=>"000111111",
106320=>"000000000",
106321=>"001010011",
106322=>"000000110",
106323=>"011011111",
106324=>"111111111",
106325=>"000000000",
106326=>"100100111",
106327=>"111111000",
106328=>"000000000",
106329=>"010001001",
106330=>"000000000",
106331=>"011000100",
106332=>"001000000",
106333=>"010010000",
106334=>"001111011",
106335=>"110111111",
106336=>"110000100",
106337=>"010000000",
106338=>"111011000",
106339=>"001000000",
106340=>"000000000",
106341=>"000011111",
106342=>"011111111",
106343=>"010010010",
106344=>"000000000",
106345=>"111100111",
106346=>"111000000",
106347=>"100000000",
106348=>"111111011",
106349=>"001011111",
106350=>"111000000",
106351=>"111000101",
106352=>"111110011",
106353=>"000000111",
106354=>"111111111",
106355=>"111111111",
106356=>"101101111",
106357=>"100100111",
106358=>"111101000",
106359=>"111111111",
106360=>"010111110",
106361=>"000000001",
106362=>"000001111",
106363=>"101111000",
106364=>"111111110",
106365=>"101111110",
106366=>"111000000",
106367=>"000111000",
106368=>"111000111",
106369=>"000000000",
106370=>"000000000",
106371=>"000000000",
106372=>"111111100",
106373=>"100011111",
106374=>"011000010",
106375=>"110100000",
106376=>"000101000",
106377=>"000100000",
106378=>"111111111",
106379=>"101000111",
106380=>"000000111",
106381=>"000000000",
106382=>"111111100",
106383=>"100000101",
106384=>"111001010",
106385=>"001000000",
106386=>"000000000",
106387=>"000000111",
106388=>"000100100",
106389=>"111000000",
106390=>"000000000",
106391=>"111110010",
106392=>"111111101",
106393=>"000111001",
106394=>"000011001",
106395=>"111111000",
106396=>"101000111",
106397=>"001000000",
106398=>"000101101",
106399=>"000010001",
106400=>"101100000",
106401=>"111111101",
106402=>"001000000",
106403=>"000000000",
106404=>"000000010",
106405=>"110000001",
106406=>"001000001",
106407=>"000000000",
106408=>"000000000",
106409=>"000101100",
106410=>"000000000",
106411=>"110100111",
106412=>"101101111",
106413=>"100110000",
106414=>"011111110",
106415=>"111111111",
106416=>"000000000",
106417=>"000000010",
106418=>"111011000",
106419=>"111110100",
106420=>"011110100",
106421=>"000010111",
106422=>"010010000",
106423=>"101101010",
106424=>"011001000",
106425=>"111001011",
106426=>"111110101",
106427=>"000000000",
106428=>"100000011",
106429=>"000111011",
106430=>"000000000",
106431=>"000000100",
106432=>"010001111",
106433=>"000000111",
106434=>"101001000",
106435=>"100111000",
106436=>"000111111",
106437=>"100001000",
106438=>"011111000",
106439=>"011010000",
106440=>"000101101",
106441=>"111111111",
106442=>"110101111",
106443=>"000000100",
106444=>"111111111",
106445=>"110111000",
106446=>"000000000",
106447=>"111110000",
106448=>"111111000",
106449=>"111011000",
106450=>"100101111",
106451=>"011011010",
106452=>"000000001",
106453=>"111011011",
106454=>"111111010",
106455=>"000111011",
106456=>"000000000",
106457=>"000111101",
106458=>"001001000",
106459=>"010111111",
106460=>"110100000",
106461=>"011111111",
106462=>"111111111",
106463=>"001000001",
106464=>"000011010",
106465=>"111111111",
106466=>"111111111",
106467=>"111110111",
106468=>"010010010",
106469=>"110100000",
106470=>"001111110",
106471=>"100100001",
106472=>"111101111",
106473=>"111000000",
106474=>"111111111",
106475=>"111111111",
106476=>"000000000",
106477=>"101111111",
106478=>"111000000",
106479=>"110101111",
106480=>"001111011",
106481=>"001000000",
106482=>"000000100",
106483=>"001000011",
106484=>"111101001",
106485=>"000111111",
106486=>"011011111",
106487=>"000000000",
106488=>"000000000",
106489=>"111001000",
106490=>"011110101",
106491=>"111100010",
106492=>"000001000",
106493=>"011100101",
106494=>"001111110",
106495=>"111111110",
106496=>"011001001",
106497=>"000000111",
106498=>"110011111",
106499=>"000001001",
106500=>"100000000",
106501=>"000000000",
106502=>"000001010",
106503=>"010000011",
106504=>"100000000",
106505=>"101101101",
106506=>"010101001",
106507=>"000000110",
106508=>"010010000",
106509=>"110101100",
106510=>"000011011",
106511=>"111111000",
106512=>"100011111",
106513=>"001001000",
106514=>"010011110",
106515=>"000101111",
106516=>"000001110",
106517=>"011000000",
106518=>"111101101",
106519=>"111000000",
106520=>"111011000",
106521=>"110101010",
106522=>"111000001",
106523=>"111000100",
106524=>"000001010",
106525=>"000000000",
106526=>"111000000",
106527=>"001101000",
106528=>"110111110",
106529=>"111111000",
106530=>"000010000",
106531=>"000000000",
106532=>"110011001",
106533=>"001011111",
106534=>"010001101",
106535=>"111110001",
106536=>"110101010",
106537=>"010110001",
106538=>"101110010",
106539=>"000000011",
106540=>"001011111",
106541=>"000000110",
106542=>"101001001",
106543=>"001001010",
106544=>"000000011",
106545=>"111111100",
106546=>"000000110",
106547=>"101000000",
106548=>"001111111",
106549=>"101111111",
106550=>"111000000",
106551=>"111111001",
106552=>"101000010",
106553=>"001001111",
106554=>"000001000",
106555=>"110000110",
106556=>"011111001",
106557=>"001101001",
106558=>"111111101",
106559=>"001011011",
106560=>"011011111",
106561=>"000111111",
106562=>"100110111",
106563=>"000101111",
106564=>"010010001",
106565=>"111111000",
106566=>"001010111",
106567=>"111011110",
106568=>"000000010",
106569=>"000011110",
106570=>"011011000",
106571=>"011001000",
106572=>"001111111",
106573=>"011101110",
106574=>"011111100",
106575=>"101111111",
106576=>"101000000",
106577=>"001000000",
106578=>"001111111",
106579=>"011000100",
106580=>"000001011",
106581=>"111001100",
106582=>"000011011",
106583=>"001000111",
106584=>"100000001",
106585=>"110110110",
106586=>"000110100",
106587=>"111111111",
106588=>"111100000",
106589=>"001001001",
106590=>"110111011",
106591=>"001000100",
106592=>"111111111",
106593=>"110000100",
106594=>"110111110",
106595=>"011111111",
106596=>"100101100",
106597=>"000100100",
106598=>"000111110",
106599=>"111101001",
106600=>"000101000",
106601=>"110000000",
106602=>"011000111",
106603=>"000000001",
106604=>"010001000",
106605=>"000000011",
106606=>"000000100",
106607=>"001001000",
106608=>"100111101",
106609=>"111101000",
106610=>"110100110",
106611=>"000001111",
106612=>"100111110",
106613=>"000000000",
106614=>"011111111",
106615=>"111111010",
106616=>"100000110",
106617=>"111111111",
106618=>"010111111",
106619=>"000000000",
106620=>"011001010",
106621=>"100000000",
106622=>"000000010",
106623=>"000000000",
106624=>"111110010",
106625=>"100010010",
106626=>"100111000",
106627=>"001111010",
106628=>"000000010",
106629=>"001111001",
106630=>"000100111",
106631=>"110100111",
106632=>"011111100",
106633=>"000001001",
106634=>"110010110",
106635=>"010011001",
106636=>"111101100",
106637=>"000010111",
106638=>"000010010",
106639=>"010001010",
106640=>"111101111",
106641=>"000000111",
106642=>"100001000",
106643=>"010001000",
106644=>"111000000",
106645=>"101000101",
106646=>"110111100",
106647=>"001011001",
106648=>"111101110",
106649=>"000110111",
106650=>"001000001",
106651=>"000110000",
106652=>"101000100",
106653=>"001000000",
106654=>"100000000",
106655=>"000001000",
106656=>"100111000",
106657=>"101010000",
106658=>"101111111",
106659=>"110010110",
106660=>"111001100",
106661=>"011111111",
106662=>"100110110",
106663=>"011111111",
106664=>"111000000",
106665=>"000101111",
106666=>"001110110",
106667=>"000000101",
106668=>"100101011",
106669=>"101000101",
106670=>"010001011",
106671=>"110110111",
106672=>"000000000",
106673=>"011011111",
106674=>"111101101",
106675=>"000001100",
106676=>"110100111",
106677=>"111111111",
106678=>"000111100",
106679=>"000010110",
106680=>"100101101",
106681=>"111001000",
106682=>"111111000",
106683=>"110101111",
106684=>"000110010",
106685=>"000010111",
106686=>"100100000",
106687=>"100000000",
106688=>"000000000",
106689=>"110000110",
106690=>"000101111",
106691=>"110100100",
106692=>"010111010",
106693=>"111111100",
106694=>"101000011",
106695=>"010010000",
106696=>"000111110",
106697=>"001101000",
106698=>"111111101",
106699=>"111111000",
106700=>"011101111",
106701=>"100100111",
106702=>"111010111",
106703=>"111011110",
106704=>"000001101",
106705=>"010111011",
106706=>"011111000",
106707=>"000100000",
106708=>"010111011",
106709=>"100000100",
106710=>"000000110",
106711=>"111000001",
106712=>"000000111",
106713=>"111000000",
106714=>"111111100",
106715=>"000000000",
106716=>"111001011",
106717=>"001001000",
106718=>"000101001",
106719=>"111011001",
106720=>"110011101",
106721=>"000000000",
106722=>"000000001",
106723=>"000010110",
106724=>"010100111",
106725=>"000000000",
106726=>"001011101",
106727=>"111001011",
106728=>"111111000",
106729=>"010010011",
106730=>"000100000",
106731=>"101111110",
106732=>"001000110",
106733=>"000000000",
106734=>"000000000",
106735=>"000110000",
106736=>"000000100",
106737=>"110000000",
106738=>"111101000",
106739=>"001000001",
106740=>"111100100",
106741=>"001000001",
106742=>"000010111",
106743=>"010111101",
106744=>"110010101",
106745=>"000000101",
106746=>"100000000",
106747=>"111011000",
106748=>"111010000",
106749=>"000000011",
106750=>"100000011",
106751=>"110110111",
106752=>"001000010",
106753=>"111111111",
106754=>"001011001",
106755=>"100110110",
106756=>"001011111",
106757=>"001011010",
106758=>"110111100",
106759=>"000011010",
106760=>"001001001",
106761=>"011011001",
106762=>"000101001",
106763=>"011011010",
106764=>"011001001",
106765=>"110111010",
106766=>"111000000",
106767=>"000011000",
106768=>"000000010",
106769=>"110011111",
106770=>"100001110",
106771=>"010000100",
106772=>"100010100",
106773=>"100110000",
106774=>"010011011",
106775=>"000001011",
106776=>"000000000",
106777=>"000000100",
106778=>"110010110",
106779=>"011001011",
106780=>"000000100",
106781=>"100100000",
106782=>"010010011",
106783=>"000000110",
106784=>"011011001",
106785=>"000011011",
106786=>"001111111",
106787=>"000001011",
106788=>"011011010",
106789=>"000010110",
106790=>"011110000",
106791=>"010010011",
106792=>"001111011",
106793=>"000100110",
106794=>"011010011",
106795=>"100001011",
106796=>"101100000",
106797=>"100110111",
106798=>"110011111",
106799=>"000100010",
106800=>"000001000",
106801=>"000111001",
106802=>"011010100",
106803=>"000100100",
106804=>"000001000",
106805=>"100100000",
106806=>"101100000",
106807=>"110001011",
106808=>"000010011",
106809=>"011000110",
106810=>"100100110",
106811=>"001000001",
106812=>"001001011",
106813=>"000110111",
106814=>"011011011",
106815=>"110010001",
106816=>"011001001",
106817=>"000011110",
106818=>"111101110",
106819=>"011011011",
106820=>"001100110",
106821=>"000000010",
106822=>"011000000",
106823=>"101101000",
106824=>"111110101",
106825=>"110000011",
106826=>"010010011",
106827=>"100110000",
106828=>"111011001",
106829=>"000011011",
106830=>"011000000",
106831=>"011011110",
106832=>"011010000",
106833=>"100111111",
106834=>"111111100",
106835=>"100111011",
106836=>"011010110",
106837=>"000001001",
106838=>"001011101",
106839=>"010001011",
106840=>"001111101",
106841=>"100110100",
106842=>"100111111",
106843=>"111111001",
106844=>"001001000",
106845=>"001101101",
106846=>"111110010",
106847=>"011011011",
106848=>"010011011",
106849=>"010000000",
106850=>"011001001",
106851=>"100100010",
106852=>"011001011",
106853=>"111100101",
106854=>"011100000",
106855=>"100100100",
106856=>"000101000",
106857=>"001110100",
106858=>"110010111",
106859=>"011110011",
106860=>"000010000",
106861=>"100100100",
106862=>"010001011",
106863=>"110011010",
106864=>"011110011",
106865=>"000001011",
106866=>"000010010",
106867=>"000100000",
106868=>"101111111",
106869=>"010010010",
106870=>"011110110",
106871=>"110000000",
106872=>"000010011",
106873=>"100100101",
106874=>"110011110",
106875=>"100101001",
106876=>"111011011",
106877=>"101000000",
106878=>"011100001",
106879=>"111001000",
106880=>"010011011",
106881=>"000000001",
106882=>"100001011",
106883=>"100100000",
106884=>"101101100",
106885=>"110000000",
106886=>"000000111",
106887=>"111010000",
106888=>"001111010",
106889=>"000100000",
106890=>"101100101",
106891=>"101001000",
106892=>"000000000",
106893=>"011011011",
106894=>"110001111",
106895=>"001001000",
106896=>"101111110",
106897=>"011011001",
106898=>"111011010",
106899=>"011011011",
106900=>"101001001",
106901=>"011001011",
106902=>"100110100",
106903=>"001001001",
106904=>"010010010",
106905=>"001100100",
106906=>"011001001",
106907=>"111111011",
106908=>"111000111",
106909=>"011011011",
106910=>"101011000",
106911=>"011010010",
106912=>"111011010",
106913=>"100100110",
106914=>"111000000",
106915=>"000100100",
106916=>"100110100",
106917=>"010000000",
106918=>"001000111",
106919=>"001011100",
106920=>"100100111",
106921=>"011011111",
106922=>"001011011",
106923=>"011001001",
106924=>"000000111",
106925=>"000001000",
106926=>"011000010",
106927=>"100111110",
106928=>"011001001",
106929=>"000010110",
106930=>"100011111",
106931=>"000001001",
106932=>"100101101",
106933=>"100100101",
106934=>"100010111",
106935=>"011011011",
106936=>"010000000",
106937=>"000000001",
106938=>"101100110",
106939=>"111011000",
106940=>"100110100",
106941=>"001001111",
106942=>"000000001",
106943=>"000100110",
106944=>"101001011",
106945=>"100110001",
106946=>"111011000",
106947=>"000110001",
106948=>"000100111",
106949=>"110011110",
106950=>"101001001",
106951=>"100000001",
106952=>"100010010",
106953=>"001000010",
106954=>"110110111",
106955=>"000000100",
106956=>"011011000",
106957=>"011010001",
106958=>"100100100",
106959=>"010011001",
106960=>"111110100",
106961=>"111110111",
106962=>"000111110",
106963=>"111100001",
106964=>"011011011",
106965=>"000000000",
106966=>"011001011",
106967=>"111110001",
106968=>"000010110",
106969=>"110110100",
106970=>"001001001",
106971=>"100100100",
106972=>"111111011",
106973=>"010100111",
106974=>"001110110",
106975=>"110010000",
106976=>"111111110",
106977=>"111100111",
106978=>"101100000",
106979=>"011011011",
106980=>"010010000",
106981=>"000110110",
106982=>"111001001",
106983=>"011111011",
106984=>"011111000",
106985=>"000000000",
106986=>"110110000",
106987=>"001000011",
106988=>"010011011",
106989=>"100110110",
106990=>"000001100",
106991=>"000001011",
106992=>"000000000",
106993=>"000001111",
106994=>"011001001",
106995=>"000000000",
106996=>"001011011",
106997=>"000100100",
106998=>"000000000",
106999=>"010100001",
107000=>"011011011",
107001=>"100000000",
107002=>"111111111",
107003=>"111100100",
107004=>"001001001",
107005=>"000000000",
107006=>"111000000",
107007=>"111010011",
107008=>"001001011",
107009=>"111111111",
107010=>"111101111",
107011=>"101101000",
107012=>"111111111",
107013=>"111001110",
107014=>"011111001",
107015=>"001010111",
107016=>"010111111",
107017=>"001000011",
107018=>"001100100",
107019=>"000111001",
107020=>"011010000",
107021=>"010111010",
107022=>"100110110",
107023=>"110000010",
107024=>"000001011",
107025=>"010100111",
107026=>"111101101",
107027=>"001001000",
107028=>"111111111",
107029=>"101000101",
107030=>"101100111",
107031=>"110100100",
107032=>"101101110",
107033=>"001111000",
107034=>"000011010",
107035=>"000111101",
107036=>"000000110",
107037=>"111000000",
107038=>"100101101",
107039=>"000111010",
107040=>"001101111",
107041=>"111111010",
107042=>"000100001",
107043=>"111111010",
107044=>"101011110",
107045=>"100100110",
107046=>"100100011",
107047=>"000000100",
107048=>"100111110",
107049=>"011011111",
107050=>"001001000",
107051=>"000000000",
107052=>"010011001",
107053=>"110111001",
107054=>"111101010",
107055=>"101101110",
107056=>"100001111",
107057=>"000111111",
107058=>"001000010",
107059=>"100000001",
107060=>"101000000",
107061=>"000111111",
107062=>"000000100",
107063=>"000000000",
107064=>"101101111",
107065=>"000000010",
107066=>"011010111",
107067=>"000000101",
107068=>"010111110",
107069=>"010111000",
107070=>"000000000",
107071=>"110101111",
107072=>"000100000",
107073=>"000000110",
107074=>"101101111",
107075=>"001000010",
107076=>"110000110",
107077=>"001000000",
107078=>"110010000",
107079=>"000101000",
107080=>"111111000",
107081=>"101111111",
107082=>"100000101",
107083=>"101001110",
107084=>"000000110",
107085=>"000111111",
107086=>"001111111",
107087=>"000011111",
107088=>"000000111",
107089=>"110000100",
107090=>"001101000",
107091=>"011000000",
107092=>"101101100",
107093=>"011011011",
107094=>"111111111",
107095=>"000000000",
107096=>"010110100",
107097=>"000010100",
107098=>"100100111",
107099=>"001010111",
107100=>"001001111",
107101=>"000010010",
107102=>"110011101",
107103=>"100010111",
107104=>"000010010",
107105=>"000111111",
107106=>"100000111",
107107=>"001011110",
107108=>"000111111",
107109=>"011100000",
107110=>"110111000",
107111=>"110000011",
107112=>"011110000",
107113=>"110000100",
107114=>"010000000",
107115=>"111110000",
107116=>"110110000",
107117=>"100100100",
107118=>"011000110",
107119=>"000000000",
107120=>"000111111",
107121=>"100101100",
107122=>"000001001",
107123=>"001000001",
107124=>"000000000",
107125=>"111000000",
107126=>"000000000",
107127=>"000000101",
107128=>"101001000",
107129=>"110111100",
107130=>"011000001",
107131=>"001000000",
107132=>"000011011",
107133=>"111100010",
107134=>"111001110",
107135=>"101000011",
107136=>"110000000",
107137=>"111101000",
107138=>"010010011",
107139=>"111111000",
107140=>"001111000",
107141=>"111000000",
107142=>"010001011",
107143=>"000110110",
107144=>"000110110",
107145=>"100001101",
107146=>"111100100",
107147=>"010010000",
107148=>"110011001",
107149=>"000010010",
107150=>"111110101",
107151=>"001001001",
107152=>"110110110",
107153=>"111111010",
107154=>"101100110",
107155=>"100101001",
107156=>"001101011",
107157=>"101000101",
107158=>"000000001",
107159=>"010111011",
107160=>"000111101",
107161=>"101000100",
107162=>"000111110",
107163=>"000000010",
107164=>"010010010",
107165=>"101101110",
107166=>"110000100",
107167=>"111101000",
107168=>"011101100",
107169=>"100000001",
107170=>"111010000",
107171=>"101101000",
107172=>"000111100",
107173=>"110000000",
107174=>"110000111",
107175=>"000010010",
107176=>"010010101",
107177=>"000001001",
107178=>"011011111",
107179=>"101000010",
107180=>"111110000",
107181=>"000000110",
107182=>"000100110",
107183=>"000010000",
107184=>"010101101",
107185=>"011011100",
107186=>"000111111",
107187=>"000001011",
107188=>"011011010",
107189=>"111100110",
107190=>"011011000",
107191=>"111101010",
107192=>"110111011",
107193=>"000110011",
107194=>"111000111",
107195=>"000111010",
107196=>"000110000",
107197=>"010111111",
107198=>"011001010",
107199=>"000101111",
107200=>"000001000",
107201=>"000100000",
107202=>"011000010",
107203=>"100101011",
107204=>"000000000",
107205=>"000000000",
107206=>"111011111",
107207=>"001000010",
107208=>"000000111",
107209=>"001000000",
107210=>"111000000",
107211=>"010110111",
107212=>"000101111",
107213=>"000110110",
107214=>"001000000",
107215=>"010111000",
107216=>"111111011",
107217=>"110010110",
107218=>"000000000",
107219=>"011000000",
107220=>"001110110",
107221=>"111110000",
107222=>"101100111",
107223=>"010000000",
107224=>"111000001",
107225=>"011010010",
107226=>"110100001",
107227=>"101000111",
107228=>"101001110",
107229=>"010000000",
107230=>"111001000",
107231=>"001100110",
107232=>"001111111",
107233=>"101101000",
107234=>"100001101",
107235=>"011011011",
107236=>"101101101",
107237=>"110110000",
107238=>"011010000",
107239=>"000000110",
107240=>"111000001",
107241=>"000000101",
107242=>"100000000",
107243=>"000000011",
107244=>"010010001",
107245=>"001000101",
107246=>"110001000",
107247=>"111000000",
107248=>"000000100",
107249=>"000000011",
107250=>"010101001",
107251=>"110110110",
107252=>"110110110",
107253=>"101000101",
107254=>"000000000",
107255=>"000001111",
107256=>"101000101",
107257=>"010000000",
107258=>"111111111",
107259=>"000000000",
107260=>"010010111",
107261=>"100010001",
107262=>"011010110",
107263=>"000101000",
107264=>"000000110",
107265=>"000100010",
107266=>"000101110",
107267=>"000000000",
107268=>"011001111",
107269=>"101101001",
107270=>"110110110",
107271=>"111110000",
107272=>"000000111",
107273=>"111000000",
107274=>"000000110",
107275=>"000000000",
107276=>"000000111",
107277=>"101111001",
107278=>"000000110",
107279=>"001000111",
107280=>"111111000",
107281=>"111111000",
107282=>"000111011",
107283=>"100111110",
107284=>"000110110",
107285=>"110111111",
107286=>"011110111",
107287=>"110111000",
107288=>"110000000",
107289=>"010111000",
107290=>"111111111",
107291=>"110010100",
107292=>"111101111",
107293=>"000110110",
107294=>"111111110",
107295=>"000001101",
107296=>"000101110",
107297=>"000100000",
107298=>"011000000",
107299=>"000100110",
107300=>"000010100",
107301=>"101011110",
107302=>"000000111",
107303=>"000111110",
107304=>"011110000",
107305=>"011000110",
107306=>"101101101",
107307=>"110010000",
107308=>"000001111",
107309=>"101110111",
107310=>"101111110",
107311=>"010110001",
107312=>"001001100",
107313=>"000101111",
107314=>"111000010",
107315=>"111000000",
107316=>"000010111",
107317=>"010000000",
107318=>"000100100",
107319=>"000000000",
107320=>"111111011",
107321=>"000001111",
107322=>"111001000",
107323=>"111111011",
107324=>"000111111",
107325=>"111001000",
107326=>"001001111",
107327=>"001110101",
107328=>"111010110",
107329=>"101001000",
107330=>"101000000",
107331=>"100111011",
107332=>"000101110",
107333=>"000001111",
107334=>"111000101",
107335=>"001001000",
107336=>"000110110",
107337=>"111111000",
107338=>"001000111",
107339=>"001101100",
107340=>"110111111",
107341=>"011001011",
107342=>"100010110",
107343=>"000000110",
107344=>"001111111",
107345=>"111111000",
107346=>"000001110",
107347=>"000011011",
107348=>"000000000",
107349=>"111111111",
107350=>"000010111",
107351=>"111110000",
107352=>"100111110",
107353=>"110111111",
107354=>"000100101",
107355=>"100110111",
107356=>"001111110",
107357=>"001101101",
107358=>"111111111",
107359=>"011111101",
107360=>"000110111",
107361=>"000000000",
107362=>"000000011",
107363=>"011011111",
107364=>"000001001",
107365=>"111111000",
107366=>"000110000",
107367=>"001000000",
107368=>"111111000",
107369=>"111111000",
107370=>"000000011",
107371=>"001001110",
107372=>"000111110",
107373=>"111000000",
107374=>"000100100",
107375=>"000000000",
107376=>"000011011",
107377=>"111000000",
107378=>"100010011",
107379=>"001001111",
107380=>"100100111",
107381=>"000001111",
107382=>"111000000",
107383=>"000000111",
107384=>"111101111",
107385=>"010001111",
107386=>"000000110",
107387=>"000100111",
107388=>"001011011",
107389=>"000000100",
107390=>"101111111",
107391=>"000001111",
107392=>"001010110",
107393=>"000010000",
107394=>"011110111",
107395=>"111000000",
107396=>"000000000",
107397=>"100001000",
107398=>"100011110",
107399=>"000000000",
107400=>"000010000",
107401=>"000000000",
107402=>"000000001",
107403=>"001000100",
107404=>"110111000",
107405=>"111111000",
107406=>"111100101",
107407=>"000001010",
107408=>"000000011",
107409=>"000000110",
107410=>"111111001",
107411=>"111010000",
107412=>"000000000",
107413=>"111111000",
107414=>"111111111",
107415=>"000101101",
107416=>"000110111",
107417=>"011111000",
107418=>"000000010",
107419=>"111000100",
107420=>"000001001",
107421=>"010111001",
107422=>"001110111",
107423=>"000000100",
107424=>"001111110",
107425=>"111110110",
107426=>"000001000",
107427=>"110101000",
107428=>"111111110",
107429=>"001011111",
107430=>"101001111",
107431=>"001111111",
107432=>"111111110",
107433=>"110111111",
107434=>"111000011",
107435=>"000000011",
107436=>"111100001",
107437=>"000000010",
107438=>"000101100",
107439=>"001101111",
107440=>"000111111",
107441=>"011001000",
107442=>"010001111",
107443=>"010001010",
107444=>"000111100",
107445=>"111111111",
107446=>"000000101",
107447=>"000001010",
107448=>"000111111",
107449=>"001001010",
107450=>"000001111",
107451=>"000001111",
107452=>"111001111",
107453=>"111110001",
107454=>"110011011",
107455=>"111110110",
107456=>"000111000",
107457=>"000000100",
107458=>"111111111",
107459=>"000001111",
107460=>"000001111",
107461=>"000010111",
107462=>"000110001",
107463=>"101101110",
107464=>"010000001",
107465=>"010101111",
107466=>"111111100",
107467=>"000000110",
107468=>"000111011",
107469=>"001111100",
107470=>"110110111",
107471=>"111110111",
107472=>"111010011",
107473=>"000011111",
107474=>"011000010",
107475=>"101111101",
107476=>"000111111",
107477=>"000001010",
107478=>"000011111",
107479=>"111101100",
107480=>"000100111",
107481=>"000000111",
107482=>"001101101",
107483=>"111000000",
107484=>"110111111",
107485=>"000001000",
107486=>"000101111",
107487=>"111101111",
107488=>"111000001",
107489=>"000000000",
107490=>"111101011",
107491=>"001011111",
107492=>"001001110",
107493=>"110111011",
107494=>"111001111",
107495=>"011111111",
107496=>"111111111",
107497=>"000000100",
107498=>"000000001",
107499=>"001000000",
107500=>"000111111",
107501=>"011101000",
107502=>"111000000",
107503=>"000000110",
107504=>"000000101",
107505=>"001111111",
107506=>"000001110",
107507=>"110111110",
107508=>"000001011",
107509=>"001000100",
107510=>"100000111",
107511=>"111000010",
107512=>"111111000",
107513=>"111111111",
107514=>"111000010",
107515=>"000110111",
107516=>"000010111",
107517=>"000111000",
107518=>"000000011",
107519=>"000000110",
107520=>"011000101",
107521=>"000000100",
107522=>"111101100",
107523=>"000000010",
107524=>"001001111",
107525=>"110101111",
107526=>"110111101",
107527=>"000011010",
107528=>"000110111",
107529=>"110000000",
107530=>"001011100",
107531=>"111001000",
107532=>"001010011",
107533=>"000010011",
107534=>"000000010",
107535=>"111111011",
107536=>"000110010",
107537=>"000000101",
107538=>"000000000",
107539=>"111111101",
107540=>"111110101",
107541=>"111101001",
107542=>"100111111",
107543=>"010010111",
107544=>"100000111",
107545=>"000100110",
107546=>"000000000",
107547=>"000001010",
107548=>"100100111",
107549=>"101000101",
107550=>"010100101",
107551=>"000100101",
107552=>"000000100",
107553=>"010110010",
107554=>"000000000",
107555=>"000111010",
107556=>"000100110",
107557=>"111011011",
107558=>"000011000",
107559=>"000010000",
107560=>"111111000",
107561=>"010010111",
107562=>"011001000",
107563=>"101101011",
107564=>"000011011",
107565=>"010010101",
107566=>"010111111",
107567=>"000110010",
107568=>"101100110",
107569=>"001111110",
107570=>"000000010",
107571=>"000100100",
107572=>"000001000",
107573=>"110110000",
107574=>"100101001",
107575=>"001000000",
107576=>"010111111",
107577=>"000001000",
107578=>"011000100",
107579=>"101101000",
107580=>"000001101",
107581=>"000111110",
107582=>"101101111",
107583=>"011110100",
107584=>"101001001",
107585=>"010000111",
107586=>"111101001",
107587=>"001001100",
107588=>"110110110",
107589=>"001000000",
107590=>"000101111",
107591=>"000010110",
107592=>"000011110",
107593=>"111110010",
107594=>"111111011",
107595=>"011000100",
107596=>"000000000",
107597=>"001101111",
107598=>"110111111",
107599=>"111111111",
107600=>"000000000",
107601=>"110011110",
107602=>"010010000",
107603=>"010011001",
107604=>"000101101",
107605=>"000001011",
107606=>"001111100",
107607=>"101000100",
107608=>"110100000",
107609=>"000011111",
107610=>"100101110",
107611=>"000000011",
107612=>"111101101",
107613=>"100001011",
107614=>"111111111",
107615=>"100001001",
107616=>"000110011",
107617=>"001101101",
107618=>"010101111",
107619=>"000110100",
107620=>"000110111",
107621=>"011011001",
107622=>"000110100",
107623=>"111000000",
107624=>"011100100",
107625=>"010000110",
107626=>"010000000",
107627=>"010110000",
107628=>"000011010",
107629=>"100110100",
107630=>"000001100",
107631=>"000101000",
107632=>"101111111",
107633=>"010010001",
107634=>"001100100",
107635=>"000000000",
107636=>"111111111",
107637=>"001000000",
107638=>"000110111",
107639=>"011000110",
107640=>"111001111",
107641=>"000010100",
107642=>"000000101",
107643=>"111000000",
107644=>"001011011",
107645=>"010100000",
107646=>"000101011",
107647=>"001000100",
107648=>"010010000",
107649=>"111100000",
107650=>"010010010",
107651=>"000010000",
107652=>"111111000",
107653=>"000001110",
107654=>"111100000",
107655=>"100110110",
107656=>"111111010",
107657=>"011000000",
107658=>"011010111",
107659=>"010010000",
107660=>"111000100",
107661=>"101001000",
107662=>"111000100",
107663=>"011001000",
107664=>"100110110",
107665=>"001101101",
107666=>"000000010",
107667=>"111111111",
107668=>"101010110",
107669=>"010000000",
107670=>"111111100",
107671=>"000111010",
107672=>"100010010",
107673=>"101000110",
107674=>"011101100",
107675=>"101101010",
107676=>"000000000",
107677=>"100000100",
107678=>"111010110",
107679=>"111101000",
107680=>"101101111",
107681=>"101100100",
107682=>"000110000",
107683=>"010000000",
107684=>"010100011",
107685=>"010110000",
107686=>"000000001",
107687=>"000010010",
107688=>"010010110",
107689=>"011010110",
107690=>"111111111",
107691=>"101101000",
107692=>"000010001",
107693=>"000000110",
107694=>"100101011",
107695=>"010010010",
107696=>"000100000",
107697=>"101011011",
107698=>"001011000",
107699=>"000001110",
107700=>"000010011",
107701=>"010000101",
107702=>"011011000",
107703=>"011001000",
107704=>"000110110",
107705=>"011000011",
107706=>"011111111",
107707=>"001000000",
107708=>"011111010",
107709=>"111110011",
107710=>"000011001",
107711=>"000000001",
107712=>"000000000",
107713=>"101101100",
107714=>"111010010",
107715=>"001011001",
107716=>"000000000",
107717=>"100100100",
107718=>"000010010",
107719=>"000001000",
107720=>"111100010",
107721=>"101111111",
107722=>"111110000",
107723=>"110101101",
107724=>"000000100",
107725=>"100110010",
107726=>"101000000",
107727=>"000000101",
107728=>"111000000",
107729=>"100110111",
107730=>"011011000",
107731=>"100111000",
107732=>"000001000",
107733=>"000000100",
107734=>"111010010",
107735=>"010111000",
107736=>"000000111",
107737=>"000001011",
107738=>"101110100",
107739=>"111000000",
107740=>"001001110",
107741=>"111100101",
107742=>"110010010",
107743=>"110000010",
107744=>"111000000",
107745=>"111000100",
107746=>"111000010",
107747=>"000111111",
107748=>"101101111",
107749=>"100011000",
107750=>"111111010",
107751=>"011111101",
107752=>"101101000",
107753=>"000000101",
107754=>"100101001",
107755=>"111001001",
107756=>"001000000",
107757=>"111011000",
107758=>"001000000",
107759=>"000000111",
107760=>"110110000",
107761=>"011001001",
107762=>"000101111",
107763=>"010110110",
107764=>"000110111",
107765=>"111101101",
107766=>"010000100",
107767=>"111110111",
107768=>"010000000",
107769=>"110010010",
107770=>"011011000",
107771=>"101101011",
107772=>"101111011",
107773=>"110111100",
107774=>"100111111",
107775=>"010100000",
107776=>"100100100",
107777=>"010010101",
107778=>"010111111",
107779=>"111111111",
107780=>"011011011",
107781=>"111111010",
107782=>"000010000",
107783=>"100000111",
107784=>"111111011",
107785=>"101100111",
107786=>"001001000",
107787=>"000100000",
107788=>"010111011",
107789=>"000000000",
107790=>"111100101",
107791=>"000000001",
107792=>"011111111",
107793=>"001000000",
107794=>"101011010",
107795=>"111000100",
107796=>"000010010",
107797=>"111111111",
107798=>"000100010",
107799=>"101000100",
107800=>"010000111",
107801=>"010101000",
107802=>"010000000",
107803=>"101000100",
107804=>"101111011",
107805=>"100001101",
107806=>"001101000",
107807=>"110100101",
107808=>"010111110",
107809=>"010010010",
107810=>"111100101",
107811=>"001000000",
107812=>"000011011",
107813=>"011001000",
107814=>"000011010",
107815=>"110100100",
107816=>"010111111",
107817=>"101001101",
107818=>"101100100",
107819=>"000000000",
107820=>"111011111",
107821=>"101000001",
107822=>"000000000",
107823=>"000000000",
107824=>"000111111",
107825=>"011110000",
107826=>"100000100",
107827=>"000011001",
107828=>"000000000",
107829=>"000000011",
107830=>"100000001",
107831=>"000101100",
107832=>"110110100",
107833=>"100101111",
107834=>"111111011",
107835=>"000100110",
107836=>"001011011",
107837=>"000111111",
107838=>"000000010",
107839=>"000000100",
107840=>"111000110",
107841=>"100000000",
107842=>"100111000",
107843=>"011110000",
107844=>"110111111",
107845=>"000000111",
107846=>"111001111",
107847=>"111101111",
107848=>"101011010",
107849=>"011010010",
107850=>"111100101",
107851=>"001000000",
107852=>"111011101",
107853=>"000100000",
107854=>"100111111",
107855=>"000111101",
107856=>"100000111",
107857=>"110111111",
107858=>"110111010",
107859=>"010111101",
107860=>"111000000",
107861=>"111011010",
107862=>"000001001",
107863=>"111101001",
107864=>"000001011",
107865=>"000110100",
107866=>"011011011",
107867=>"000111000",
107868=>"000111010",
107869=>"010110000",
107870=>"111111010",
107871=>"011110110",
107872=>"000100100",
107873=>"000101001",
107874=>"001000000",
107875=>"111111111",
107876=>"000011010",
107877=>"111111100",
107878=>"010000010",
107879=>"100101100",
107880=>"011001000",
107881=>"000000000",
107882=>"011000000",
107883=>"111111111",
107884=>"000000010",
107885=>"000011100",
107886=>"000000000",
107887=>"111011010",
107888=>"100110110",
107889=>"001000000",
107890=>"000000100",
107891=>"100100000",
107892=>"101111000",
107893=>"101000011",
107894=>"110011000",
107895=>"110100000",
107896=>"111001000",
107897=>"011011001",
107898=>"000000000",
107899=>"111111000",
107900=>"110001111",
107901=>"101001100",
107902=>"111101110",
107903=>"010010011",
107904=>"000000000",
107905=>"110011010",
107906=>"011001111",
107907=>"100000110",
107908=>"011001011",
107909=>"101001000",
107910=>"101100010",
107911=>"000100100",
107912=>"001011011",
107913=>"100001001",
107914=>"100000111",
107915=>"111111111",
107916=>"010011000",
107917=>"100110111",
107918=>"010000010",
107919=>"001001011",
107920=>"000000000",
107921=>"010111100",
107922=>"000000000",
107923=>"111101001",
107924=>"000001101",
107925=>"000111111",
107926=>"111111111",
107927=>"000101100",
107928=>"000000000",
107929=>"010101000",
107930=>"011111111",
107931=>"000000111",
107932=>"010101101",
107933=>"111000000",
107934=>"101000000",
107935=>"111000000",
107936=>"111110010",
107937=>"110010000",
107938=>"111101010",
107939=>"111111111",
107940=>"111010000",
107941=>"011001000",
107942=>"101111111",
107943=>"000011010",
107944=>"100000000",
107945=>"000011111",
107946=>"000010010",
107947=>"100100110",
107948=>"000000110",
107949=>"000111101",
107950=>"011111000",
107951=>"010010000",
107952=>"001000000",
107953=>"010111000",
107954=>"100000000",
107955=>"100010011",
107956=>"110101001",
107957=>"110000011",
107958=>"010000010",
107959=>"010011100",
107960=>"110111100",
107961=>"011001001",
107962=>"000100111",
107963=>"001010111",
107964=>"110110001",
107965=>"010111111",
107966=>"100100000",
107967=>"100000101",
107968=>"010010000",
107969=>"000000000",
107970=>"010010001",
107971=>"001001000",
107972=>"000100101",
107973=>"110001110",
107974=>"000100111",
107975=>"111011000",
107976=>"110010011",
107977=>"100000000",
107978=>"101110100",
107979=>"101000100",
107980=>"000100100",
107981=>"010110110",
107982=>"000000001",
107983=>"111111001",
107984=>"010000100",
107985=>"100110000",
107986=>"011111111",
107987=>"111101111",
107988=>"000000000",
107989=>"011001000",
107990=>"001000000",
107991=>"000011111",
107992=>"101100000",
107993=>"000000001",
107994=>"011010011",
107995=>"111000000",
107996=>"001001111",
107997=>"100101101",
107998=>"100000101",
107999=>"000000000",
108000=>"110010000",
108001=>"000010011",
108002=>"101100000",
108003=>"011001000",
108004=>"011000000",
108005=>"010011111",
108006=>"000100010",
108007=>"100011100",
108008=>"000000000",
108009=>"000000101",
108010=>"100000000",
108011=>"111111111",
108012=>"000111000",
108013=>"000101110",
108014=>"000110010",
108015=>"001000000",
108016=>"000100111",
108017=>"110110110",
108018=>"111101011",
108019=>"001001011",
108020=>"000011011",
108021=>"111011100",
108022=>"001000000",
108023=>"100000000",
108024=>"000100000",
108025=>"111111111",
108026=>"000000000",
108027=>"011000000",
108028=>"000000000",
108029=>"000010000",
108030=>"110100110",
108031=>"000000000",
108032=>"000110101",
108033=>"111111001",
108034=>"000010011",
108035=>"000000000",
108036=>"011000100",
108037=>"100000001",
108038=>"000000000",
108039=>"011000000",
108040=>"101101100",
108041=>"000000000",
108042=>"010111111",
108043=>"111001100",
108044=>"010111011",
108045=>"010111001",
108046=>"111100100",
108047=>"110111011",
108048=>"100000100",
108049=>"010111111",
108050=>"000011011",
108051=>"111000000",
108052=>"001111010",
108053=>"000000000",
108054=>"111100000",
108055=>"011111100",
108056=>"000000111",
108057=>"010011111",
108058=>"000000000",
108059=>"000111111",
108060=>"000111011",
108061=>"000000000",
108062=>"111111000",
108063=>"011111000",
108064=>"100000000",
108065=>"111111111",
108066=>"111000000",
108067=>"111000000",
108068=>"111111100",
108069=>"000011010",
108070=>"010111111",
108071=>"000101001",
108072=>"011111111",
108073=>"011111111",
108074=>"000000111",
108075=>"000000000",
108076=>"010111111",
108077=>"000111000",
108078=>"101000011",
108079=>"111101101",
108080=>"100000000",
108081=>"010110000",
108082=>"000000110",
108083=>"011000001",
108084=>"000010010",
108085=>"111111111",
108086=>"000011000",
108087=>"000000000",
108088=>"011000000",
108089=>"111001000",
108090=>"000000001",
108091=>"110000000",
108092=>"000001001",
108093=>"001111111",
108094=>"111000000",
108095=>"000000000",
108096=>"010111010",
108097=>"010000110",
108098=>"000000000",
108099=>"111000000",
108100=>"010111111",
108101=>"000000000",
108102=>"111111011",
108103=>"000000111",
108104=>"011011110",
108105=>"000000000",
108106=>"000000010",
108107=>"101100100",
108108=>"000000100",
108109=>"000011001",
108110=>"110011000",
108111=>"011111111",
108112=>"010111010",
108113=>"001111111",
108114=>"000100000",
108115=>"111001000",
108116=>"000000000",
108117=>"001101000",
108118=>"111111001",
108119=>"111000000",
108120=>"001110000",
108121=>"010111111",
108122=>"010010010",
108123=>"010101100",
108124=>"000000000",
108125=>"110000000",
108126=>"111111010",
108127=>"111101000",
108128=>"100000100",
108129=>"100000000",
108130=>"101011010",
108131=>"001111001",
108132=>"010111001",
108133=>"011111111",
108134=>"000000000",
108135=>"000000001",
108136=>"000000000",
108137=>"000000000",
108138=>"011100100",
108139=>"101011010",
108140=>"000001111",
108141=>"000000000",
108142=>"101100101",
108143=>"010010000",
108144=>"111110110",
108145=>"000000111",
108146=>"001111000",
108147=>"111001111",
108148=>"001100100",
108149=>"000101000",
108150=>"111101000",
108151=>"000010000",
108152=>"101001101",
108153=>"110111000",
108154=>"010010111",
108155=>"010011001",
108156=>"011001001",
108157=>"100000000",
108158=>"100000000",
108159=>"100000000",
108160=>"110000000",
108161=>"000010010",
108162=>"000000000",
108163=>"111110111",
108164=>"010100000",
108165=>"000000100",
108166=>"000000010",
108167=>"011110100",
108168=>"100111111",
108169=>"001001000",
108170=>"000000000",
108171=>"101101001",
108172=>"100000000",
108173=>"100001101",
108174=>"000000101",
108175=>"110000000",
108176=>"010011110",
108177=>"010010000",
108178=>"011101111",
108179=>"101110110",
108180=>"011110000",
108181=>"000010000",
108182=>"000111010",
108183=>"000000000",
108184=>"000101111",
108185=>"010010001",
108186=>"000111111",
108187=>"000000000",
108188=>"100000101",
108189=>"000000000",
108190=>"000000111",
108191=>"101000100",
108192=>"111010110",
108193=>"111111110",
108194=>"111011000",
108195=>"111111111",
108196=>"001100000",
108197=>"110111000",
108198=>"110110111",
108199=>"011101100",
108200=>"111011010",
108201=>"101000100",
108202=>"111111111",
108203=>"111111111",
108204=>"111111111",
108205=>"100100101",
108206=>"100111010",
108207=>"101111011",
108208=>"100000000",
108209=>"100111110",
108210=>"010100000",
108211=>"011000000",
108212=>"010111000",
108213=>"010011111",
108214=>"110000000",
108215=>"000010011",
108216=>"000110110",
108217=>"110001001",
108218=>"000000111",
108219=>"011111111",
108220=>"000000111",
108221=>"000111001",
108222=>"110100100",
108223=>"000011110",
108224=>"011111011",
108225=>"000000101",
108226=>"111111101",
108227=>"111100111",
108228=>"010001111",
108229=>"101110111",
108230=>"110111000",
108231=>"000000000",
108232=>"111111111",
108233=>"000110000",
108234=>"110111111",
108235=>"000111011",
108236=>"111100100",
108237=>"100110100",
108238=>"111111111",
108239=>"000000000",
108240=>"101000001",
108241=>"000110100",
108242=>"101001001",
108243=>"000111001",
108244=>"101101001",
108245=>"001011111",
108246=>"000000000",
108247=>"100001000",
108248=>"011000000",
108249=>"010110010",
108250=>"111011101",
108251=>"000110110",
108252=>"110011000",
108253=>"011001100",
108254=>"000000000",
108255=>"111111111",
108256=>"010111011",
108257=>"010111111",
108258=>"000000000",
108259=>"111111111",
108260=>"111000101",
108261=>"101100000",
108262=>"101000000",
108263=>"011101000",
108264=>"011111111",
108265=>"111111110",
108266=>"000011011",
108267=>"111111111",
108268=>"000011111",
108269=>"111000000",
108270=>"100111010",
108271=>"100000000",
108272=>"100111111",
108273=>"101001001",
108274=>"111101000",
108275=>"110111010",
108276=>"101001101",
108277=>"011111111",
108278=>"001000100",
108279=>"000000100",
108280=>"111100000",
108281=>"011000000",
108282=>"000011111",
108283=>"111111000",
108284=>"000111000",
108285=>"111000000",
108286=>"011111001",
108287=>"000000000",
108288=>"011100100",
108289=>"111010000",
108290=>"111100101",
108291=>"001000111",
108292=>"010000000",
108293=>"000001111",
108294=>"001111111",
108295=>"010111111",
108296=>"000001111",
108297=>"000101111",
108298=>"111010000",
108299=>"001101100",
108300=>"000000111",
108301=>"111111111",
108302=>"000111110",
108303=>"101111110",
108304=>"111111000",
108305=>"011110000",
108306=>"010000110",
108307=>"001000001",
108308=>"111110110",
108309=>"000000111",
108310=>"101011111",
108311=>"011010000",
108312=>"000000111",
108313=>"001111111",
108314=>"100111111",
108315=>"111110000",
108316=>"110111111",
108317=>"100000000",
108318=>"101000000",
108319=>"100111111",
108320=>"111001001",
108321=>"111111111",
108322=>"000110111",
108323=>"000111111",
108324=>"000000100",
108325=>"011000010",
108326=>"011000010",
108327=>"000011001",
108328=>"110000110",
108329=>"111111000",
108330=>"000110110",
108331=>"000011111",
108332=>"111111010",
108333=>"111000000",
108334=>"111000000",
108335=>"000011111",
108336=>"000000000",
108337=>"100100000",
108338=>"111111111",
108339=>"001100000",
108340=>"111111000",
108341=>"000000000",
108342=>"011000010",
108343=>"000001111",
108344=>"101010111",
108345=>"000000001",
108346=>"000010000",
108347=>"000111110",
108348=>"000001110",
108349=>"111000110",
108350=>"000000001",
108351=>"000001100",
108352=>"100000000",
108353=>"001101111",
108354=>"000111111",
108355=>"000101111",
108356=>"000000000",
108357=>"101000000",
108358=>"110010000",
108359=>"111110011",
108360=>"110001111",
108361=>"101111010",
108362=>"100001111",
108363=>"001001011",
108364=>"001000101",
108365=>"100000000",
108366=>"011001101",
108367=>"000100000",
108368=>"000000000",
108369=>"111101111",
108370=>"101111111",
108371=>"001000000",
108372=>"011010000",
108373=>"010110011",
108374=>"110011011",
108375=>"000000000",
108376=>"001111111",
108377=>"000000011",
108378=>"111111000",
108379=>"000000111",
108380=>"110000000",
108381=>"001111111",
108382=>"111000000",
108383=>"001000110",
108384=>"000111111",
108385=>"010111111",
108386=>"000101111",
108387=>"111001000",
108388=>"100001101",
108389=>"011011111",
108390=>"111111100",
108391=>"000100000",
108392=>"000000111",
108393=>"101000100",
108394=>"011111111",
108395=>"010010111",
108396=>"110010110",
108397=>"111111000",
108398=>"000001111",
108399=>"111111111",
108400=>"111111011",
108401=>"000011000",
108402=>"000000000",
108403=>"000000000",
108404=>"000000000",
108405=>"000101001",
108406=>"111111111",
108407=>"000111111",
108408=>"111000000",
108409=>"101010111",
108410=>"011110111",
108411=>"000000111",
108412=>"100001000",
108413=>"100000000",
108414=>"110000011",
108415=>"000000111",
108416=>"000000000",
108417=>"000000111",
108418=>"100111111",
108419=>"111111110",
108420=>"000000010",
108421=>"000000101",
108422=>"110100000",
108423=>"000000000",
108424=>"011010111",
108425=>"111000000",
108426=>"011011000",
108427=>"000000101",
108428=>"111001111",
108429=>"001101111",
108430=>"100110111",
108431=>"000001111",
108432=>"111111011",
108433=>"111011111",
108434=>"011000000",
108435=>"111100000",
108436=>"111000000",
108437=>"000111111",
108438=>"001100010",
108439=>"101100111",
108440=>"000000100",
108441=>"000001000",
108442=>"010110111",
108443=>"000001000",
108444=>"100100111",
108445=>"100101111",
108446=>"010010011",
108447=>"000111111",
108448=>"000001011",
108449=>"010000000",
108450=>"110101111",
108451=>"000110101",
108452=>"111101110",
108453=>"110000010",
108454=>"101000110",
108455=>"000000000",
108456=>"111111011",
108457=>"101100010",
108458=>"000101111",
108459=>"001011000",
108460=>"111110111",
108461=>"000001111",
108462=>"100001011",
108463=>"000000111",
108464=>"001100000",
108465=>"100100111",
108466=>"101101000",
108467=>"000110111",
108468=>"111100000",
108469=>"011000000",
108470=>"100011001",
108471=>"011100000",
108472=>"000110111",
108473=>"111011000",
108474=>"000000000",
108475=>"111110111",
108476=>"000100111",
108477=>"000111111",
108478=>"000000110",
108479=>"000000000",
108480=>"010010000",
108481=>"000001000",
108482=>"001001000",
108483=>"001011011",
108484=>"000000000",
108485=>"011000100",
108486=>"010000000",
108487=>"001111010",
108488=>"000111111",
108489=>"001001011",
108490=>"001111100",
108491=>"000011000",
108492=>"011000000",
108493=>"100100010",
108494=>"000000000",
108495=>"000001111",
108496=>"000000000",
108497=>"011011111",
108498=>"000000111",
108499=>"111100010",
108500=>"000110111",
108501=>"110011000",
108502=>"111000000",
108503=>"100000000",
108504=>"111000000",
108505=>"001111111",
108506=>"000000100",
108507=>"000001111",
108508=>"111010110",
108509=>"100100111",
108510=>"101111010",
108511=>"111111000",
108512=>"111100101",
108513=>"100110111",
108514=>"000000001",
108515=>"010011011",
108516=>"011000000",
108517=>"000000111",
108518=>"001000111",
108519=>"110000111",
108520=>"000000010",
108521=>"111101001",
108522=>"111010000",
108523=>"101111111",
108524=>"000010101",
108525=>"001000000",
108526=>"011000000",
108527=>"000100100",
108528=>"001111101",
108529=>"011101000",
108530=>"001101011",
108531=>"111101100",
108532=>"001000011",
108533=>"111000000",
108534=>"000000111",
108535=>"111101000",
108536=>"011000111",
108537=>"110000110",
108538=>"100111111",
108539=>"111000010",
108540=>"000100010",
108541=>"000001011",
108542=>"001001111",
108543=>"000011010",
108544=>"111010010",
108545=>"111001000",
108546=>"101101111",
108547=>"111010000",
108548=>"110111110",
108549=>"001111110",
108550=>"000111100",
108551=>"001011110",
108552=>"010011001",
108553=>"000101110",
108554=>"101001001",
108555=>"000000100",
108556=>"011000000",
108557=>"100101001",
108558=>"011110100",
108559=>"001000000",
108560=>"000110001",
108561=>"001000000",
108562=>"101010010",
108563=>"011111001",
108564=>"101101101",
108565=>"000000101",
108566=>"111010111",
108567=>"000000000",
108568=>"000111101",
108569=>"110111101",
108570=>"011111101",
108571=>"010101100",
108572=>"000000100",
108573=>"111100101",
108574=>"001011100",
108575=>"111000000",
108576=>"010111111",
108577=>"100000001",
108578=>"111101101",
108579=>"000011000",
108580=>"010011010",
108581=>"011011111",
108582=>"100101111",
108583=>"111111111",
108584=>"100101111",
108585=>"000000010",
108586=>"111100000",
108587=>"100000000",
108588=>"011000010",
108589=>"000000000",
108590=>"111000000",
108591=>"010010000",
108592=>"000010100",
108593=>"010111011",
108594=>"001010111",
108595=>"111111101",
108596=>"001000000",
108597=>"000001100",
108598=>"001011000",
108599=>"110010000",
108600=>"101011001",
108601=>"111111000",
108602=>"100100011",
108603=>"000000111",
108604=>"111010011",
108605=>"001010111",
108606=>"100101101",
108607=>"010011101",
108608=>"101010111",
108609=>"101111111",
108610=>"011111111",
108611=>"100010011",
108612=>"010111011",
108613=>"000000111",
108614=>"111111011",
108615=>"011011011",
108616=>"100010011",
108617=>"111001101",
108618=>"011100000",
108619=>"011000110",
108620=>"010101111",
108621=>"010110111",
108622=>"000110111",
108623=>"101101000",
108624=>"010010001",
108625=>"111111111",
108626=>"011000000",
108627=>"011011001",
108628=>"010100110",
108629=>"111110001",
108630=>"101010001",
108631=>"001101101",
108632=>"111111011",
108633=>"011010110",
108634=>"111100000",
108635=>"110000000",
108636=>"011000101",
108637=>"101100110",
108638=>"111101111",
108639=>"001010100",
108640=>"010010110",
108641=>"011011000",
108642=>"100100110",
108643=>"111011000",
108644=>"111000000",
108645=>"110010110",
108646=>"111001001",
108647=>"100100100",
108648=>"010010111",
108649=>"000111111",
108650=>"000111111",
108651=>"000000000",
108652=>"000011001",
108653=>"000000000",
108654=>"110111111",
108655=>"000011011",
108656=>"011011111",
108657=>"000111111",
108658=>"110110011",
108659=>"011111111",
108660=>"000111000",
108661=>"000000000",
108662=>"010111001",
108663=>"001101101",
108664=>"001101111",
108665=>"101011100",
108666=>"111101100",
108667=>"001011011",
108668=>"100010001",
108669=>"101110110",
108670=>"000010111",
108671=>"111010111",
108672=>"000111110",
108673=>"001010000",
108674=>"000101100",
108675=>"111011000",
108676=>"000010010",
108677=>"000000000",
108678=>"110110111",
108679=>"111011110",
108680=>"110110110",
108681=>"011010111",
108682=>"100111000",
108683=>"011000010",
108684=>"110101111",
108685=>"100110111",
108686=>"111010111",
108687=>"000110010",
108688=>"111110011",
108689=>"100111111",
108690=>"110100011",
108691=>"111111101",
108692=>"010111000",
108693=>"000101101",
108694=>"101110000",
108695=>"001001010",
108696=>"111111010",
108697=>"011000000",
108698=>"111110111",
108699=>"000110000",
108700=>"010111101",
108701=>"000010011",
108702=>"110100001",
108703=>"001000000",
108704=>"000010101",
108705=>"011110100",
108706=>"000000000",
108707=>"101111111",
108708=>"010110111",
108709=>"010110001",
108710=>"110010101",
108711=>"111101101",
108712=>"111111001",
108713=>"000001111",
108714=>"100100000",
108715=>"000010001",
108716=>"111101011",
108717=>"000100111",
108718=>"000010000",
108719=>"111000001",
108720=>"110000000",
108721=>"001000011",
108722=>"101111111",
108723=>"110111001",
108724=>"111010110",
108725=>"000000011",
108726=>"111001000",
108727=>"001111100",
108728=>"000010110",
108729=>"110011001",
108730=>"010111111",
108731=>"111101000",
108732=>"101000000",
108733=>"001111111",
108734=>"110110110",
108735=>"101001101",
108736=>"111100000",
108737=>"111000000",
108738=>"011010000",
108739=>"010010010",
108740=>"000000000",
108741=>"011000000",
108742=>"101011000",
108743=>"111000000",
108744=>"101111101",
108745=>"111110101",
108746=>"010000000",
108747=>"011010111",
108748=>"000000000",
108749=>"101010100",
108750=>"110000000",
108751=>"010111000",
108752=>"010110000",
108753=>"110110110",
108754=>"111111101",
108755=>"001000000",
108756=>"111000101",
108757=>"100010000",
108758=>"111101000",
108759=>"010010000",
108760=>"101000000",
108761=>"111000101",
108762=>"110100001",
108763=>"111101101",
108764=>"000010101",
108765=>"000000000",
108766=>"111011111",
108767=>"001101000",
108768=>"000111000",
108769=>"000000000",
108770=>"101100000",
108771=>"011011011",
108772=>"000101101",
108773=>"010010010",
108774=>"000011111",
108775=>"000010000",
108776=>"100111111",
108777=>"010000101",
108778=>"101101100",
108779=>"111101000",
108780=>"000101101",
108781=>"000111100",
108782=>"000101111",
108783=>"000010000",
108784=>"000000000",
108785=>"111000001",
108786=>"001000101",
108787=>"011011000",
108788=>"001001010",
108789=>"111000001",
108790=>"000000100",
108791=>"111111111",
108792=>"101100101",
108793=>"111111101",
108794=>"010110101",
108795=>"111111000",
108796=>"010010000",
108797=>"111000110",
108798=>"011011101",
108799=>"010000000",
108800=>"001101000",
108801=>"000010010",
108802=>"001000111",
108803=>"000000101",
108804=>"001011000",
108805=>"110111111",
108806=>"001111000",
108807=>"000001111",
108808=>"000000000",
108809=>"000000000",
108810=>"110100100",
108811=>"110111000",
108812=>"000000000",
108813=>"110110100",
108814=>"011111111",
108815=>"111111111",
108816=>"000000000",
108817=>"000100000",
108818=>"000000010",
108819=>"011010000",
108820=>"101010000",
108821=>"111001111",
108822=>"110100111",
108823=>"010111101",
108824=>"000000000",
108825=>"111110110",
108826=>"000010011",
108827=>"000000111",
108828=>"000000101",
108829=>"000000010",
108830=>"011010011",
108831=>"000010010",
108832=>"110000111",
108833=>"000010000",
108834=>"111001111",
108835=>"000000000",
108836=>"001000001",
108837=>"100110100",
108838=>"000100000",
108839=>"111101001",
108840=>"101010111",
108841=>"100100000",
108842=>"000100000",
108843=>"010000000",
108844=>"000010100",
108845=>"011010000",
108846=>"111010010",
108847=>"111111011",
108848=>"110110000",
108849=>"100001011",
108850=>"011010000",
108851=>"000101101",
108852=>"111111000",
108853=>"110000110",
108854=>"111111011",
108855=>"010111111",
108856=>"000011011",
108857=>"000000101",
108858=>"000000111",
108859=>"111101100",
108860=>"100110110",
108861=>"111111010",
108862=>"000000000",
108863=>"011011100",
108864=>"000111101",
108865=>"010111000",
108866=>"100101001",
108867=>"111111000",
108868=>"010000000",
108869=>"000100000",
108870=>"000111100",
108871=>"101111111",
108872=>"010011011",
108873=>"000010000",
108874=>"010000000",
108875=>"000001010",
108876=>"010010000",
108877=>"011011010",
108878=>"000100000",
108879=>"000001000",
108880=>"000111111",
108881=>"111110000",
108882=>"011010100",
108883=>"000110000",
108884=>"100000010",
108885=>"110000001",
108886=>"010011110",
108887=>"010000111",
108888=>"000110111",
108889=>"000001111",
108890=>"111111011",
108891=>"100100111",
108892=>"010000000",
108893=>"010000011",
108894=>"111001000",
108895=>"101100101",
108896=>"000110111",
108897=>"000111111",
108898=>"111100111",
108899=>"001101110",
108900=>"000010000",
108901=>"111100110",
108902=>"100110011",
108903=>"111011011",
108904=>"101000011",
108905=>"101101111",
108906=>"110101101",
108907=>"000111111",
108908=>"010000101",
108909=>"101101101",
108910=>"111101001",
108911=>"000111111",
108912=>"001111110",
108913=>"000000111",
108914=>"010101110",
108915=>"011000000",
108916=>"010100000",
108917=>"100101101",
108918=>"000101100",
108919=>"010110111",
108920=>"000100100",
108921=>"011101111",
108922=>"011111111",
108923=>"001001001",
108924=>"100100010",
108925=>"000010000",
108926=>"001101111",
108927=>"000000110",
108928=>"000001101",
108929=>"011100000",
108930=>"010010010",
108931=>"000000001",
108932=>"000010000",
108933=>"001001111",
108934=>"001011000",
108935=>"100100110",
108936=>"100100011",
108937=>"111101100",
108938=>"101101000",
108939=>"000010111",
108940=>"000110111",
108941=>"101101111",
108942=>"010101111",
108943=>"000001001",
108944=>"011001011",
108945=>"001111111",
108946=>"100000000",
108947=>"000111111",
108948=>"100101111",
108949=>"000000111",
108950=>"010011110",
108951=>"000010000",
108952=>"111101001",
108953=>"011011000",
108954=>"100010010",
108955=>"111101101",
108956=>"111101100",
108957=>"111011110",
108958=>"101000010",
108959=>"000000000",
108960=>"010000100",
108961=>"101000000",
108962=>"101101111",
108963=>"000110000",
108964=>"010111111",
108965=>"011100110",
108966=>"000000110",
108967=>"000110100",
108968=>"010010000",
108969=>"100100001",
108970=>"101000000",
108971=>"110101000",
108972=>"000000011",
108973=>"000100100",
108974=>"110100100",
108975=>"101111000",
108976=>"000000010",
108977=>"110101011",
108978=>"011110000",
108979=>"100110110",
108980=>"100111011",
108981=>"110011010",
108982=>"000001001",
108983=>"011000010",
108984=>"001001011",
108985=>"001001011",
108986=>"000011011",
108987=>"011110000",
108988=>"000000000",
108989=>"111111111",
108990=>"000100101",
108991=>"000011010",
108992=>"010010000",
108993=>"000001101",
108994=>"101010000",
108995=>"011010111",
108996=>"010111000",
108997=>"111111110",
108998=>"000111111",
108999=>"111100111",
109000=>"100100000",
109001=>"000001011",
109002=>"111100101",
109003=>"000100110",
109004=>"001100000",
109005=>"101001011",
109006=>"100000010",
109007=>"111000101",
109008=>"100111000",
109009=>"000110110",
109010=>"101010111",
109011=>"010000111",
109012=>"000010111",
109013=>"000000000",
109014=>"010000101",
109015=>"101000011",
109016=>"110111000",
109017=>"000111111",
109018=>"001000001",
109019=>"101101101",
109020=>"001000110",
109021=>"001000000",
109022=>"000111111",
109023=>"000010000",
109024=>"100101000",
109025=>"111101000",
109026=>"111001001",
109027=>"011001001",
109028=>"000000000",
109029=>"000010101",
109030=>"111101101",
109031=>"111010100",
109032=>"100101101",
109033=>"111000000",
109034=>"111001001",
109035=>"000000110",
109036=>"000000000",
109037=>"101010000",
109038=>"111000000",
109039=>"111000011",
109040=>"100000011",
109041=>"111011010",
109042=>"010000000",
109043=>"001110110",
109044=>"110110000",
109045=>"111001101",
109046=>"000010010",
109047=>"100100010",
109048=>"111110110",
109049=>"000000101",
109050=>"111110110",
109051=>"101100001",
109052=>"111000100",
109053=>"010101000",
109054=>"100100111",
109055=>"111001100",
109056=>"011011001",
109057=>"000001100",
109058=>"100000101",
109059=>"010100100",
109060=>"010001011",
109061=>"111110000",
109062=>"101000111",
109063=>"000010011",
109064=>"000011111",
109065=>"000000111",
109066=>"101001001",
109067=>"001000011",
109068=>"000000000",
109069=>"100111101",
109070=>"100001011",
109071=>"110001111",
109072=>"100110101",
109073=>"100100010",
109074=>"111110111",
109075=>"111100100",
109076=>"110101111",
109077=>"000100000",
109078=>"110100101",
109079=>"101101111",
109080=>"000000000",
109081=>"011000000",
109082=>"000011000",
109083=>"011011111",
109084=>"000100111",
109085=>"010011000",
109086=>"111101101",
109087=>"100100000",
109088=>"000000100",
109089=>"111100010",
109090=>"111101001",
109091=>"000011000",
109092=>"011011001",
109093=>"110111011",
109094=>"000010010",
109095=>"000001110",
109096=>"101000101",
109097=>"000111111",
109098=>"100000000",
109099=>"100000100",
109100=>"111000101",
109101=>"000101111",
109102=>"011000101",
109103=>"010100100",
109104=>"001000110",
109105=>"101100011",
109106=>"000010111",
109107=>"000100001",
109108=>"000000111",
109109=>"000000000",
109110=>"100100111",
109111=>"000000000",
109112=>"011000011",
109113=>"101100111",
109114=>"100000110",
109115=>"000100000",
109116=>"010010000",
109117=>"111111000",
109118=>"100100011",
109119=>"011111110",
109120=>"011111111",
109121=>"110111111",
109122=>"111111011",
109123=>"010010000",
109124=>"011111101",
109125=>"111101101",
109126=>"001011111",
109127=>"010000110",
109128=>"101001111",
109129=>"000000000",
109130=>"001000101",
109131=>"111000011",
109132=>"111111111",
109133=>"101001001",
109134=>"100000000",
109135=>"101111111",
109136=>"100000100",
109137=>"110111111",
109138=>"101111111",
109139=>"001101101",
109140=>"000011011",
109141=>"011111111",
109142=>"111010110",
109143=>"000111111",
109144=>"100000011",
109145=>"011110100",
109146=>"100100000",
109147=>"110110000",
109148=>"000101100",
109149=>"001000001",
109150=>"010111111",
109151=>"100010001",
109152=>"000111010",
109153=>"011111000",
109154=>"101111010",
109155=>"001000111",
109156=>"000000001",
109157=>"100001010",
109158=>"000000111",
109159=>"100000000",
109160=>"111101000",
109161=>"111010111",
109162=>"111011101",
109163=>"010001101",
109164=>"010010101",
109165=>"000100100",
109166=>"100000000",
109167=>"111000001",
109168=>"100111011",
109169=>"000001011",
109170=>"000001011",
109171=>"111111001",
109172=>"111111111",
109173=>"000000101",
109174=>"010000011",
109175=>"101101111",
109176=>"011001011",
109177=>"111111000",
109178=>"111101101",
109179=>"111101100",
109180=>"100000011",
109181=>"110100100",
109182=>"000101010",
109183=>"111110110",
109184=>"111101100",
109185=>"111000010",
109186=>"011011110",
109187=>"111011101",
109188=>"000101101",
109189=>"111001011",
109190=>"011011111",
109191=>"000000100",
109192=>"100100100",
109193=>"011111100",
109194=>"100100111",
109195=>"010000000",
109196=>"000000000",
109197=>"001111100",
109198=>"011010010",
109199=>"001000000",
109200=>"010000000",
109201=>"010010000",
109202=>"000000000",
109203=>"101101111",
109204=>"000000111",
109205=>"000001111",
109206=>"010111111",
109207=>"000011011",
109208=>"110111000",
109209=>"100000111",
109210=>"000000010",
109211=>"000011010",
109212=>"000100010",
109213=>"011000000",
109214=>"010000110",
109215=>"000000110",
109216=>"001110100",
109217=>"010000010",
109218=>"100111111",
109219=>"111111111",
109220=>"111111000",
109221=>"011011001",
109222=>"110110011",
109223=>"111111011",
109224=>"010000101",
109225=>"000010111",
109226=>"100111111",
109227=>"010000000",
109228=>"111111011",
109229=>"101000110",
109230=>"100000010",
109231=>"111100101",
109232=>"000100000",
109233=>"000100000",
109234=>"000000000",
109235=>"111001000",
109236=>"110110100",
109237=>"111100000",
109238=>"100110100",
109239=>"000000000",
109240=>"110110110",
109241=>"000001001",
109242=>"110000100",
109243=>"111000000",
109244=>"111000011",
109245=>"110011010",
109246=>"111111001",
109247=>"101100110",
109248=>"100000000",
109249=>"101000101",
109250=>"000000101",
109251=>"001110100",
109252=>"101001001",
109253=>"100000111",
109254=>"010110100",
109255=>"100000101",
109256=>"100000010",
109257=>"000100000",
109258=>"111101000",
109259=>"111101000",
109260=>"111100000",
109261=>"001000111",
109262=>"101101111",
109263=>"010111000",
109264=>"000000011",
109265=>"110110111",
109266=>"000000000",
109267=>"111111111",
109268=>"000001101",
109269=>"100110000",
109270=>"100110111",
109271=>"000111111",
109272=>"100100111",
109273=>"111000000",
109274=>"101101001",
109275=>"000000000",
109276=>"111011111",
109277=>"000011111",
109278=>"111111111",
109279=>"100101110",
109280=>"000000000",
109281=>"000000100",
109282=>"100100111",
109283=>"001111100",
109284=>"101000000",
109285=>"010010011",
109286=>"010110111",
109287=>"010001000",
109288=>"000111101",
109289=>"100111111",
109290=>"111100100",
109291=>"110100100",
109292=>"000011010",
109293=>"101011010",
109294=>"000000000",
109295=>"000010000",
109296=>"111111100",
109297=>"000000011",
109298=>"010001101",
109299=>"010001011",
109300=>"111110111",
109301=>"100101111",
109302=>"000000000",
109303=>"110000001",
109304=>"000000111",
109305=>"100001000",
109306=>"100100101",
109307=>"000000111",
109308=>"111010000",
109309=>"000000000",
109310=>"110110100",
109311=>"100000011",
109312=>"111000100",
109313=>"010011010",
109314=>"000000101",
109315=>"110010000",
109316=>"111001100",
109317=>"100100111",
109318=>"111000011",
109319=>"111011111",
109320=>"011101111",
109321=>"101100100",
109322=>"000010010",
109323=>"100101000",
109324=>"000000100",
109325=>"000000010",
109326=>"101001000",
109327=>"101001111",
109328=>"111001001",
109329=>"101000000",
109330=>"101101111",
109331=>"000000001",
109332=>"000000010",
109333=>"000000100",
109334=>"000010011",
109335=>"001111000",
109336=>"000000000",
109337=>"000000100",
109338=>"100100000",
109339=>"111000000",
109340=>"100110101",
109341=>"111111111",
109342=>"001000001",
109343=>"011010010",
109344=>"000000110",
109345=>"110101111",
109346=>"000010110",
109347=>"000000111",
109348=>"001001111",
109349=>"110000001",
109350=>"000010000",
109351=>"111111111",
109352=>"100100010",
109353=>"100000000",
109354=>"101101001",
109355=>"100000111",
109356=>"000011101",
109357=>"010010000",
109358=>"010010010",
109359=>"010000000",
109360=>"111101101",
109361=>"011000110",
109362=>"101000111",
109363=>"100000101",
109364=>"010010010",
109365=>"000111111",
109366=>"000011010",
109367=>"011010000",
109368=>"100001111",
109369=>"011011000",
109370=>"101101101",
109371=>"101100111",
109372=>"111111011",
109373=>"111111011",
109374=>"001000000",
109375=>"010100110",
109376=>"000000111",
109377=>"000000100",
109378=>"111000000",
109379=>"111001100",
109380=>"111111000",
109381=>"111100101",
109382=>"000100100",
109383=>"111001000",
109384=>"111111111",
109385=>"111111011",
109386=>"010010000",
109387=>"111011101",
109388=>"101000101",
109389=>"000100110",
109390=>"110110000",
109391=>"000100111",
109392=>"010010010",
109393=>"111111010",
109394=>"111111010",
109395=>"101101100",
109396=>"000011111",
109397=>"100110110",
109398=>"100111111",
109399=>"000100010",
109400=>"101110110",
109401=>"001100100",
109402=>"000001001",
109403=>"111100111",
109404=>"110100000",
109405=>"111011011",
109406=>"111101011",
109407=>"110100001",
109408=>"000000000",
109409=>"001000000",
109410=>"100001101",
109411=>"000100000",
109412=>"110000001",
109413=>"111011111",
109414=>"011010011",
109415=>"111100010",
109416=>"001111111",
109417=>"101000110",
109418=>"101101111",
109419=>"111101101",
109420=>"101111111",
109421=>"101100000",
109422=>"010000000",
109423=>"010100101",
109424=>"000000000",
109425=>"111100101",
109426=>"000010110",
109427=>"010111011",
109428=>"010010000",
109429=>"001000101",
109430=>"010000001",
109431=>"000000100",
109432=>"001000000",
109433=>"011000000",
109434=>"011011100",
109435=>"010000011",
109436=>"110111110",
109437=>"111100110",
109438=>"001101111",
109439=>"001101000",
109440=>"101000111",
109441=>"110011011",
109442=>"100000111",
109443=>"011000011",
109444=>"000000000",
109445=>"101111111",
109446=>"000100110",
109447=>"000010001",
109448=>"010110000",
109449=>"010111111",
109450=>"001000000",
109451=>"111000100",
109452=>"011100010",
109453=>"000000111",
109454=>"100100101",
109455=>"000000000",
109456=>"110100110",
109457=>"001100000",
109458=>"001101111",
109459=>"010111111",
109460=>"001010000",
109461=>"000000100",
109462=>"000110001",
109463=>"000100100",
109464=>"000101111",
109465=>"100111111",
109466=>"100000101",
109467=>"100101101",
109468=>"011101101",
109469=>"100100101",
109470=>"000001111",
109471=>"110111111",
109472=>"011011011",
109473=>"101011111",
109474=>"010011101",
109475=>"101100110",
109476=>"111011000",
109477=>"100000111",
109478=>"111111000",
109479=>"000101100",
109480=>"010111101",
109481=>"000111100",
109482=>"101101100",
109483=>"000101100",
109484=>"000010010",
109485=>"001100101",
109486=>"010000011",
109487=>"110011000",
109488=>"011000000",
109489=>"011011011",
109490=>"111100000",
109491=>"110001100",
109492=>"111011110",
109493=>"100100111",
109494=>"000000011",
109495=>"100100101",
109496=>"111111111",
109497=>"001011001",
109498=>"110000011",
109499=>"010101101",
109500=>"000000111",
109501=>"101101001",
109502=>"100001011",
109503=>"000010111",
109504=>"001100000",
109505=>"000100111",
109506=>"110010000",
109507=>"000000000",
109508=>"010100110",
109509=>"010001000",
109510=>"000101011",
109511=>"000000000",
109512=>"010111111",
109513=>"000011010",
109514=>"000010100",
109515=>"000100111",
109516=>"011100100",
109517=>"111011010",
109518=>"000000000",
109519=>"010101111",
109520=>"001101011",
109521=>"010000011",
109522=>"110100000",
109523=>"000000011",
109524=>"101001000",
109525=>"110110000",
109526=>"111111100",
109527=>"000010110",
109528=>"000110101",
109529=>"011111000",
109530=>"100100110",
109531=>"101100101",
109532=>"000000000",
109533=>"111010111",
109534=>"000000010",
109535=>"111101011",
109536=>"000101111",
109537=>"010001000",
109538=>"111110000",
109539=>"110001001",
109540=>"101100100",
109541=>"111111110",
109542=>"110111111",
109543=>"000100100",
109544=>"111001000",
109545=>"001000001",
109546=>"010011000",
109547=>"100100000",
109548=>"010010100",
109549=>"000111110",
109550=>"001000000",
109551=>"111101101",
109552=>"100101111",
109553=>"011101000",
109554=>"010010000",
109555=>"110100111",
109556=>"010000001",
109557=>"000010011",
109558=>"101100101",
109559=>"100000110",
109560=>"101101111",
109561=>"100111111",
109562=>"111000000",
109563=>"000100000",
109564=>"000101111",
109565=>"111100000",
109566=>"110000000",
109567=>"100010000",
109568=>"010000100",
109569=>"100101000",
109570=>"001001001",
109571=>"000001111",
109572=>"110111001",
109573=>"000010010",
109574=>"000111111",
109575=>"101111111",
109576=>"010000000",
109577=>"111111000",
109578=>"000000010",
109579=>"111110101",
109580=>"000110110",
109581=>"010011010",
109582=>"111111111",
109583=>"110000000",
109584=>"111101011",
109585=>"001111111",
109586=>"001000010",
109587=>"000101111",
109588=>"000000001",
109589=>"000111111",
109590=>"111100000",
109591=>"110111111",
109592=>"000000001",
109593=>"111111111",
109594=>"111101110",
109595=>"111111011",
109596=>"111111111",
109597=>"111111000",
109598=>"000000000",
109599=>"000000101",
109600=>"010100000",
109601=>"010000001",
109602=>"111010111",
109603=>"111000000",
109604=>"100101000",
109605=>"100000001",
109606=>"111100000",
109607=>"110000000",
109608=>"111110011",
109609=>"111111000",
109610=>"111111111",
109611=>"110111110",
109612=>"000111000",
109613=>"000000000",
109614=>"111111000",
109615=>"110111000",
109616=>"101011000",
109617=>"000000000",
109618=>"000000100",
109619=>"000111111",
109620=>"111111000",
109621=>"111110101",
109622=>"001001011",
109623=>"000111011",
109624=>"000000101",
109625=>"000000111",
109626=>"000000111",
109627=>"111111111",
109628=>"110000001",
109629=>"001111111",
109630=>"000111111",
109631=>"011000000",
109632=>"111111111",
109633=>"000000000",
109634=>"000010000",
109635=>"111011000",
109636=>"001000000",
109637=>"000000000",
109638=>"111110110",
109639=>"000111111",
109640=>"000000000",
109641=>"011000000",
109642=>"000010000",
109643=>"111111111",
109644=>"001111111",
109645=>"000100000",
109646=>"000000000",
109647=>"110011011",
109648=>"111110110",
109649=>"000011111",
109650=>"000000011",
109651=>"000100110",
109652=>"000010000",
109653=>"100001001",
109654=>"101110000",
109655=>"000111111",
109656=>"000000101",
109657=>"001000101",
109658=>"101101000",
109659=>"000111111",
109660=>"000011000",
109661=>"000001011",
109662=>"010000000",
109663=>"011111100",
109664=>"111110111",
109665=>"001000000",
109666=>"000111111",
109667=>"110011001",
109668=>"100100001",
109669=>"100011001",
109670=>"000000001",
109671=>"010101001",
109672=>"111011111",
109673=>"000110111",
109674=>"000000010",
109675=>"000100101",
109676=>"111101001",
109677=>"000110111",
109678=>"111111110",
109679=>"110111110",
109680=>"110111110",
109681=>"001111111",
109682=>"100110110",
109683=>"000000010",
109684=>"000000101",
109685=>"000000101",
109686=>"111111111",
109687=>"000000001",
109688=>"000111111",
109689=>"000000000",
109690=>"000000000",
109691=>"101000111",
109692=>"011111111",
109693=>"000001011",
109694=>"000000000",
109695=>"111001000",
109696=>"110000001",
109697=>"111111010",
109698=>"111000000",
109699=>"101000000",
109700=>"101001000",
109701=>"000000000",
109702=>"011000000",
109703=>"101111101",
109704=>"001100110",
109705=>"111111111",
109706=>"111010010",
109707=>"000101001",
109708=>"111101000",
109709=>"110110100",
109710=>"000111101",
109711=>"111111100",
109712=>"000000111",
109713=>"100000100",
109714=>"000001001",
109715=>"111111101",
109716=>"001101111",
109717=>"111111001",
109718=>"010010010",
109719=>"100000000",
109720=>"111111111",
109721=>"000001001",
109722=>"111111111",
109723=>"111111110",
109724=>"100110000",
109725=>"111111111",
109726=>"000010101",
109727=>"111111111",
109728=>"000000000",
109729=>"111111010",
109730=>"111111111",
109731=>"111010101",
109732=>"000010011",
109733=>"101111111",
109734=>"000001000",
109735=>"111111101",
109736=>"110010000",
109737=>"010000000",
109738=>"011011011",
109739=>"101101111",
109740=>"010000011",
109741=>"000000001",
109742=>"001001001",
109743=>"000010010",
109744=>"000000010",
109745=>"110110100",
109746=>"000000011",
109747=>"111111111",
109748=>"000000011",
109749=>"000000000",
109750=>"100100110",
109751=>"010101000",
109752=>"000000100",
109753=>"100111110",
109754=>"111001001",
109755=>"111111101",
109756=>"111100101",
109757=>"000000000",
109758=>"110110010",
109759=>"111111000",
109760=>"000010010",
109761=>"101111111",
109762=>"010000000",
109763=>"001011001",
109764=>"110111110",
109765=>"010010001",
109766=>"000000011",
109767=>"000110010",
109768=>"111111111",
109769=>"000000010",
109770=>"011011010",
109771=>"000000101",
109772=>"110101110",
109773=>"111111101",
109774=>"111111111",
109775=>"111111111",
109776=>"000000000",
109777=>"000010000",
109778=>"111111111",
109779=>"110110101",
109780=>"111101111",
109781=>"111111111",
109782=>"000000000",
109783=>"101001110",
109784=>"001111001",
109785=>"011000000",
109786=>"000001011",
109787=>"111111111",
109788=>"111011000",
109789=>"000000000",
109790=>"110111100",
109791=>"000000001",
109792=>"111111000",
109793=>"111110000",
109794=>"000000000",
109795=>"111111111",
109796=>"000111101",
109797=>"110111101",
109798=>"100000111",
109799=>"001000000",
109800=>"000000000",
109801=>"110111000",
109802=>"000001011",
109803=>"011001000",
109804=>"111110000",
109805=>"111001000",
109806=>"010011001",
109807=>"111111011",
109808=>"111111111",
109809=>"010001100",
109810=>"011110000",
109811=>"000000000",
109812=>"000100011",
109813=>"111111001",
109814=>"101101111",
109815=>"101111100",
109816=>"111101101",
109817=>"000000000",
109818=>"111111111",
109819=>"110010001",
109820=>"111111111",
109821=>"111111111",
109822=>"101011111",
109823=>"111111111",
109824=>"000010000",
109825=>"011010100",
109826=>"100000000",
109827=>"110000000",
109828=>"011111001",
109829=>"110000001",
109830=>"000000111",
109831=>"011111111",
109832=>"000100111",
109833=>"111010111",
109834=>"110110101",
109835=>"001111010",
109836=>"000111100",
109837=>"100000011",
109838=>"000100100",
109839=>"000000000",
109840=>"001010110",
109841=>"010000011",
109842=>"000100101",
109843=>"000000111",
109844=>"100000100",
109845=>"111101111",
109846=>"111011010",
109847=>"111000010",
109848=>"011000111",
109849=>"101011000",
109850=>"000011111",
109851=>"000000100",
109852=>"111010000",
109853=>"101100111",
109854=>"100101000",
109855=>"000010010",
109856=>"000000110",
109857=>"000100010",
109858=>"111001000",
109859=>"000000010",
109860=>"010110110",
109861=>"111110000",
109862=>"000110011",
109863=>"111101101",
109864=>"010011111",
109865=>"000011010",
109866=>"001000011",
109867=>"111111010",
109868=>"101111101",
109869=>"111101111",
109870=>"110000111",
109871=>"111100000",
109872=>"111000110",
109873=>"111001100",
109874=>"110111000",
109875=>"101011111",
109876=>"011000111",
109877=>"000111111",
109878=>"010000011",
109879=>"100101001",
109880=>"100011111",
109881=>"000000010",
109882=>"001000000",
109883=>"111111111",
109884=>"100110110",
109885=>"010010010",
109886=>"000000100",
109887=>"111111111",
109888=>"000000010",
109889=>"101111100",
109890=>"110000000",
109891=>"011011100",
109892=>"101101111",
109893=>"001001000",
109894=>"101000011",
109895=>"110000000",
109896=>"110101111",
109897=>"010111111",
109898=>"000100000",
109899=>"000010110",
109900=>"111111111",
109901=>"000011000",
109902=>"100110100",
109903=>"000000000",
109904=>"010011000",
109905=>"000000001",
109906=>"111011000",
109907=>"001010111",
109908=>"000000010",
109909=>"101110100",
109910=>"010001001",
109911=>"100000010",
109912=>"000001001",
109913=>"001111011",
109914=>"000011010",
109915=>"110000000",
109916=>"111111000",
109917=>"100100100",
109918=>"111101111",
109919=>"100101111",
109920=>"111101101",
109921=>"001000000",
109922=>"001101000",
109923=>"000111111",
109924=>"000011001",
109925=>"110110000",
109926=>"111111111",
109927=>"001001000",
109928=>"101111010",
109929=>"010101011",
109930=>"000010111",
109931=>"111000100",
109932=>"111110101",
109933=>"101111111",
109934=>"101100001",
109935=>"111010101",
109936=>"010011101",
109937=>"100011111",
109938=>"011000010",
109939=>"100100100",
109940=>"100111111",
109941=>"101000000",
109942=>"111010010",
109943=>"101101101",
109944=>"011000101",
109945=>"111010000",
109946=>"111000000",
109947=>"000010000",
109948=>"101110010",
109949=>"000000011",
109950=>"111011111",
109951=>"100101011",
109952=>"010000000",
109953=>"000011000",
109954=>"111000111",
109955=>"111001111",
109956=>"111111111",
109957=>"000000101",
109958=>"011011000",
109959=>"000011011",
109960=>"110110110",
109961=>"001011000",
109962=>"000000000",
109963=>"001000111",
109964=>"111100100",
109965=>"001000001",
109966=>"000101111",
109967=>"100000000",
109968=>"011011101",
109969=>"000010111",
109970=>"000000011",
109971=>"000010111",
109972=>"000100111",
109973=>"010111111",
109974=>"111111110",
109975=>"100000000",
109976=>"101001110",
109977=>"000001011",
109978=>"100010000",
109979=>"001000101",
109980=>"100000111",
109981=>"000000000",
109982=>"111000110",
109983=>"000111111",
109984=>"011011001",
109985=>"111111011",
109986=>"000000111",
109987=>"110000111",
109988=>"111010010",
109989=>"000000000",
109990=>"000001111",
109991=>"000101000",
109992=>"110000011",
109993=>"011000000",
109994=>"011010000",
109995=>"010100100",
109996=>"000010000",
109997=>"011111000",
109998=>"000100101",
109999=>"101101101",
110000=>"111011101",
110001=>"000110110",
110002=>"001001111",
110003=>"011001000",
110004=>"110110111",
110005=>"110100011",
110006=>"001001100",
110007=>"101111000",
110008=>"001011001",
110009=>"000110011",
110010=>"010010000",
110011=>"001111111",
110012=>"100101101",
110013=>"011011111",
110014=>"101011100",
110015=>"011111000",
110016=>"111111100",
110017=>"011011000",
110018=>"010010101",
110019=>"001100000",
110020=>"111101111",
110021=>"110110001",
110022=>"010010111",
110023=>"000100111",
110024=>"100111111",
110025=>"000100111",
110026=>"100111011",
110027=>"000100111",
110028=>"111100100",
110029=>"000000010",
110030=>"010111010",
110031=>"111101111",
110032=>"001010000",
110033=>"001010000",
110034=>"000000111",
110035=>"000110000",
110036=>"111000101",
110037=>"010011011",
110038=>"000011010",
110039=>"111010111",
110040=>"100101111",
110041=>"110100000",
110042=>"001000000",
110043=>"111000001",
110044=>"100111011",
110045=>"101100000",
110046=>"111101111",
110047=>"010000111",
110048=>"111000100",
110049=>"000111001",
110050=>"101000101",
110051=>"010001100",
110052=>"000000000",
110053=>"111101000",
110054=>"010111001",
110055=>"011011101",
110056=>"111100100",
110057=>"111111111",
110058=>"011011000",
110059=>"111000101",
110060=>"011001011",
110061=>"111010000",
110062=>"000000000",
110063=>"001010000",
110064=>"100100111",
110065=>"011111100",
110066=>"000010011",
110067=>"111111111",
110068=>"000101011",
110069=>"001111101",
110070=>"000000000",
110071=>"111101001",
110072=>"010111001",
110073=>"110001110",
110074=>"010010110",
110075=>"011010111",
110076=>"110111011",
110077=>"111101111",
110078=>"100111001",
110079=>"000010000",
110080=>"001000000",
110081=>"000001111",
110082=>"000110000",
110083=>"111000101",
110084=>"110111110",
110085=>"111110000",
110086=>"110000000",
110087=>"001000011",
110088=>"011011000",
110089=>"000000000",
110090=>"011011101",
110091=>"111110100",
110092=>"000001111",
110093=>"011010000",
110094=>"000011011",
110095=>"110000000",
110096=>"101000110",
110097=>"111111000",
110098=>"011101101",
110099=>"000011011",
110100=>"001000011",
110101=>"000111111",
110102=>"110000000",
110103=>"110010010",
110104=>"000000000",
110105=>"000000110",
110106=>"011010000",
110107=>"010000100",
110108=>"101100111",
110109=>"011100100",
110110=>"000000000",
110111=>"000000101",
110112=>"000000000",
110113=>"000000010",
110114=>"010101001",
110115=>"111011010",
110116=>"100100100",
110117=>"101111110",
110118=>"011011111",
110119=>"111111010",
110120=>"110110111",
110121=>"101000111",
110122=>"111111000",
110123=>"111111111",
110124=>"111011001",
110125=>"000010010",
110126=>"111110000",
110127=>"110010000",
110128=>"010000010",
110129=>"101100100",
110130=>"011000000",
110131=>"111000010",
110132=>"000010000",
110133=>"101111011",
110134=>"001011011",
110135=>"000000000",
110136=>"011000000",
110137=>"001101000",
110138=>"000000100",
110139=>"010010000",
110140=>"111011011",
110141=>"111101010",
110142=>"000111011",
110143=>"011001111",
110144=>"010101000",
110145=>"000101111",
110146=>"111001111",
110147=>"011011111",
110148=>"101000000",
110149=>"001000000",
110150=>"000000000",
110151=>"000000101",
110152=>"101100110",
110153=>"101001000",
110154=>"001000000",
110155=>"101011010",
110156=>"111010111",
110157=>"101111011",
110158=>"001001111",
110159=>"000011111",
110160=>"000111111",
110161=>"001000000",
110162=>"001101111",
110163=>"011100000",
110164=>"000101111",
110165=>"111000000",
110166=>"001001001",
110167=>"111111111",
110168=>"100110110",
110169=>"000100101",
110170=>"000110110",
110171=>"011100011",
110172=>"111111101",
110173=>"110001001",
110174=>"010111000",
110175=>"010110010",
110176=>"000110010",
110177=>"111111000",
110178=>"000010111",
110179=>"000001001",
110180=>"101101000",
110181=>"111000101",
110182=>"111111010",
110183=>"000100101",
110184=>"010000000",
110185=>"010000001",
110186=>"000000000",
110187=>"001111101",
110188=>"111110000",
110189=>"111000000",
110190=>"000000111",
110191=>"000010010",
110192=>"110111110",
110193=>"011010000",
110194=>"110110100",
110195=>"110011001",
110196=>"000000111",
110197=>"111100010",
110198=>"110100110",
110199=>"001111111",
110200=>"000010111",
110201=>"000000000",
110202=>"010000110",
110203=>"111000000",
110204=>"001000101",
110205=>"111000000",
110206=>"000001000",
110207=>"000100111",
110208=>"000000010",
110209=>"110000000",
110210=>"111111000",
110211=>"101111101",
110212=>"000000001",
110213=>"111110010",
110214=>"100110111",
110215=>"100100011",
110216=>"001101101",
110217=>"000110111",
110218=>"000111111",
110219=>"010111000",
110220=>"110111111",
110221=>"000111110",
110222=>"111101000",
110223=>"000010000",
110224=>"111101100",
110225=>"100100101",
110226=>"010100100",
110227=>"001000100",
110228=>"000110011",
110229=>"111110000",
110230=>"001000000",
110231=>"011001000",
110232=>"111101111",
110233=>"101111111",
110234=>"000001001",
110235=>"000000000",
110236=>"000000000",
110237=>"111111111",
110238=>"001000000",
110239=>"000111111",
110240=>"101100001",
110241=>"010000000",
110242=>"101101000",
110243=>"111111100",
110244=>"101000111",
110245=>"011011100",
110246=>"001101011",
110247=>"111110111",
110248=>"111111100",
110249=>"101001111",
110250=>"000000000",
110251=>"110110110",
110252=>"110101111",
110253=>"000111111",
110254=>"001001001",
110255=>"000111111",
110256=>"111100010",
110257=>"000001111",
110258=>"000000000",
110259=>"000110100",
110260=>"111100101",
110261=>"000111110",
110262=>"000101011",
110263=>"110001111",
110264=>"111110000",
110265=>"000011110",
110266=>"111111000",
110267=>"110001111",
110268=>"111111110",
110269=>"000111111",
110270=>"110111011",
110271=>"011000000",
110272=>"000000111",
110273=>"110110000",
110274=>"010000100",
110275=>"000110100",
110276=>"111000011",
110277=>"100100001",
110278=>"011000110",
110279=>"000010110",
110280=>"001111010",
110281=>"100111111",
110282=>"100101010",
110283=>"111111010",
110284=>"011001000",
110285=>"100000111",
110286=>"000000001",
110287=>"010000111",
110288=>"111101111",
110289=>"100011111",
110290=>"000011111",
110291=>"010100010",
110292=>"000010111",
110293=>"100000000",
110294=>"101100101",
110295=>"010100000",
110296=>"101100111",
110297=>"011111101",
110298=>"101110111",
110299=>"110111010",
110300=>"011000001",
110301=>"000111111",
110302=>"000101100",
110303=>"010000010",
110304=>"000010111",
110305=>"000111111",
110306=>"111111111",
110307=>"000111111",
110308=>"000010111",
110309=>"101001011",
110310=>"111011111",
110311=>"100000111",
110312=>"110011100",
110313=>"000010010",
110314=>"110100100",
110315=>"110001100",
110316=>"000110000",
110317=>"011011111",
110318=>"010000000",
110319=>"000000010",
110320=>"000000000",
110321=>"001001110",
110322=>"101000001",
110323=>"111011000",
110324=>"110000000",
110325=>"000101001",
110326=>"000010011",
110327=>"000100000",
110328=>"111000000",
110329=>"111000000",
110330=>"101101111",
110331=>"000111111",
110332=>"001011111",
110333=>"110100100",
110334=>"111111100",
110335=>"000100111",
110336=>"011011101",
110337=>"110011001",
110338=>"001000000",
110339=>"110000011",
110340=>"010100100",
110341=>"000000110",
110342=>"110110011",
110343=>"110111111",
110344=>"000001001",
110345=>"000111101",
110346=>"000100110",
110347=>"111111100",
110348=>"001111111",
110349=>"000000111",
110350=>"000000010",
110351=>"111111001",
110352=>"100111000",
110353=>"111000000",
110354=>"000101000",
110355=>"111001000",
110356=>"111111011",
110357=>"111001111",
110358=>"011111110",
110359=>"111111111",
110360=>"001001001",
110361=>"001110111",
110362=>"101001101",
110363=>"000110000",
110364=>"101000001",
110365=>"111111000",
110366=>"110111111",
110367=>"001111010",
110368=>"100110000",
110369=>"000000000",
110370=>"000000100",
110371=>"111101111",
110372=>"110001001",
110373=>"010011110",
110374=>"111001001",
110375=>"001110110",
110376=>"111110101",
110377=>"001111111",
110378=>"001101111",
110379=>"100000000",
110380=>"111000100",
110381=>"111000110",
110382=>"110000101",
110383=>"000100100",
110384=>"111000000",
110385=>"110100100",
110386=>"000000001",
110387=>"011110110",
110388=>"101110000",
110389=>"110111110",
110390=>"000011011",
110391=>"110111001",
110392=>"111111111",
110393=>"000001001",
110394=>"000000101",
110395=>"110000000",
110396=>"000100110",
110397=>"111111111",
110398=>"111000001",
110399=>"010011111",
110400=>"001000100",
110401=>"101100000",
110402=>"000000101",
110403=>"001110011",
110404=>"000001000",
110405=>"010110001",
110406=>"101011000",
110407=>"000001000",
110408=>"111000000",
110409=>"000000110",
110410=>"110001111",
110411=>"000000110",
110412=>"111001001",
110413=>"101001000",
110414=>"001001011",
110415=>"111001001",
110416=>"000010110",
110417=>"111110111",
110418=>"010101001",
110419=>"011000100",
110420=>"010000000",
110421=>"101111111",
110422=>"100011001",
110423=>"001010110",
110424=>"101001110",
110425=>"000101111",
110426=>"000101101",
110427=>"101001001",
110428=>"100000000",
110429=>"000000000",
110430=>"000110110",
110431=>"000000100",
110432=>"001000000",
110433=>"100010011",
110434=>"001000000",
110435=>"100111111",
110436=>"000000000",
110437=>"000001010",
110438=>"000111111",
110439=>"000111001",
110440=>"000100111",
110441=>"111000001",
110442=>"000000111",
110443=>"111110110",
110444=>"111010011",
110445=>"011000000",
110446=>"011000111",
110447=>"111001111",
110448=>"110100100",
110449=>"000001101",
110450=>"001111100",
110451=>"000000111",
110452=>"101001111",
110453=>"011000000",
110454=>"000001111",
110455=>"110110001",
110456=>"001010011",
110457=>"011011000",
110458=>"011000011",
110459=>"000000110",
110460=>"000110111",
110461=>"100100000",
110462=>"000001010",
110463=>"000000111",
110464=>"001000110",
110465=>"100100001",
110466=>"111000000",
110467=>"111000001",
110468=>"111101011",
110469=>"000100010",
110470=>"011011101",
110471=>"000000000",
110472=>"001001001",
110473=>"010010010",
110474=>"010000000",
110475=>"000000000",
110476=>"000110001",
110477=>"101111000",
110478=>"000110110",
110479=>"001000001",
110480=>"011101101",
110481=>"000111110",
110482=>"111000001",
110483=>"100101101",
110484=>"000110110",
110485=>"100000100",
110486=>"000110000",
110487=>"000000001",
110488=>"111111111",
110489=>"111011000",
110490=>"001111111",
110491=>"000010000",
110492=>"110000101",
110493=>"010110110",
110494=>"000001111",
110495=>"101001001",
110496=>"000000111",
110497=>"010111110",
110498=>"000000000",
110499=>"001000100",
110500=>"111000000",
110501=>"101001011",
110502=>"000000000",
110503=>"000001111",
110504=>"111111010",
110505=>"010000001",
110506=>"001000000",
110507=>"001000000",
110508=>"011000000",
110509=>"101000000",
110510=>"100111011",
110511=>"000110000",
110512=>"100000110",
110513=>"111011101",
110514=>"111010110",
110515=>"000000100",
110516=>"010011010",
110517=>"110100110",
110518=>"111101000",
110519=>"000110111",
110520=>"101011001",
110521=>"000000100",
110522=>"000101001",
110523=>"110011100",
110524=>"111111111",
110525=>"111111111",
110526=>"000100100",
110527=>"011101111",
110528=>"000110000",
110529=>"001000000",
110530=>"001111011",
110531=>"001001111",
110532=>"000000111",
110533=>"101100001",
110534=>"110110101",
110535=>"010111111",
110536=>"010000101",
110537=>"111001001",
110538=>"000000001",
110539=>"111111110",
110540=>"000101110",
110541=>"100000011",
110542=>"011001000",
110543=>"001000111",
110544=>"010001000",
110545=>"000000001",
110546=>"000000000",
110547=>"111100100",
110548=>"111111111",
110549=>"101001011",
110550=>"001001000",
110551=>"000000000",
110552=>"001001011",
110553=>"000000001",
110554=>"000000011",
110555=>"011000111",
110556=>"110111001",
110557=>"110100110",
110558=>"111001001",
110559=>"110111111",
110560=>"111000001",
110561=>"011110110",
110562=>"000110110",
110563=>"000001001",
110564=>"000000000",
110565=>"101000001",
110566=>"100000000",
110567=>"011111000",
110568=>"000101101",
110569=>"110001000",
110570=>"011111110",
110571=>"111000000",
110572=>"000000001",
110573=>"111111111",
110574=>"111001000",
110575=>"111000001",
110576=>"110101001",
110577=>"011110010",
110578=>"111000000",
110579=>"101001101",
110580=>"110110001",
110581=>"000001111",
110582=>"100000000",
110583=>"001001011",
110584=>"000010111",
110585=>"101111011",
110586=>"111001001",
110587=>"101110000",
110588=>"111111001",
110589=>"000010000",
110590=>"010010011",
110591=>"111001001",
110592=>"111000101",
110593=>"100111111",
110594=>"000000111",
110595=>"000011010",
110596=>"001001111",
110597=>"101100010",
110598=>"000100111",
110599=>"111010001",
110600=>"100010000",
110601=>"000111111",
110602=>"000011011",
110603=>"010111101",
110604=>"111000000",
110605=>"000101111",
110606=>"100111111",
110607=>"001010010",
110608=>"010110000",
110609=>"000000000",
110610=>"111110000",
110611=>"000000000",
110612=>"101011000",
110613=>"110000000",
110614=>"101000010",
110615=>"010000001",
110616=>"110111000",
110617=>"000100000",
110618=>"000000001",
110619=>"000111010",
110620=>"001101000",
110621=>"111111000",
110622=>"111000110",
110623=>"000000111",
110624=>"000010000",
110625=>"000011111",
110626=>"111010001",
110627=>"111111001",
110628=>"100001111",
110629=>"001001000",
110630=>"000101010",
110631=>"101001111",
110632=>"000000010",
110633=>"010100101",
110634=>"111000111",
110635=>"000101011",
110636=>"111101001",
110637=>"111111000",
110638=>"101111111",
110639=>"011011111",
110640=>"111001101",
110641=>"001101011",
110642=>"111111111",
110643=>"111010000",
110644=>"011001111",
110645=>"111000000",
110646=>"000000000",
110647=>"001111111",
110648=>"110101000",
110649=>"001000111",
110650=>"000000110",
110651=>"101000001",
110652=>"101001001",
110653=>"000101101",
110654=>"000000110",
110655=>"101100110",
110656=>"111010000",
110657=>"010000000",
110658=>"100000011",
110659=>"101011101",
110660=>"101000000",
110661=>"010000001",
110662=>"000100111",
110663=>"111111111",
110664=>"111011001",
110665=>"010111010",
110666=>"111101111",
110667=>"000000111",
110668=>"111010111",
110669=>"011110111",
110670=>"100101101",
110671=>"111111110",
110672=>"000001111",
110673=>"000010000",
110674=>"111111111",
110675=>"100110000",
110676=>"000100010",
110677=>"110111111",
110678=>"000000111",
110679=>"110111010",
110680=>"010000000",
110681=>"000001000",
110682=>"001011111",
110683=>"100100101",
110684=>"111010000",
110685=>"000001000",
110686=>"111111000",
110687=>"011111111",
110688=>"000000000",
110689=>"111111111",
110690=>"100000000",
110691=>"100100101",
110692=>"111010000",
110693=>"000000100",
110694=>"100111111",
110695=>"001111111",
110696=>"101000010",
110697=>"110000000",
110698=>"111111100",
110699=>"110000000",
110700=>"101000110",
110701=>"111111000",
110702=>"111000001",
110703=>"001111111",
110704=>"001111111",
110705=>"000101110",
110706=>"110000000",
110707=>"010000001",
110708=>"111000000",
110709=>"001000000",
110710=>"011001111",
110711=>"000000111",
110712=>"110111010",
110713=>"000000111",
110714=>"111110101",
110715=>"110111000",
110716=>"011110100",
110717=>"111000010",
110718=>"111111111",
110719=>"000101111",
110720=>"111000000",
110721=>"000111000",
110722=>"111111000",
110723=>"111010011",
110724=>"001110111",
110725=>"000100000",
110726=>"000100000",
110727=>"110100000",
110728=>"100011111",
110729=>"000110000",
110730=>"010010000",
110731=>"000111101",
110732=>"000000000",
110733=>"000111011",
110734=>"111000000",
110735=>"000010011",
110736=>"101111001",
110737=>"111101010",
110738=>"000001101",
110739=>"010111000",
110740=>"111111010",
110741=>"100111000",
110742=>"010001101",
110743=>"010100100",
110744=>"010011010",
110745=>"111010011",
110746=>"000001000",
110747=>"100111110",
110748=>"010011001",
110749=>"111011000",
110750=>"010111111",
110751=>"000000011",
110752=>"011101111",
110753=>"110000000",
110754=>"001111101",
110755=>"000000000",
110756=>"111001001",
110757=>"000000001",
110758=>"111011001",
110759=>"100011001",
110760=>"111111111",
110761=>"111011001",
110762=>"111000101",
110763=>"000000111",
110764=>"010010111",
110765=>"000010111",
110766=>"000001011",
110767=>"000000011",
110768=>"101100000",
110769=>"011000000",
110770=>"110000000",
110771=>"001000110",
110772=>"111111010",
110773=>"010011111",
110774=>"111000000",
110775=>"110000000",
110776=>"001000100",
110777=>"001011000",
110778=>"111111111",
110779=>"000000100",
110780=>"011001100",
110781=>"111000111",
110782=>"011001001",
110783=>"010000111",
110784=>"000100010",
110785=>"000010110",
110786=>"111011000",
110787=>"100100110",
110788=>"110000111",
110789=>"110110011",
110790=>"011000000",
110791=>"101111100",
110792=>"111111101",
110793=>"001000000",
110794=>"000000000",
110795=>"110000000",
110796=>"000010010",
110797=>"110010001",
110798=>"000001110",
110799=>"110011000",
110800=>"111111010",
110801=>"011000111",
110802=>"010111111",
110803=>"111111111",
110804=>"100111111",
110805=>"000100000",
110806=>"001111111",
110807=>"010111111",
110808=>"000000000",
110809=>"001000000",
110810=>"101100100",
110811=>"110110110",
110812=>"011000100",
110813=>"000110111",
110814=>"000000000",
110815=>"111001100",
110816=>"000100110",
110817=>"110111111",
110818=>"111000000",
110819=>"000100111",
110820=>"000000011",
110821=>"001111010",
110822=>"111111110",
110823=>"001000100",
110824=>"111101101",
110825=>"010111000",
110826=>"000110110",
110827=>"111000111",
110828=>"110111111",
110829=>"111011001",
110830=>"000000010",
110831=>"111000000",
110832=>"000001000",
110833=>"111111110",
110834=>"001001101",
110835=>"110111000",
110836=>"101001011",
110837=>"000111111",
110838=>"000000111",
110839=>"111111000",
110840=>"111011000",
110841=>"000101010",
110842=>"000010001",
110843=>"001011000",
110844=>"010000000",
110845=>"000010000",
110846=>"110100010",
110847=>"111111111",
110848=>"000000001",
110849=>"110001111",
110850=>"000000110",
110851=>"010101001",
110852=>"100100110",
110853=>"001000110",
110854=>"110000111",
110855=>"111111111",
110856=>"001001111",
110857=>"111000011",
110858=>"001111110",
110859=>"000000100",
110860=>"000000000",
110861=>"000110110",
110862=>"000000011",
110863=>"111111000",
110864=>"111111110",
110865=>"110111111",
110866=>"101000000",
110867=>"011111111",
110868=>"111111000",
110869=>"001001011",
110870=>"010100000",
110871=>"010011111",
110872=>"000000011",
110873=>"011001000",
110874=>"000100000",
110875=>"000000000",
110876=>"000100000",
110877=>"100100111",
110878=>"000001111",
110879=>"010101000",
110880=>"011111000",
110881=>"000010000",
110882=>"011111111",
110883=>"010011111",
110884=>"000110010",
110885=>"101001110",
110886=>"000110010",
110887=>"100111110",
110888=>"011111010",
110889=>"000001000",
110890=>"000000000",
110891=>"000000000",
110892=>"010011011",
110893=>"101101000",
110894=>"111111111",
110895=>"001000000",
110896=>"000111000",
110897=>"111011111",
110898=>"110111000",
110899=>"000011111",
110900=>"111111110",
110901=>"111101101",
110902=>"110110010",
110903=>"001000111",
110904=>"000001000",
110905=>"001000000",
110906=>"100110111",
110907=>"010110000",
110908=>"010011001",
110909=>"010000111",
110910=>"010000111",
110911=>"110000000",
110912=>"111011010",
110913=>"000011111",
110914=>"010000111",
110915=>"101101111",
110916=>"111110111",
110917=>"111001000",
110918=>"001000000",
110919=>"111000000",
110920=>"010111111",
110921=>"010110110",
110922=>"111111001",
110923=>"111111111",
110924=>"000000000",
110925=>"011011110",
110926=>"001001001",
110927=>"000000000",
110928=>"010000000",
110929=>"110111110",
110930=>"111000000",
110931=>"001001000",
110932=>"100000111",
110933=>"111110110",
110934=>"010011001",
110935=>"101111000",
110936=>"000000000",
110937=>"000000000",
110938=>"000000100",
110939=>"011011011",
110940=>"000000000",
110941=>"111110000",
110942=>"000000000",
110943=>"001100100",
110944=>"000000000",
110945=>"010110100",
110946=>"000110111",
110947=>"111101000",
110948=>"001111101",
110949=>"100000101",
110950=>"110110110",
110951=>"001000000",
110952=>"110001000",
110953=>"001001111",
110954=>"100000000",
110955=>"101000010",
110956=>"000000000",
110957=>"101111001",
110958=>"101000111",
110959=>"100111111",
110960=>"110110110",
110961=>"000000000",
110962=>"000000100",
110963=>"000000111",
110964=>"010110111",
110965=>"111000111",
110966=>"100000000",
110967=>"001101111",
110968=>"010000110",
110969=>"000000000",
110970=>"000111111",
110971=>"111111101",
110972=>"011001010",
110973=>"100000000",
110974=>"111111011",
110975=>"100111001",
110976=>"000000000",
110977=>"111000000",
110978=>"000000000",
110979=>"000001110",
110980=>"001000111",
110981=>"000000110",
110982=>"100110110",
110983=>"000101001",
110984=>"011011111",
110985=>"000010111",
110986=>"111111111",
110987=>"001001010",
110988=>"010000000",
110989=>"110000111",
110990=>"001001000",
110991=>"000000110",
110992=>"111101101",
110993=>"000000111",
110994=>"111111111",
110995=>"001000110",
110996=>"100010000",
110997=>"101000000",
110998=>"111001001",
110999=>"110110000",
111000=>"011101110",
111001=>"110100010",
111002=>"000000010",
111003=>"111000011",
111004=>"111100000",
111005=>"111111111",
111006=>"011111111",
111007=>"101000001",
111008=>"000000000",
111009=>"111100000",
111010=>"000000100",
111011=>"000001110",
111012=>"101001111",
111013=>"110000000",
111014=>"011111011",
111015=>"100001111",
111016=>"111001000",
111017=>"000001101",
111018=>"000000000",
111019=>"101001000",
111020=>"011000111",
111021=>"000000000",
111022=>"101101100",
111023=>"011000110",
111024=>"000000000",
111025=>"000100101",
111026=>"010110000",
111027=>"010000100",
111028=>"111111111",
111029=>"000101111",
111030=>"001000000",
111031=>"111101111",
111032=>"101100100",
111033=>"111111100",
111034=>"001111101",
111035=>"011111111",
111036=>"000110010",
111037=>"010010000",
111038=>"110000001",
111039=>"001000000",
111040=>"111101100",
111041=>"001000111",
111042=>"000111101",
111043=>"101100110",
111044=>"001000000",
111045=>"111101000",
111046=>"010011000",
111047=>"111111110",
111048=>"110000000",
111049=>"000101111",
111050=>"001000000",
111051=>"111111111",
111052=>"111000101",
111053=>"100100001",
111054=>"100101101",
111055=>"101111111",
111056=>"000010110",
111057=>"010010000",
111058=>"111111000",
111059=>"111101101",
111060=>"000000100",
111061=>"111011111",
111062=>"101000000",
111063=>"100000100",
111064=>"000000001",
111065=>"100111011",
111066=>"100000000",
111067=>"111111110",
111068=>"000000011",
111069=>"110111110",
111070=>"001000000",
111071=>"001110100",
111072=>"000000000",
111073=>"000010111",
111074=>"111111000",
111075=>"011111111",
111076=>"111011111",
111077=>"111101111",
111078=>"000000000",
111079=>"011011011",
111080=>"111111100",
111081=>"111011110",
111082=>"010111111",
111083=>"101111010",
111084=>"111111111",
111085=>"001000000",
111086=>"010010000",
111087=>"111111111",
111088=>"000000000",
111089=>"011001000",
111090=>"101000000",
111091=>"110000000",
111092=>"001010110",
111093=>"000100110",
111094=>"111101000",
111095=>"000011111",
111096=>"101111011",
111097=>"111111111",
111098=>"000000000",
111099=>"101000000",
111100=>"010111011",
111101=>"000111001",
111102=>"001011011",
111103=>"010010011",
111104=>"000100100",
111105=>"000000000",
111106=>"000000001",
111107=>"000011101",
111108=>"110100000",
111109=>"011110000",
111110=>"111010000",
111111=>"100100111",
111112=>"010011001",
111113=>"111111000",
111114=>"000000001",
111115=>"110111111",
111116=>"000000100",
111117=>"111111000",
111118=>"100100000",
111119=>"111111111",
111120=>"001000100",
111121=>"101000101",
111122=>"001000001",
111123=>"111111010",
111124=>"111101111",
111125=>"001000000",
111126=>"000011111",
111127=>"000001000",
111128=>"010101100",
111129=>"100100000",
111130=>"110011000",
111131=>"000000000",
111132=>"100000000",
111133=>"010001000",
111134=>"111010000",
111135=>"010010010",
111136=>"000111001",
111137=>"111101111",
111138=>"101101111",
111139=>"101100110",
111140=>"010100000",
111141=>"000011011",
111142=>"111110000",
111143=>"111111000",
111144=>"000000010",
111145=>"000100111",
111146=>"111111000",
111147=>"100011111",
111148=>"111111100",
111149=>"000100101",
111150=>"100000010",
111151=>"010000111",
111152=>"111000000",
111153=>"011011000",
111154=>"111101101",
111155=>"111101111",
111156=>"100000000",
111157=>"111101111",
111158=>"000000000",
111159=>"111111001",
111160=>"101111111",
111161=>"111101000",
111162=>"101110011",
111163=>"110000011",
111164=>"111000000",
111165=>"110111010",
111166=>"000100000",
111167=>"001011010",
111168=>"010101111",
111169=>"000011001",
111170=>"000000101",
111171=>"110011001",
111172=>"111111011",
111173=>"010111111",
111174=>"010011000",
111175=>"111111001",
111176=>"011011110",
111177=>"000000111",
111178=>"101100110",
111179=>"111111111",
111180=>"101111000",
111181=>"011111101",
111182=>"110110000",
111183=>"000000101",
111184=>"100001001",
111185=>"000000111",
111186=>"010010000",
111187=>"011000000",
111188=>"000000000",
111189=>"000100000",
111190=>"011011000",
111191=>"000010000",
111192=>"111111110",
111193=>"000001001",
111194=>"110011011",
111195=>"010110001",
111196=>"000000011",
111197=>"001001111",
111198=>"000000000",
111199=>"111110000",
111200=>"010011010",
111201=>"101000100",
111202=>"000100100",
111203=>"111111000",
111204=>"010010010",
111205=>"000100100",
111206=>"000000111",
111207=>"010000000",
111208=>"100111111",
111209=>"111100011",
111210=>"000000010",
111211=>"111111101",
111212=>"101000000",
111213=>"111000111",
111214=>"000000111",
111215=>"111000111",
111216=>"101101000",
111217=>"000000111",
111218=>"000000000",
111219=>"111111000",
111220=>"000011111",
111221=>"000100100",
111222=>"100000111",
111223=>"111111111",
111224=>"111001000",
111225=>"000011010",
111226=>"011111110",
111227=>"000000111",
111228=>"000000110",
111229=>"110100000",
111230=>"000000111",
111231=>"010110100",
111232=>"101100100",
111233=>"000010011",
111234=>"111000000",
111235=>"111111001",
111236=>"111110010",
111237=>"101101111",
111238=>"010100110",
111239=>"110100100",
111240=>"111100100",
111241=>"000000000",
111242=>"000111110",
111243=>"111000101",
111244=>"000011111",
111245=>"010101111",
111246=>"000100111",
111247=>"111001110",
111248=>"100100111",
111249=>"101111011",
111250=>"001000010",
111251=>"111100000",
111252=>"110000000",
111253=>"001001101",
111254=>"111111101",
111255=>"111101111",
111256=>"001111010",
111257=>"000010011",
111258=>"111111000",
111259=>"100101100",
111260=>"011111111",
111261=>"011111111",
111262=>"110101101",
111263=>"110111000",
111264=>"011010001",
111265=>"000001100",
111266=>"111101111",
111267=>"011001000",
111268=>"110100100",
111269=>"011010000",
111270=>"111110000",
111271=>"001000100",
111272=>"111011100",
111273=>"000011111",
111274=>"101111111",
111275=>"101111000",
111276=>"000000101",
111277=>"011000001",
111278=>"100111001",
111279=>"111000111",
111280=>"100100111",
111281=>"110101100",
111282=>"000000111",
111283=>"000000100",
111284=>"111110111",
111285=>"000010000",
111286=>"110110110",
111287=>"000000101",
111288=>"111111001",
111289=>"001000001",
111290=>"000000100",
111291=>"000100111",
111292=>"110000011",
111293=>"000111111",
111294=>"110110000",
111295=>"101110111",
111296=>"000000101",
111297=>"000000000",
111298=>"101011111",
111299=>"111100100",
111300=>"101100011",
111301=>"000010111",
111302=>"111111000",
111303=>"000000000",
111304=>"000010000",
111305=>"000000000",
111306=>"100000100",
111307=>"010001111",
111308=>"000000000",
111309=>"100100000",
111310=>"100111010",
111311=>"000111010",
111312=>"111011000",
111313=>"111111110",
111314=>"110000001",
111315=>"011101010",
111316=>"100000001",
111317=>"000000010",
111318=>"100111110",
111319=>"000000011",
111320=>"000000110",
111321=>"101100100",
111322=>"110011100",
111323=>"101100101",
111324=>"000100111",
111325=>"100111111",
111326=>"111111000",
111327=>"011111000",
111328=>"000001010",
111329=>"000000101",
111330=>"000010000",
111331=>"010000000",
111332=>"100111001",
111333=>"000100111",
111334=>"011111111",
111335=>"011111100",
111336=>"111101000",
111337=>"101101010",
111338=>"001100111",
111339=>"101101101",
111340=>"000000100",
111341=>"010111000",
111342=>"011010101",
111343=>"000000000",
111344=>"111111010",
111345=>"000011111",
111346=>"111011000",
111347=>"011011100",
111348=>"111110000",
111349=>"111111010",
111350=>"101100000",
111351=>"110101011",
111352=>"000000111",
111353=>"000001111",
111354=>"110100111",
111355=>"000000000",
111356=>"010111000",
111357=>"000000000",
111358=>"110100110",
111359=>"000000000",
111360=>"001001010",
111361=>"000101110",
111362=>"000000001",
111363=>"000000000",
111364=>"101111111",
111365=>"000001001",
111366=>"011111111",
111367=>"111111111",
111368=>"000000001",
111369=>"010110101",
111370=>"001011011",
111371=>"001000111",
111372=>"000000000",
111373=>"000000000",
111374=>"000011110",
111375=>"101111001",
111376=>"110100111",
111377=>"000010011",
111378=>"000001001",
111379=>"101101100",
111380=>"101000100",
111381=>"000111000",
111382=>"111111110",
111383=>"111111000",
111384=>"101001000",
111385=>"111001001",
111386=>"000000000",
111387=>"000000101",
111388=>"101101111",
111389=>"101000001",
111390=>"010010011",
111391=>"010111110",
111392=>"111101101",
111393=>"111111111",
111394=>"000010111",
111395=>"111110000",
111396=>"010001101",
111397=>"100111010",
111398=>"110011001",
111399=>"111110000",
111400=>"000000000",
111401=>"000001010",
111402=>"111111111",
111403=>"010001101",
111404=>"000100100",
111405=>"101010000",
111406=>"111101111",
111407=>"011110111",
111408=>"111000000",
111409=>"111110110",
111410=>"001101000",
111411=>"100000000",
111412=>"101000111",
111413=>"111111111",
111414=>"110111111",
111415=>"000000000",
111416=>"111000000",
111417=>"000000010",
111418=>"000000000",
111419=>"101110111",
111420=>"111001000",
111421=>"111111000",
111422=>"001000101",
111423=>"111111011",
111424=>"001101111",
111425=>"010101110",
111426=>"000000000",
111427=>"011011100",
111428=>"111010111",
111429=>"101000000",
111430=>"110011001",
111431=>"101010111",
111432=>"000011100",
111433=>"000110101",
111434=>"100000000",
111435=>"111110000",
111436=>"001000110",
111437=>"000100011",
111438=>"101001010",
111439=>"001101100",
111440=>"001110111",
111441=>"111111000",
111442=>"010110011",
111443=>"011000000",
111444=>"000000000",
111445=>"111111100",
111446=>"101001111",
111447=>"000010100",
111448=>"000000011",
111449=>"001001110",
111450=>"000011011",
111451=>"001100100",
111452=>"111110000",
111453=>"000000000",
111454=>"111111111",
111455=>"110000000",
111456=>"111111111",
111457=>"011001000",
111458=>"000000101",
111459=>"100010010",
111460=>"000001100",
111461=>"000000000",
111462=>"000000000",
111463=>"011111111",
111464=>"101010111",
111465=>"101001011",
111466=>"000001111",
111467=>"100111000",
111468=>"001101100",
111469=>"010111111",
111470=>"000011000",
111471=>"000000110",
111472=>"110011011",
111473=>"000000111",
111474=>"011011110",
111475=>"100111000",
111476=>"111111111",
111477=>"000000000",
111478=>"000010101",
111479=>"000010111",
111480=>"001010111",
111481=>"000111111",
111482=>"001111000",
111483=>"101101100",
111484=>"111100000",
111485=>"110100001",
111486=>"111111111",
111487=>"101000000",
111488=>"110001000",
111489=>"100100000",
111490=>"111111110",
111491=>"000100101",
111492=>"000101111",
111493=>"000000000",
111494=>"110110111",
111495=>"111110100",
111496=>"001111111",
111497=>"110100111",
111498=>"111110000",
111499=>"111111111",
111500=>"010010000",
111501=>"001000001",
111502=>"111100011",
111503=>"000001001",
111504=>"111111001",
111505=>"000000111",
111506=>"110101000",
111507=>"000000001",
111508=>"000000100",
111509=>"000000111",
111510=>"000010010",
111511=>"000001011",
111512=>"011011001",
111513=>"001000001",
111514=>"111111010",
111515=>"100100001",
111516=>"000000100",
111517=>"001000111",
111518=>"111000000",
111519=>"011111101",
111520=>"101111100",
111521=>"100101111",
111522=>"001000100",
111523=>"000010001",
111524=>"010000000",
111525=>"101001000",
111526=>"000110000",
111527=>"001000100",
111528=>"111111000",
111529=>"001001000",
111530=>"000110110",
111531=>"000000000",
111532=>"000000001",
111533=>"000000100",
111534=>"000101011",
111535=>"000111110",
111536=>"000000010",
111537=>"100000001",
111538=>"111000000",
111539=>"000100110",
111540=>"001011111",
111541=>"101011101",
111542=>"011101111",
111543=>"001000101",
111544=>"010100000",
111545=>"011011111",
111546=>"111111000",
111547=>"010010101",
111548=>"010000000",
111549=>"111010010",
111550=>"011011111",
111551=>"000000101",
111552=>"000010000",
111553=>"000011001",
111554=>"101110000",
111555=>"001001111",
111556=>"011111000",
111557=>"001000100",
111558=>"000000010",
111559=>"110111011",
111560=>"100101111",
111561=>"010111001",
111562=>"111111111",
111563=>"101101000",
111564=>"000000100",
111565=>"101111101",
111566=>"101001101",
111567=>"111111101",
111568=>"001000111",
111569=>"001011000",
111570=>"001101000",
111571=>"000100101",
111572=>"010011000",
111573=>"110100110",
111574=>"000000010",
111575=>"000100100",
111576=>"111110110",
111577=>"111001100",
111578=>"111101101",
111579=>"111010000",
111580=>"110111101",
111581=>"000001111",
111582=>"000101101",
111583=>"110000000",
111584=>"000110101",
111585=>"000000110",
111586=>"000000111",
111587=>"111111011",
111588=>"000010111",
111589=>"000000101",
111590=>"101001110",
111591=>"011111100",
111592=>"101101000",
111593=>"011000000",
111594=>"000110110",
111595=>"110111010",
111596=>"100000111",
111597=>"100101001",
111598=>"100000000",
111599=>"111001000",
111600=>"110101010",
111601=>"100101001",
111602=>"010000000",
111603=>"100101111",
111604=>"100100100",
111605=>"000110010",
111606=>"111111000",
111607=>"001101111",
111608=>"111111000",
111609=>"010000000",
111610=>"110100111",
111611=>"101100000",
111612=>"111110000",
111613=>"100110011",
111614=>"001111101",
111615=>"001000111",
111616=>"111110101",
111617=>"000000000",
111618=>"100000111",
111619=>"010000000",
111620=>"100100110",
111621=>"001000111",
111622=>"001111001",
111623=>"000110111",
111624=>"111001000",
111625=>"110100111",
111626=>"110000000",
111627=>"101100000",
111628=>"111100111",
111629=>"000000100",
111630=>"011110100",
111631=>"111111000",
111632=>"000000001",
111633=>"100100000",
111634=>"000010111",
111635=>"000110000",
111636=>"110110100",
111637=>"111101111",
111638=>"000001111",
111639=>"011111111",
111640=>"110000000",
111641=>"111111101",
111642=>"000101100",
111643=>"100100111",
111644=>"000100110",
111645=>"001010010",
111646=>"101111000",
111647=>"111000000",
111648=>"000111101",
111649=>"010000001",
111650=>"001000010",
111651=>"010010010",
111652=>"000100011",
111653=>"010010010",
111654=>"011011000",
111655=>"000000000",
111656=>"111100110",
111657=>"111101111",
111658=>"000000110",
111659=>"100000100",
111660=>"100100110",
111661=>"110010011",
111662=>"010000000",
111663=>"001011010",
111664=>"111111000",
111665=>"110110111",
111666=>"101111111",
111667=>"000110101",
111668=>"111010000",
111669=>"000000111",
111670=>"001000000",
111671=>"010111000",
111672=>"111001000",
111673=>"010111001",
111674=>"101101111",
111675=>"101000110",
111676=>"001111001",
111677=>"111111000",
111678=>"000000000",
111679=>"111101001",
111680=>"000100100",
111681=>"000000101",
111682=>"111111000",
111683=>"000110000",
111684=>"101111111",
111685=>"111101011",
111686=>"001100100",
111687=>"001100101",
111688=>"000100101",
111689=>"010111010",
111690=>"000000111",
111691=>"100001001",
111692=>"001111101",
111693=>"110110110",
111694=>"011001111",
111695=>"101000111",
111696=>"000000100",
111697=>"101111100",
111698=>"100100110",
111699=>"001100010",
111700=>"000000110",
111701=>"110110100",
111702=>"011011000",
111703=>"110010000",
111704=>"000000101",
111705=>"100000101",
111706=>"100000010",
111707=>"010000001",
111708=>"010111000",
111709=>"001001000",
111710=>"010010010",
111711=>"010001011",
111712=>"100100111",
111713=>"001010000",
111714=>"000000111",
111715=>"000110100",
111716=>"111100000",
111717=>"100100001",
111718=>"110111110",
111719=>"110111000",
111720=>"010010110",
111721=>"100101111",
111722=>"010111011",
111723=>"110110011",
111724=>"111111111",
111725=>"100101111",
111726=>"000100110",
111727=>"001101111",
111728=>"010100000",
111729=>"110001001",
111730=>"110000000",
111731=>"001111000",
111732=>"100111011",
111733=>"001100111",
111734=>"110001111",
111735=>"101000101",
111736=>"000000110",
111737=>"000000010",
111738=>"001111110",
111739=>"111101011",
111740=>"110110010",
111741=>"100000000",
111742=>"110010111",
111743=>"000010000",
111744=>"010000000",
111745=>"101101010",
111746=>"000000000",
111747=>"001000110",
111748=>"000111111",
111749=>"010010000",
111750=>"110100110",
111751=>"011011000",
111752=>"111011000",
111753=>"110010010",
111754=>"001011010",
111755=>"000100101",
111756=>"000000101",
111757=>"000000001",
111758=>"011111000",
111759=>"000000100",
111760=>"011011011",
111761=>"000010010",
111762=>"111000001",
111763=>"101101111",
111764=>"010010111",
111765=>"000000000",
111766=>"010010000",
111767=>"111100100",
111768=>"000000000",
111769=>"010000110",
111770=>"111011010",
111771=>"101000000",
111772=>"010000111",
111773=>"101000111",
111774=>"111010000",
111775=>"110000111",
111776=>"101111001",
111777=>"001001111",
111778=>"111111000",
111779=>"111111011",
111780=>"000000000",
111781=>"100100100",
111782=>"001101100",
111783=>"001001001",
111784=>"010101111",
111785=>"000000010",
111786=>"111101100",
111787=>"100100111",
111788=>"000001000",
111789=>"000010100",
111790=>"111011001",
111791=>"100111111",
111792=>"111000101",
111793=>"100000001",
111794=>"111111101",
111795=>"101110100",
111796=>"001011001",
111797=>"111111000",
111798=>"001000100",
111799=>"111110010",
111800=>"001011000",
111801=>"101100000",
111802=>"010111111",
111803=>"000011111",
111804=>"101101110",
111805=>"101111111",
111806=>"001000100",
111807=>"001100111",
111808=>"010010000",
111809=>"000000111",
111810=>"000111001",
111811=>"100100100",
111812=>"010011000",
111813=>"110100100",
111814=>"010000000",
111815=>"000000100",
111816=>"000000001",
111817=>"101001111",
111818=>"111011010",
111819=>"111100000",
111820=>"111011111",
111821=>"101011001",
111822=>"000000000",
111823=>"000001000",
111824=>"000000100",
111825=>"111111111",
111826=>"111111111",
111827=>"111111100",
111828=>"100000000",
111829=>"000000000",
111830=>"000100000",
111831=>"001111111",
111832=>"010111011",
111833=>"000111011",
111834=>"101101110",
111835=>"100000111",
111836=>"000100000",
111837=>"000000100",
111838=>"000111100",
111839=>"010110000",
111840=>"010010110",
111841=>"000000111",
111842=>"001101111",
111843=>"111000011",
111844=>"000000100",
111845=>"101101110",
111846=>"000000101",
111847=>"010110110",
111848=>"000000101",
111849=>"010111001",
111850=>"011010010",
111851=>"111101101",
111852=>"000000111",
111853=>"000000111",
111854=>"000000000",
111855=>"000000101",
111856=>"001000000",
111857=>"011000001",
111858=>"000000111",
111859=>"000100100",
111860=>"010001001",
111861=>"000010110",
111862=>"000000000",
111863=>"100000101",
111864=>"101000011",
111865=>"000001010",
111866=>"111101111",
111867=>"100110000",
111868=>"111111000",
111869=>"011111011",
111870=>"011011011",
111871=>"000000000",
111872=>"011010011",
111873=>"100100000",
111874=>"101000111",
111875=>"000001111",
111876=>"101001000",
111877=>"000001010",
111878=>"111101111",
111879=>"111111100",
111880=>"010110110",
111881=>"111110110",
111882=>"000100110",
111883=>"000100010",
111884=>"000000111",
111885=>"010010010",
111886=>"100011011",
111887=>"101000000",
111888=>"101100110",
111889=>"111111111",
111890=>"101010101",
111891=>"111101000",
111892=>"111111111",
111893=>"010111000",
111894=>"101101101",
111895=>"111011001",
111896=>"000000010",
111897=>"100100110",
111898=>"000011001",
111899=>"010011011",
111900=>"101001100",
111901=>"111010101",
111902=>"010001000",
111903=>"000010111",
111904=>"000110010",
111905=>"000101010",
111906=>"010111000",
111907=>"101100101",
111908=>"010001011",
111909=>"010000100",
111910=>"010110010",
111911=>"011011001",
111912=>"010111010",
111913=>"101100010",
111914=>"001000000",
111915=>"111100000",
111916=>"110100111",
111917=>"000111111",
111918=>"011010000",
111919=>"000101001",
111920=>"110011110",
111921=>"000001001",
111922=>"111111100",
111923=>"110011111",
111924=>"100000101",
111925=>"100000000",
111926=>"011011000",
111927=>"010000000",
111928=>"011010010",
111929=>"101000000",
111930=>"000111010",
111931=>"000001101",
111932=>"011000110",
111933=>"111111000",
111934=>"000000010",
111935=>"001110110",
111936=>"111111100",
111937=>"001101110",
111938=>"111010110",
111939=>"001000000",
111940=>"111101101",
111941=>"001111100",
111942=>"111000101",
111943=>"100000000",
111944=>"000110111",
111945=>"010010000",
111946=>"110000101",
111947=>"110100101",
111948=>"111111010",
111949=>"010001010",
111950=>"000100111",
111951=>"001101111",
111952=>"101111000",
111953=>"010001000",
111954=>"010000100",
111955=>"011001101",
111956=>"101101100",
111957=>"000000111",
111958=>"011001010",
111959=>"100000100",
111960=>"111111110",
111961=>"000100110",
111962=>"001001000",
111963=>"110100011",
111964=>"000000000",
111965=>"000000000",
111966=>"111001111",
111967=>"000000001",
111968=>"101100000",
111969=>"000000001",
111970=>"000000000",
111971=>"101110000",
111972=>"000000111",
111973=>"000100010",
111974=>"011001001",
111975=>"010010110",
111976=>"000001101",
111977=>"111111000",
111978=>"000000000",
111979=>"111000000",
111980=>"010111110",
111981=>"101111010",
111982=>"111100100",
111983=>"000000111",
111984=>"000001000",
111985=>"000101111",
111986=>"011110100",
111987=>"111000000",
111988=>"000000000",
111989=>"011000100",
111990=>"101110010",
111991=>"101000000",
111992=>"001010111",
111993=>"011100000",
111994=>"101101101",
111995=>"000011010",
111996=>"100100001",
111997=>"110000000",
111998=>"111001001",
111999=>"000010000",
112000=>"111101100",
112001=>"100101101",
112002=>"111000000",
112003=>"101100010",
112004=>"011011111",
112005=>"111001001",
112006=>"100000001",
112007=>"011100100",
112008=>"001011001",
112009=>"111001000",
112010=>"111100000",
112011=>"010000100",
112012=>"110110011",
112013=>"111111010",
112014=>"110000111",
112015=>"010000000",
112016=>"011011010",
112017=>"011001000",
112018=>"111110001",
112019=>"010000000",
112020=>"100010000",
112021=>"000000010",
112022=>"101100101",
112023=>"000001111",
112024=>"110001010",
112025=>"011000000",
112026=>"111111001",
112027=>"100000010",
112028=>"111001000",
112029=>"111001011",
112030=>"010111110",
112031=>"101100101",
112032=>"100110111",
112033=>"000000000",
112034=>"011000000",
112035=>"011000000",
112036=>"010001011",
112037=>"011011001",
112038=>"111111100",
112039=>"111100101",
112040=>"100101101",
112041=>"101100000",
112042=>"000010000",
112043=>"001101000",
112044=>"101100110",
112045=>"010010010",
112046=>"110110100",
112047=>"000001010",
112048=>"100000010",
112049=>"110111001",
112050=>"111011111",
112051=>"000000100",
112052=>"111111000",
112053=>"111000111",
112054=>"111110100",
112055=>"010111101",
112056=>"010110010",
112057=>"000010101",
112058=>"010010000",
112059=>"101000110",
112060=>"011100000",
112061=>"111111010",
112062=>"110011011",
112063=>"101011100",
112064=>"100100101",
112065=>"101000000",
112066=>"010000000",
112067=>"001100110",
112068=>"101101101",
112069=>"110010001",
112070=>"011000011",
112071=>"111001000",
112072=>"000000110",
112073=>"111111000",
112074=>"000101111",
112075=>"000000101",
112076=>"011011010",
112077=>"001000000",
112078=>"101000000",
112079=>"000100111",
112080=>"000010010",
112081=>"010001110",
112082=>"010010111",
112083=>"101101111",
112084=>"110010010",
112085=>"111001000",
112086=>"100111111",
112087=>"000001111",
112088=>"000000001",
112089=>"000001111",
112090=>"011001111",
112091=>"101101100",
112092=>"001101111",
112093=>"101111011",
112094=>"111111000",
112095=>"010111111",
112096=>"010101100",
112097=>"001000000",
112098=>"111111011",
112099=>"011101111",
112100=>"110100000",
112101=>"111111000",
112102=>"111010000",
112103=>"001011010",
112104=>"111000111",
112105=>"000111111",
112106=>"001001001",
112107=>"101100101",
112108=>"000101101",
112109=>"101110010",
112110=>"000110000",
112111=>"101101000",
112112=>"111111001",
112113=>"000110100",
112114=>"010001101",
112115=>"001000110",
112116=>"110110111",
112117=>"100000000",
112118=>"000010001",
112119=>"010000000",
112120=>"111111111",
112121=>"110000110",
112122=>"100111111",
112123=>"000001101",
112124=>"001000101",
112125=>"010110111",
112126=>"111000010",
112127=>"001001011",
112128=>"110100101",
112129=>"011010000",
112130=>"001001101",
112131=>"000000101",
112132=>"110011010",
112133=>"110110000",
112134=>"000000101",
112135=>"111011101",
112136=>"000100111",
112137=>"010010000",
112138=>"011100100",
112139=>"111100000",
112140=>"000111111",
112141=>"101111011",
112142=>"100111111",
112143=>"101001111",
112144=>"001010111",
112145=>"000000101",
112146=>"000010101",
112147=>"101010000",
112148=>"000100110",
112149=>"110111000",
112150=>"000100010",
112151=>"101000100",
112152=>"000001001",
112153=>"111000110",
112154=>"101111111",
112155=>"000101111",
112156=>"000010111",
112157=>"100000000",
112158=>"001000001",
112159=>"101101100",
112160=>"001000100",
112161=>"000101111",
112162=>"000010000",
112163=>"010011010",
112164=>"000100110",
112165=>"110110110",
112166=>"011111000",
112167=>"111000000",
112168=>"010011010",
112169=>"110111111",
112170=>"010100010",
112171=>"011101111",
112172=>"111000110",
112173=>"000000010",
112174=>"111011110",
112175=>"010000010",
112176=>"111000000",
112177=>"000101111",
112178=>"000000101",
112179=>"000010010",
112180=>"000101000",
112181=>"011001000",
112182=>"100110110",
112183=>"011001011",
112184=>"111101000",
112185=>"000010100",
112186=>"111000000",
112187=>"010011100",
112188=>"000000000",
112189=>"110111000",
112190=>"001100100",
112191=>"100100110",
112192=>"111111110",
112193=>"111111000",
112194=>"110000100",
112195=>"001001000",
112196=>"000000000",
112197=>"001001001",
112198=>"010000010",
112199=>"111111100",
112200=>"000000111",
112201=>"000000011",
112202=>"000000101",
112203=>"101101111",
112204=>"000000100",
112205=>"100011011",
112206=>"000100111",
112207=>"101001111",
112208=>"000100111",
112209=>"111010000",
112210=>"100000000",
112211=>"000000000",
112212=>"101000000",
112213=>"011001111",
112214=>"001011011",
112215=>"110010010",
112216=>"110100111",
112217=>"000000010",
112218=>"001110000",
112219=>"111000000",
112220=>"000000000",
112221=>"001001011",
112222=>"001001011",
112223=>"001000000",
112224=>"101000000",
112225=>"011110110",
112226=>"000000111",
112227=>"100011000",
112228=>"110101000",
112229=>"110110000",
112230=>"111111000",
112231=>"101101000",
112232=>"000000000",
112233=>"010010110",
112234=>"000000110",
112235=>"000111110",
112236=>"011111000",
112237=>"010010000",
112238=>"011000100",
112239=>"111111110",
112240=>"001101011",
112241=>"111101010",
112242=>"001001001",
112243=>"000000001",
112244=>"010000010",
112245=>"000000000",
112246=>"111001111",
112247=>"101111111",
112248=>"110111110",
112249=>"000000100",
112250=>"000010111",
112251=>"111110111",
112252=>"000110111",
112253=>"010010000",
112254=>"000000000",
112255=>"000101111",
112256=>"111101000",
112257=>"010001000",
112258=>"100000111",
112259=>"000101110",
112260=>"000010110",
112261=>"111100100",
112262=>"111011001",
112263=>"100000000",
112264=>"110111011",
112265=>"101111111",
112266=>"101010100",
112267=>"100101100",
112268=>"000011010",
112269=>"100101000",
112270=>"010011111",
112271=>"001001001",
112272=>"101100100",
112273=>"001001001",
112274=>"000000000",
112275=>"000000101",
112276=>"000010110",
112277=>"010000111",
112278=>"101110101",
112279=>"001011010",
112280=>"010001101",
112281=>"111100000",
112282=>"111111100",
112283=>"000000011",
112284=>"100000011",
112285=>"001000000",
112286=>"000100011",
112287=>"011000000",
112288=>"101000011",
112289=>"101101011",
112290=>"000010100",
112291=>"111001000",
112292=>"000100000",
112293=>"111000100",
112294=>"000000000",
112295=>"000000000",
112296=>"000000110",
112297=>"000110111",
112298=>"111111110",
112299=>"100000100",
112300=>"010110110",
112301=>"000001111",
112302=>"000100110",
112303=>"111000111",
112304=>"011000000",
112305=>"100000001",
112306=>"111011111",
112307=>"000000010",
112308=>"011011000",
112309=>"000010010",
112310=>"110101000",
112311=>"000011000",
112312=>"000000001",
112313=>"000010111",
112314=>"101000010",
112315=>"000100111",
112316=>"111010000",
112317=>"111111000",
112318=>"001011011",
112319=>"101111010",
112320=>"101000101",
112321=>"111000000",
112322=>"100110011",
112323=>"101111010",
112324=>"000010000",
112325=>"001000000",
112326=>"000000010",
112327=>"010010001",
112328=>"001010000",
112329=>"111101001",
112330=>"111111000",
112331=>"101111110",
112332=>"110010000",
112333=>"000011111",
112334=>"101111011",
112335=>"000111010",
112336=>"111111010",
112337=>"110100110",
112338=>"101000100",
112339=>"100111111",
112340=>"010010001",
112341=>"101111101",
112342=>"010000111",
112343=>"101010011",
112344=>"001000000",
112345=>"000000110",
112346=>"101000111",
112347=>"010000000",
112348=>"001111001",
112349=>"111111000",
112350=>"111101000",
112351=>"001010110",
112352=>"101101101",
112353=>"100100111",
112354=>"010111110",
112355=>"000110111",
112356=>"101000001",
112357=>"110100000",
112358=>"111100101",
112359=>"001011011",
112360=>"011000000",
112361=>"010011110",
112362=>"110000001",
112363=>"000010000",
112364=>"011111000",
112365=>"111111000",
112366=>"111111000",
112367=>"110000000",
112368=>"001110000",
112369=>"001000111",
112370=>"011000000",
112371=>"100000110",
112372=>"101001011",
112373=>"101111111",
112374=>"000010000",
112375=>"011100101",
112376=>"001000000",
112377=>"101000000",
112378=>"110001111",
112379=>"000101111",
112380=>"010010111",
112381=>"111101001",
112382=>"011110000",
112383=>"001000101",
112384=>"111110111",
112385=>"011000000",
112386=>"101000000",
112387=>"000100111",
112388=>"100011011",
112389=>"001011111",
112390=>"000011111",
112391=>"111111101",
112392=>"000011010",
112393=>"001000101",
112394=>"001000100",
112395=>"101100000",
112396=>"000011111",
112397=>"000110010",
112398=>"101100110",
112399=>"000000100",
112400=>"111000100",
112401=>"010010000",
112402=>"101000000",
112403=>"111111000",
112404=>"011000000",
112405=>"111001010",
112406=>"001110110",
112407=>"001011010",
112408=>"111101101",
112409=>"000000001",
112410=>"000011010",
112411=>"101000000",
112412=>"101100000",
112413=>"000001000",
112414=>"000111101",
112415=>"000010010",
112416=>"010000000",
112417=>"100111111",
112418=>"000000111",
112419=>"000111111",
112420=>"110110110",
112421=>"111001011",
112422=>"000011110",
112423=>"000000110",
112424=>"011011011",
112425=>"000000111",
112426=>"100100000",
112427=>"010000001",
112428=>"011000100",
112429=>"100100010",
112430=>"000000111",
112431=>"000001001",
112432=>"001000111",
112433=>"011011001",
112434=>"100110000",
112435=>"111111111",
112436=>"111001101",
112437=>"111101101",
112438=>"110110011",
112439=>"111100000",
112440=>"000000011",
112441=>"101100000",
112442=>"000001100",
112443=>"110000111",
112444=>"000100000",
112445=>"111111011",
112446=>"000000000",
112447=>"001011100",
112448=>"100000111",
112449=>"001000100",
112450=>"001000000",
112451=>"101111111",
112452=>"000101001",
112453=>"000000000",
112454=>"111001000",
112455=>"000011010",
112456=>"000100111",
112457=>"111100000",
112458=>"001101100",
112459=>"101000000",
112460=>"111100101",
112461=>"011011011",
112462=>"100100000",
112463=>"000000000",
112464=>"100110110",
112465=>"110111111",
112466=>"000011010",
112467=>"000011001",
112468=>"111000000",
112469=>"011110110",
112470=>"011011011",
112471=>"101000000",
112472=>"000010100",
112473=>"000001001",
112474=>"111100001",
112475=>"001011011",
112476=>"100000000",
112477=>"011010000",
112478=>"100111011",
112479=>"011101101",
112480=>"000000000",
112481=>"111110111",
112482=>"111100000",
112483=>"110110000",
112484=>"110000010",
112485=>"001000100",
112486=>"111000000",
112487=>"110101101",
112488=>"010000101",
112489=>"111111001",
112490=>"100111111",
112491=>"000001110",
112492=>"011001000",
112493=>"111010010",
112494=>"001100111",
112495=>"001000100",
112496=>"111100001",
112497=>"000000011",
112498=>"001011101",
112499=>"000111111",
112500=>"000100110",
112501=>"111000100",
112502=>"101000000",
112503=>"100000010",
112504=>"000000000",
112505=>"010000001",
112506=>"010000100",
112507=>"111111011",
112508=>"011111100",
112509=>"001010000",
112510=>"111010000",
112511=>"111101101",
112512=>"000000000",
112513=>"111111110",
112514=>"101000000",
112515=>"100000111",
112516=>"010111111",
112517=>"101000000",
112518=>"111100110",
112519=>"111000001",
112520=>"000111000",
112521=>"111000000",
112522=>"011110000",
112523=>"001011110",
112524=>"000000010",
112525=>"111101001",
112526=>"111101000",
112527=>"011000101",
112528=>"110100111",
112529=>"000000110",
112530=>"110000011",
112531=>"101101111",
112532=>"010010010",
112533=>"000111111",
112534=>"001000000",
112535=>"000000011",
112536=>"111101000",
112537=>"000101010",
112538=>"000111011",
112539=>"101011000",
112540=>"011100100",
112541=>"111100100",
112542=>"000100100",
112543=>"111100100",
112544=>"000001000",
112545=>"010000000",
112546=>"111001101",
112547=>"010000000",
112548=>"010011111",
112549=>"000000001",
112550=>"000110110",
112551=>"111111101",
112552=>"000111010",
112553=>"010000000",
112554=>"001110011",
112555=>"111000100",
112556=>"000000010",
112557=>"000010010",
112558=>"111101000",
112559=>"101010111",
112560=>"000000100",
112561=>"000110000",
112562=>"000100111",
112563=>"000100100",
112564=>"110001001",
112565=>"000001101",
112566=>"000000100",
112567=>"011111000",
112568=>"000001001",
112569=>"100111111",
112570=>"111101000",
112571=>"100111101",
112572=>"110111000",
112573=>"000010111",
112574=>"000110011",
112575=>"000100111",
112576=>"101000000",
112577=>"111000111",
112578=>"000001000",
112579=>"101110111",
112580=>"110000000",
112581=>"101000100",
112582=>"111111111",
112583=>"111111011",
112584=>"011001000",
112585=>"100101000",
112586=>"000011100",
112587=>"000000000",
112588=>"111100100",
112589=>"100101101",
112590=>"101101101",
112591=>"000111111",
112592=>"100111011",
112593=>"010100110",
112594=>"011000000",
112595=>"000101010",
112596=>"111000000",
112597=>"110011011",
112598=>"000100000",
112599=>"000000011",
112600=>"111000000",
112601=>"111111101",
112602=>"000011111",
112603=>"011101101",
112604=>"001011011",
112605=>"000011011",
112606=>"000000101",
112607=>"101111111",
112608=>"000000000",
112609=>"101000111",
112610=>"000111111",
112611=>"111101001",
112612=>"111000101",
112613=>"111000101",
112614=>"000000111",
112615=>"110011000",
112616=>"111111001",
112617=>"111111111",
112618=>"001100000",
112619=>"000000000",
112620=>"010111111",
112621=>"000111111",
112622=>"010000000",
112623=>"001000010",
112624=>"110111000",
112625=>"000010001",
112626=>"000000111",
112627=>"100110111",
112628=>"011011100",
112629=>"111000000",
112630=>"000000100",
112631=>"011001000",
112632=>"001111111",
112633=>"111111001",
112634=>"001000000",
112635=>"110110000",
112636=>"111110010",
112637=>"111111100",
112638=>"101111001",
112639=>"111100100",
112640=>"001001001",
112641=>"100101000",
112642=>"101000000",
112643=>"010101101",
112644=>"111000001",
112645=>"011101101",
112646=>"111101000",
112647=>"110111110",
112648=>"011000101",
112649=>"110011000",
112650=>"111000100",
112651=>"000111111",
112652=>"111110111",
112653=>"100110010",
112654=>"100000100",
112655=>"000000111",
112656=>"000110011",
112657=>"000000000",
112658=>"000000000",
112659=>"111001100",
112660=>"111000000",
112661=>"000000111",
112662=>"001000000",
112663=>"001010010",
112664=>"111000000",
112665=>"000110110",
112666=>"000101111",
112667=>"000000000",
112668=>"001000000",
112669=>"000000101",
112670=>"110111101",
112671=>"101000111",
112672=>"101101000",
112673=>"011110001",
112674=>"101010010",
112675=>"000000110",
112676=>"111111110",
112677=>"010001000",
112678=>"000010111",
112679=>"000010111",
112680=>"110010111",
112681=>"000110010",
112682=>"000110111",
112683=>"010000000",
112684=>"000011010",
112685=>"000011111",
112686=>"000110111",
112687=>"000101100",
112688=>"110111000",
112689=>"111101001",
112690=>"000111000",
112691=>"111101000",
112692=>"110000011",
112693=>"000101001",
112694=>"010110111",
112695=>"000000110",
112696=>"110111100",
112697=>"111000001",
112698=>"000000111",
112699=>"000000000",
112700=>"000110011",
112701=>"111011111",
112702=>"000000101",
112703=>"100101110",
112704=>"111000100",
112705=>"001101000",
112706=>"101111100",
112707=>"000000011",
112708=>"000000110",
112709=>"000000001",
112710=>"000000000",
112711=>"111000000",
112712=>"000111111",
112713=>"010000000",
112714=>"111001100",
112715=>"111111101",
112716=>"111111000",
112717=>"100001111",
112718=>"101001110",
112719=>"111110111",
112720=>"111001111",
112721=>"111111000",
112722=>"100111000",
112723=>"000111000",
112724=>"000000100",
112725=>"000110111",
112726=>"111111111",
112727=>"000111010",
112728=>"110000010",
112729=>"000000001",
112730=>"110000000",
112731=>"000111101",
112732=>"000000000",
112733=>"000000000",
112734=>"000011011",
112735=>"111000000",
112736=>"000011111",
112737=>"010000000",
112738=>"111000000",
112739=>"011011000",
112740=>"001000001",
112741=>"100111010",
112742=>"000000111",
112743=>"001000000",
112744=>"011101101",
112745=>"111111111",
112746=>"101111111",
112747=>"000101111",
112748=>"000111111",
112749=>"111000010",
112750=>"111100000",
112751=>"001101000",
112752=>"000110100",
112753=>"000000111",
112754=>"000010111",
112755=>"011000000",
112756=>"001001000",
112757=>"010001100",
112758=>"000000111",
112759=>"000001000",
112760=>"110111000",
112761=>"011000100",
112762=>"010000001",
112763=>"101000001",
112764=>"000000001",
112765=>"000110000",
112766=>"000111111",
112767=>"111000011",
112768=>"011111101",
112769=>"111101000",
112770=>"000011011",
112771=>"000000111",
112772=>"111110111",
112773=>"101111000",
112774=>"100111100",
112775=>"111000100",
112776=>"100100001",
112777=>"000000001",
112778=>"111110001",
112779=>"101111011",
112780=>"111010000",
112781=>"111101000",
112782=>"100000000",
112783=>"111000001",
112784=>"011001100",
112785=>"000000000",
112786=>"000111001",
112787=>"000111101",
112788=>"111000110",
112789=>"000111000",
112790=>"111111000",
112791=>"010000001",
112792=>"110111111",
112793=>"110100000",
112794=>"000110111",
112795=>"101110000",
112796=>"111111110",
112797=>"000010010",
112798=>"111111000",
112799=>"100101111",
112800=>"011001100",
112801=>"011000000",
112802=>"000101111",
112803=>"111000000",
112804=>"000111101",
112805=>"010000001",
112806=>"000000111",
112807=>"010011111",
112808=>"000000010",
112809=>"000000100",
112810=>"100000010",
112811=>"101001001",
112812=>"001001010",
112813=>"011110111",
112814=>"000000111",
112815=>"111111111",
112816=>"000000000",
112817=>"111000011",
112818=>"000111011",
112819=>"101000100",
112820=>"000000001",
112821=>"101111010",
112822=>"000001000",
112823=>"101111011",
112824=>"001011010",
112825=>"011001001",
112826=>"011000000",
112827=>"010111110",
112828=>"010101101",
112829=>"111011011",
112830=>"000000001",
112831=>"011101000",
112832=>"010110111",
112833=>"101111000",
112834=>"111111111",
112835=>"100101111",
112836=>"000110111",
112837=>"001011001",
112838=>"010111101",
112839=>"111000000",
112840=>"011111011",
112841=>"000000000",
112842=>"101000000",
112843=>"111101100",
112844=>"000010011",
112845=>"100000110",
112846=>"111000101",
112847=>"111101000",
112848=>"100000111",
112849=>"101000100",
112850=>"011000001",
112851=>"000000000",
112852=>"000010110",
112853=>"111001111",
112854=>"111101111",
112855=>"000111011",
112856=>"000111111",
112857=>"011000111",
112858=>"101000000",
112859=>"111111000",
112860=>"000110000",
112861=>"110001010",
112862=>"010001011",
112863=>"100110111",
112864=>"111000000",
112865=>"111001111",
112866=>"111111111",
112867=>"001000100",
112868=>"111000101",
112869=>"110000000",
112870=>"000110000",
112871=>"000000000",
112872=>"100111111",
112873=>"011000101",
112874=>"001000011",
112875=>"111001000",
112876=>"000010011",
112877=>"010111111",
112878=>"111000001",
112879=>"000010111",
112880=>"000111101",
112881=>"110011111",
112882=>"000111111",
112883=>"000000110",
112884=>"011110110",
112885=>"111101000",
112886=>"101000000",
112887=>"010111111",
112888=>"000110010",
112889=>"010111101",
112890=>"001000000",
112891=>"001001111",
112892=>"000010111",
112893=>"111100000",
112894=>"100100100",
112895=>"010110110",
112896=>"001001101",
112897=>"111111000",
112898=>"000000101",
112899=>"000001000",
112900=>"000011011",
112901=>"000000110",
112902=>"000110100",
112903=>"000110110",
112904=>"000110000",
112905=>"011001101",
112906=>"010010010",
112907=>"101111000",
112908=>"100111110",
112909=>"101100000",
112910=>"000111011",
112911=>"101100000",
112912=>"110111111",
112913=>"111000111",
112914=>"100000000",
112915=>"000000010",
112916=>"110000100",
112917=>"111000000",
112918=>"000010011",
112919=>"101000111",
112920=>"001000000",
112921=>"111011000",
112922=>"000000010",
112923=>"001111111",
112924=>"101110000",
112925=>"100000000",
112926=>"111000011",
112927=>"011001000",
112928=>"010011111",
112929=>"000000110",
112930=>"111000010",
112931=>"111100011",
112932=>"100111011",
112933=>"101101010",
112934=>"111010000",
112935=>"000100100",
112936=>"111000000",
112937=>"000111100",
112938=>"000000000",
112939=>"101111010",
112940=>"100111111",
112941=>"111001111",
112942=>"000100011",
112943=>"000100001",
112944=>"111000000",
112945=>"001100100",
112946=>"111010001",
112947=>"000100110",
112948=>"101001111",
112949=>"111100111",
112950=>"000000011",
112951=>"011110000",
112952=>"111000110",
112953=>"000100110",
112954=>"100000000",
112955=>"111111111",
112956=>"011111110",
112957=>"111111101",
112958=>"000000101",
112959=>"110110111",
112960=>"100100111",
112961=>"000110110",
112962=>"001000011",
112963=>"001110100",
112964=>"000001000",
112965=>"100110100",
112966=>"000100110",
112967=>"000101101",
112968=>"111001101",
112969=>"101011111",
112970=>"000110110",
112971=>"101111111",
112972=>"000000011",
112973=>"011011110",
112974=>"000001011",
112975=>"101001110",
112976=>"000001000",
112977=>"111111111",
112978=>"111010111",
112979=>"001001000",
112980=>"110000000",
112981=>"110100110",
112982=>"001001110",
112983=>"111011101",
112984=>"000001000",
112985=>"000100110",
112986=>"011101100",
112987=>"011000000",
112988=>"010111000",
112989=>"000001001",
112990=>"111011000",
112991=>"111000000",
112992=>"000000010",
112993=>"111000111",
112994=>"000000111",
112995=>"100011111",
112996=>"000110101",
112997=>"000000101",
112998=>"000111100",
112999=>"110000000",
113000=>"110011100",
113001=>"111000111",
113002=>"000000111",
113003=>"000000110",
113004=>"010010111",
113005=>"111111000",
113006=>"000000000",
113007=>"001111110",
113008=>"110001011",
113009=>"010000000",
113010=>"001100110",
113011=>"010000000",
113012=>"000000010",
113013=>"001000000",
113014=>"000100000",
113015=>"000010000",
113016=>"000110000",
113017=>"011111010",
113018=>"110111001",
113019=>"111111101",
113020=>"101101101",
113021=>"100100000",
113022=>"110000000",
113023=>"111000000",
113024=>"000000000",
113025=>"010000010",
113026=>"010010000",
113027=>"011110110",
113028=>"101101111",
113029=>"110011100",
113030=>"001100110",
113031=>"011101100",
113032=>"011111110",
113033=>"101111110",
113034=>"011011001",
113035=>"101100000",
113036=>"111000000",
113037=>"110000000",
113038=>"111110000",
113039=>"000101000",
113040=>"001001011",
113041=>"000111111",
113042=>"111001000",
113043=>"000110101",
113044=>"011001111",
113045=>"010000101",
113046=>"010111010",
113047=>"011010100",
113048=>"110010000",
113049=>"111111101",
113050=>"111011001",
113051=>"000000000",
113052=>"000001010",
113053=>"100110010",
113054=>"000000111",
113055=>"000101111",
113056=>"000010011",
113057=>"010111111",
113058=>"000111101",
113059=>"011111000",
113060=>"100110111",
113061=>"100110010",
113062=>"110110000",
113063=>"000111100",
113064=>"010010011",
113065=>"000000010",
113066=>"111000000",
113067=>"000000000",
113068=>"010111111",
113069=>"000000111",
113070=>"100100111",
113071=>"011010000",
113072=>"110110000",
113073=>"011011011",
113074=>"000001000",
113075=>"100100001",
113076=>"111111010",
113077=>"010010000",
113078=>"010011100",
113079=>"001001000",
113080=>"110111100",
113081=>"000111010",
113082=>"010000000",
113083=>"011011110",
113084=>"010001000",
113085=>"000000000",
113086=>"011010011",
113087=>"110000000",
113088=>"001101011",
113089=>"010010011",
113090=>"111110000",
113091=>"001001110",
113092=>"000101000",
113093=>"100101101",
113094=>"110000000",
113095=>"000001101",
113096=>"000000111",
113097=>"000111010",
113098=>"010110000",
113099=>"111110010",
113100=>"000011010",
113101=>"000100000",
113102=>"010000000",
113103=>"111110111",
113104=>"001111111",
113105=>"000111111",
113106=>"111101110",
113107=>"101000000",
113108=>"011000000",
113109=>"110111100",
113110=>"000000111",
113111=>"000011111",
113112=>"111000000",
113113=>"011100000",
113114=>"000000110",
113115=>"111000000",
113116=>"010110110",
113117=>"111100000",
113118=>"111010000",
113119=>"010001101",
113120=>"000111111",
113121=>"110100101",
113122=>"111011000",
113123=>"100110111",
113124=>"000000000",
113125=>"110011111",
113126=>"000100111",
113127=>"010011011",
113128=>"000000001",
113129=>"010011000",
113130=>"111011011",
113131=>"010010000",
113132=>"111010000",
113133=>"000001000",
113134=>"111001000",
113135=>"011000000",
113136=>"110100000",
113137=>"011001111",
113138=>"001000000",
113139=>"000010001",
113140=>"110110111",
113141=>"001011010",
113142=>"001000000",
113143=>"111111000",
113144=>"010011000",
113145=>"000000000",
113146=>"111101100",
113147=>"000101111",
113148=>"010111101",
113149=>"111000000",
113150=>"010111111",
113151=>"000111111",
113152=>"100100110",
113153=>"000000110",
113154=>"011000111",
113155=>"001000100",
113156=>"001000001",
113157=>"111010000",
113158=>"111001000",
113159=>"110010111",
113160=>"001011011",
113161=>"000110010",
113162=>"001100100",
113163=>"101111010",
113164=>"111000000",
113165=>"010011000",
113166=>"110001001",
113167=>"111000001",
113168=>"000111101",
113169=>"000111100",
113170=>"111000001",
113171=>"000101111",
113172=>"001110111",
113173=>"001000110",
113174=>"111010001",
113175=>"111111111",
113176=>"110000000",
113177=>"000001111",
113178=>"000100110",
113179=>"000100000",
113180=>"100000010",
113181=>"111000000",
113182=>"111111011",
113183=>"010101000",
113184=>"011000000",
113185=>"000010000",
113186=>"111100000",
113187=>"000001000",
113188=>"010000001",
113189=>"001100110",
113190=>"101100111",
113191=>"000110010",
113192=>"010000000",
113193=>"010100010",
113194=>"000101111",
113195=>"000010110",
113196=>"010110001",
113197=>"000000110",
113198=>"101111001",
113199=>"010101111",
113200=>"111110000",
113201=>"111100000",
113202=>"000001101",
113203=>"111111110",
113204=>"011001100",
113205=>"000000000",
113206=>"001001000",
113207=>"000010000",
113208=>"111111010",
113209=>"110010111",
113210=>"111000101",
113211=>"000001111",
113212=>"011001001",
113213=>"000010000",
113214=>"000000011",
113215=>"001011111",
113216=>"111111111",
113217=>"100100100",
113218=>"001001111",
113219=>"001000101",
113220=>"100010110",
113221=>"010011001",
113222=>"111111000",
113223=>"011111100",
113224=>"100010001",
113225=>"000111110",
113226=>"000110000",
113227=>"001011101",
113228=>"111111100",
113229=>"001001000",
113230=>"010000100",
113231=>"100111111",
113232=>"111101000",
113233=>"001000000",
113234=>"000111000",
113235=>"111111000",
113236=>"000000000",
113237=>"010001101",
113238=>"110101101",
113239=>"010111111",
113240=>"001011111",
113241=>"111001001",
113242=>"010100100",
113243=>"100110110",
113244=>"000011011",
113245=>"110000001",
113246=>"110000111",
113247=>"011001000",
113248=>"000101111",
113249=>"000000110",
113250=>"101001111",
113251=>"110110001",
113252=>"111000000",
113253=>"011110001",
113254=>"000110110",
113255=>"111001000",
113256=>"110111000",
113257=>"000111111",
113258=>"110010101",
113259=>"111001110",
113260=>"000101101",
113261=>"100001011",
113262=>"111111000",
113263=>"101000000",
113264=>"111011000",
113265=>"101110110",
113266=>"100110000",
113267=>"111101111",
113268=>"111010000",
113269=>"110001000",
113270=>"000000110",
113271=>"000101111",
113272=>"110100100",
113273=>"111111110",
113274=>"010000010",
113275=>"110000000",
113276=>"110110100",
113277=>"011011000",
113278=>"001111010",
113279=>"111101101",
113280=>"111111000",
113281=>"110010000",
113282=>"000101111",
113283=>"000111100",
113284=>"111111010",
113285=>"110101100",
113286=>"000001111",
113287=>"000011101",
113288=>"110100000",
113289=>"010000000",
113290=>"111101000",
113291=>"100101000",
113292=>"110010000",
113293=>"111000001",
113294=>"101111000",
113295=>"001001111",
113296=>"111000100",
113297=>"111001000",
113298=>"000010111",
113299=>"111111001",
113300=>"111111001",
113301=>"110000110",
113302=>"110111111",
113303=>"010001001",
113304=>"000101111",
113305=>"110000111",
113306=>"111010111",
113307=>"110000101",
113308=>"110011011",
113309=>"000110110",
113310=>"101111100",
113311=>"111110110",
113312=>"110001001",
113313=>"000101000",
113314=>"001011000",
113315=>"000111111",
113316=>"111110011",
113317=>"011001001",
113318=>"011011111",
113319=>"000101001",
113320=>"000111101",
113321=>"000100111",
113322=>"111110001",
113323=>"111010010",
113324=>"111001000",
113325=>"111100111",
113326=>"011001000",
113327=>"000111111",
113328=>"110000000",
113329=>"110111000",
113330=>"010000101",
113331=>"000000100",
113332=>"110100000",
113333=>"110111101",
113334=>"000000000",
113335=>"111001011",
113336=>"100100000",
113337=>"110110111",
113338=>"100000000",
113339=>"111111000",
113340=>"101000000",
113341=>"000111111",
113342=>"100110110",
113343=>"101000000",
113344=>"111001100",
113345=>"000111111",
113346=>"111110110",
113347=>"110100000",
113348=>"000000001",
113349=>"111010010",
113350=>"111100011",
113351=>"100110111",
113352=>"111111001",
113353=>"010000000",
113354=>"111111111",
113355=>"000111111",
113356=>"101111111",
113357=>"001011001",
113358=>"111111000",
113359=>"000000000",
113360=>"000000111",
113361=>"111110101",
113362=>"010010010",
113363=>"111100100",
113364=>"101110010",
113365=>"011011100",
113366=>"111111111",
113367=>"000011110",
113368=>"000101111",
113369=>"111101100",
113370=>"011001101",
113371=>"111101000",
113372=>"110110101",
113373=>"111000111",
113374=>"101101010",
113375=>"100111110",
113376=>"000001101",
113377=>"111011000",
113378=>"111000101",
113379=>"111011000",
113380=>"000000100",
113381=>"000111010",
113382=>"111111111",
113383=>"100100001",
113384=>"010111111",
113385=>"110000000",
113386=>"100000011",
113387=>"000101111",
113388=>"111101001",
113389=>"111001101",
113390=>"000000000",
113391=>"010000000",
113392=>"111101000",
113393=>"111011111",
113394=>"100110000",
113395=>"010010101",
113396=>"011011001",
113397=>"010000000",
113398=>"100100011",
113399=>"011010000",
113400=>"000010101",
113401=>"001001100",
113402=>"111110000",
113403=>"010110101",
113404=>"111110111",
113405=>"000000111",
113406=>"011000000",
113407=>"000111010",
113408=>"111101100",
113409=>"001101100",
113410=>"001000000",
113411=>"111001001",
113412=>"010001000",
113413=>"000000001",
113414=>"111111000",
113415=>"000010110",
113416=>"111110000",
113417=>"000010000",
113418=>"001001000",
113419=>"101000100",
113420=>"111000101",
113421=>"110110001",
113422=>"001011000",
113423=>"001101110",
113424=>"010000010",
113425=>"000000001",
113426=>"000000011",
113427=>"110111110",
113428=>"111111100",
113429=>"000001001",
113430=>"111101101",
113431=>"101000011",
113432=>"100111000",
113433=>"111111000",
113434=>"010000000",
113435=>"000100101",
113436=>"000111111",
113437=>"000001101",
113438=>"110000111",
113439=>"101001000",
113440=>"000111000",
113441=>"111101111",
113442=>"111100000",
113443=>"111111010",
113444=>"011011000",
113445=>"100101100",
113446=>"110010000",
113447=>"100010010",
113448=>"001001100",
113449=>"110010000",
113450=>"001000010",
113451=>"001000111",
113452=>"111111100",
113453=>"000010110",
113454=>"111010101",
113455=>"001000111",
113456=>"001001110",
113457=>"101000000",
113458=>"000000000",
113459=>"001001101",
113460=>"000000111",
113461=>"101000000",
113462=>"100110101",
113463=>"000000111",
113464=>"010011110",
113465=>"100000000",
113466=>"010000000",
113467=>"101111000",
113468=>"100100011",
113469=>"011111101",
113470=>"000000100",
113471=>"011111000",
113472=>"101001000",
113473=>"010111101",
113474=>"111111111",
113475=>"000100110",
113476=>"100111101",
113477=>"010000010",
113478=>"111100000",
113479=>"110010110",
113480=>"111010110",
113481=>"000101111",
113482=>"000000001",
113483=>"110100000",
113484=>"010110000",
113485=>"011101000",
113486=>"001100000",
113487=>"001111111",
113488=>"101001000",
113489=>"001011111",
113490=>"111101111",
113491=>"011001101",
113492=>"001000110",
113493=>"000000010",
113494=>"100111110",
113495=>"111111000",
113496=>"010000110",
113497=>"110110010",
113498=>"100100000",
113499=>"110110000",
113500=>"000000000",
113501=>"001000000",
113502=>"010110110",
113503=>"000001000",
113504=>"110111000",
113505=>"011001111",
113506=>"010000000",
113507=>"111001000",
113508=>"001111000",
113509=>"001011101",
113510=>"000111010",
113511=>"000000000",
113512=>"111111000",
113513=>"000000010",
113514=>"110010111",
113515=>"111001011",
113516=>"000111000",
113517=>"000000111",
113518=>"111100110",
113519=>"000110110",
113520=>"101100100",
113521=>"111101101",
113522=>"011011101",
113523=>"001001000",
113524=>"010000100",
113525=>"000000000",
113526=>"111110111",
113527=>"111000000",
113528=>"000000110",
113529=>"010111010",
113530=>"111111111",
113531=>"011000111",
113532=>"110110100",
113533=>"100100100",
113534=>"011100010",
113535=>"001000000",
113536=>"111110110",
113537=>"111001000",
113538=>"110000111",
113539=>"111101110",
113540=>"100000011",
113541=>"111110110",
113542=>"001000011",
113543=>"011011000",
113544=>"101111000",
113545=>"000001101",
113546=>"000000000",
113547=>"111111111",
113548=>"001000101",
113549=>"101000001",
113550=>"001010110",
113551=>"001001000",
113552=>"111100000",
113553=>"001001001",
113554=>"110111000",
113555=>"000000111",
113556=>"011000100",
113557=>"111110110",
113558=>"110110110",
113559=>"011011011",
113560=>"001011101",
113561=>"000111111",
113562=>"010111000",
113563=>"100000110",
113564=>"010111000",
113565=>"000110111",
113566=>"000010111",
113567=>"111111101",
113568=>"111110010",
113569=>"111000111",
113570=>"111110110",
113571=>"000000000",
113572=>"010001011",
113573=>"011111100",
113574=>"011110101",
113575=>"010111010",
113576=>"000001111",
113577=>"000110111",
113578=>"001000000",
113579=>"000010001",
113580=>"111000110",
113581=>"110010000",
113582=>"100101100",
113583=>"001000000",
113584=>"001000000",
113585=>"110100000",
113586=>"011010000",
113587=>"000110000",
113588=>"101111111",
113589=>"000001101",
113590=>"100001000",
113591=>"101110111",
113592=>"001011000",
113593=>"110110101",
113594=>"110000000",
113595=>"110110000",
113596=>"100000010",
113597=>"101111111",
113598=>"110110000",
113599=>"000000101",
113600=>"110100000",
113601=>"001001100",
113602=>"010000111",
113603=>"111101000",
113604=>"000010000",
113605=>"000001011",
113606=>"000011000",
113607=>"010000000",
113608=>"101111010",
113609=>"000000000",
113610=>"001000000",
113611=>"000111111",
113612=>"000111111",
113613=>"111011001",
113614=>"101111101",
113615=>"110111100",
113616=>"001000111",
113617=>"010110100",
113618=>"111111000",
113619=>"000000111",
113620=>"000010111",
113621=>"011001110",
113622=>"110000111",
113623=>"110000000",
113624=>"110000111",
113625=>"000000001",
113626=>"111111000",
113627=>"000000101",
113628=>"000001100",
113629=>"101000000",
113630=>"000000000",
113631=>"000001010",
113632=>"000000001",
113633=>"101001111",
113634=>"001000111",
113635=>"111011100",
113636=>"111101100",
113637=>"111010000",
113638=>"111100001",
113639=>"011011011",
113640=>"000001000",
113641=>"000000111",
113642=>"001000101",
113643=>"111000001",
113644=>"000000001",
113645=>"000000000",
113646=>"010000000",
113647=>"101100100",
113648=>"101101001",
113649=>"010000010",
113650=>"110010100",
113651=>"011011110",
113652=>"111111001",
113653=>"010011000",
113654=>"000010010",
113655=>"101000110",
113656=>"000111111",
113657=>"010010110",
113658=>"111000001",
113659=>"110010000",
113660=>"101111010",
113661=>"000000110",
113662=>"100111000",
113663=>"001001111",
113664=>"100000000",
113665=>"101000000",
113666=>"000000000",
113667=>"001000111",
113668=>"000011011",
113669=>"001011111",
113670=>"111100100",
113671=>"111000100",
113672=>"000000011",
113673=>"001000000",
113674=>"100010011",
113675=>"100100110",
113676=>"010011010",
113677=>"001011000",
113678=>"100100110",
113679=>"111101011",
113680=>"111010001",
113681=>"001011111",
113682=>"101001101",
113683=>"011110000",
113684=>"011001000",
113685=>"100111010",
113686=>"000111010",
113687=>"110111111",
113688=>"111101000",
113689=>"110000000",
113690=>"100000000",
113691=>"000010010",
113692=>"100000000",
113693=>"100100111",
113694=>"000100111",
113695=>"000000100",
113696=>"111101111",
113697=>"000010100",
113698=>"100101111",
113699=>"000100001",
113700=>"010010000",
113701=>"100001000",
113702=>"111100000",
113703=>"001110101",
113704=>"011000000",
113705=>"001000011",
113706=>"101100000",
113707=>"000010111",
113708=>"000011001",
113709=>"101010010",
113710=>"010010111",
113711=>"000111101",
113712=>"101111111",
113713=>"011001000",
113714=>"111111101",
113715=>"110100000",
113716=>"000010000",
113717=>"111111111",
113718=>"101111100",
113719=>"000100101",
113720=>"000111100",
113721=>"101101101",
113722=>"111111101",
113723=>"000110000",
113724=>"000001001",
113725=>"101111101",
113726=>"000000111",
113727=>"001000010",
113728=>"100111111",
113729=>"001100110",
113730=>"000000011",
113731=>"100100000",
113732=>"000010000",
113733=>"000101110",
113734=>"010000000",
113735=>"001000111",
113736=>"101010001",
113737=>"001000000",
113738=>"101101100",
113739=>"111100101",
113740=>"000100101",
113741=>"111011001",
113742=>"101110100",
113743=>"010000000",
113744=>"111000000",
113745=>"111000100",
113746=>"000000101",
113747=>"000000001",
113748=>"000000001",
113749=>"011001101",
113750=>"000100010",
113751=>"111100100",
113752=>"000000101",
113753=>"000000101",
113754=>"000000000",
113755=>"000110010",
113756=>"010000000",
113757=>"000010000",
113758=>"010111000",
113759=>"100100100",
113760=>"100100001",
113761=>"001000000",
113762=>"000011100",
113763=>"001011001",
113764=>"011000111",
113765=>"001111111",
113766=>"110011100",
113767=>"100000011",
113768=>"110101000",
113769=>"011111111",
113770=>"111111100",
113771=>"001100100",
113772=>"000101111",
113773=>"000101110",
113774=>"000000000",
113775=>"100000100",
113776=>"000110110",
113777=>"000011100",
113778=>"010011011",
113779=>"111101111",
113780=>"011000000",
113781=>"101111010",
113782=>"000111111",
113783=>"000100011",
113784=>"000001000",
113785=>"011011101",
113786=>"111111111",
113787=>"111111101",
113788=>"011001000",
113789=>"000001000",
113790=>"111111110",
113791=>"111100110",
113792=>"100101110",
113793=>"000000000",
113794=>"000011000",
113795=>"100100111",
113796=>"000010000",
113797=>"111111111",
113798=>"000100100",
113799=>"010000000",
113800=>"001001100",
113801=>"000000110",
113802=>"111101000",
113803=>"000011111",
113804=>"111100000",
113805=>"111101111",
113806=>"000000010",
113807=>"111000001",
113808=>"101110001",
113809=>"010111101",
113810=>"000100100",
113811=>"010000000",
113812=>"111000100",
113813=>"111010000",
113814=>"100000000",
113815=>"110010001",
113816=>"101001110",
113817=>"111000000",
113818=>"000011001",
113819=>"000010011",
113820=>"111100000",
113821=>"000000000",
113822=>"001000011",
113823=>"000100101",
113824=>"010100110",
113825=>"001000101",
113826=>"100001111",
113827=>"000000101",
113828=>"000000011",
113829=>"110101101",
113830=>"100000110",
113831=>"000111111",
113832=>"100111000",
113833=>"000000110",
113834=>"000011011",
113835=>"000000010",
113836=>"010100111",
113837=>"111000001",
113838=>"100100100",
113839=>"111111111",
113840=>"110011011",
113841=>"111110001",
113842=>"000000010",
113843=>"000000001",
113844=>"001001011",
113845=>"101111000",
113846=>"000000100",
113847=>"000011111",
113848=>"000000000",
113849=>"010000000",
113850=>"111011010",
113851=>"101111111",
113852=>"110100000",
113853=>"011111111",
113854=>"010000000",
113855=>"001111111",
113856=>"111000000",
113857=>"101100000",
113858=>"111001000",
113859=>"110000000",
113860=>"100100111",
113861=>"011001111",
113862=>"000011000",
113863=>"111011101",
113864=>"010100101",
113865=>"000100111",
113866=>"000000100",
113867=>"000100000",
113868=>"111100011",
113869=>"110000100",
113870=>"000010011",
113871=>"011000010",
113872=>"100111111",
113873=>"101110110",
113874=>"100000100",
113875=>"111111111",
113876=>"000000000",
113877=>"011011011",
113878=>"000000000",
113879=>"001000001",
113880=>"100100000",
113881=>"000100000",
113882=>"110001101",
113883=>"011111111",
113884=>"110111110",
113885=>"111011011",
113886=>"101101000",
113887=>"000100111",
113888=>"100000000",
113889=>"001011011",
113890=>"011010011",
113891=>"010100101",
113892=>"001000000",
113893=>"000011010",
113894=>"111111111",
113895=>"000101100",
113896=>"010111101",
113897=>"111111000",
113898=>"001001000",
113899=>"001000000",
113900=>"100000000",
113901=>"000100100",
113902=>"101010100",
113903=>"000000111",
113904=>"000000101",
113905=>"010100011",
113906=>"100000111",
113907=>"100100000",
113908=>"001001100",
113909=>"111011000",
113910=>"000000101",
113911=>"000010010",
113912=>"011111000",
113913=>"010111011",
113914=>"111111110",
113915=>"000000111",
113916=>"100100000",
113917=>"000111110",
113918=>"111111111",
113919=>"100000100",
113920=>"010000010",
113921=>"000011111",
113922=>"000000000",
113923=>"000110111",
113924=>"111101000",
113925=>"111000010",
113926=>"111111111",
113927=>"111101101",
113928=>"000101111",
113929=>"000000100",
113930=>"000100000",
113931=>"101000100",
113932=>"110000000",
113933=>"111011011",
113934=>"010100100",
113935=>"111010000",
113936=>"100011010",
113937=>"000000110",
113938=>"000111000",
113939=>"011000011",
113940=>"010010000",
113941=>"000000111",
113942=>"000011111",
113943=>"000111111",
113944=>"111000100",
113945=>"111010000",
113946=>"000000111",
113947=>"000111111",
113948=>"101111111",
113949=>"000000011",
113950=>"010000011",
113951=>"010011111",
113952=>"111000010",
113953=>"010011000",
113954=>"000111101",
113955=>"010010000",
113956=>"000111111",
113957=>"000001011",
113958=>"000100111",
113959=>"000100000",
113960=>"011111100",
113961=>"000100000",
113962=>"100110000",
113963=>"111101001",
113964=>"111011010",
113965=>"100100000",
113966=>"000100010",
113967=>"000000101",
113968=>"101100000",
113969=>"000000011",
113970=>"000000000",
113971=>"111111100",
113972=>"000000010",
113973=>"001100100",
113974=>"011011011",
113975=>"100000100",
113976=>"111010000",
113977=>"011111011",
113978=>"000000000",
113979=>"110111000",
113980=>"111011001",
113981=>"011111000",
113982=>"100100001",
113983=>"101101110",
113984=>"111101000",
113985=>"100111111",
113986=>"111100001",
113987=>"111100000",
113988=>"111111000",
113989=>"000100100",
113990=>"111111011",
113991=>"010111111",
113992=>"000111001",
113993=>"111110111",
113994=>"000000000",
113995=>"000100001",
113996=>"000000000",
113997=>"000111111",
113998=>"111111010",
113999=>"000000000",
114000=>"010010011",
114001=>"111111110",
114002=>"111001111",
114003=>"001000000",
114004=>"100100111",
114005=>"101111111",
114006=>"001111110",
114007=>"101100111",
114008=>"000000001",
114009=>"011001000",
114010=>"101111111",
114011=>"011111111",
114012=>"000011010",
114013=>"000000000",
114014=>"001111010",
114015=>"100101100",
114016=>"111001010",
114017=>"111000000",
114018=>"101100111",
114019=>"100110110",
114020=>"000010010",
114021=>"000000001",
114022=>"000011011",
114023=>"100000000",
114024=>"111111000",
114025=>"000000001",
114026=>"010101111",
114027=>"111101000",
114028=>"000000000",
114029=>"000100110",
114030=>"010000000",
114031=>"000000011",
114032=>"111111111",
114033=>"010000000",
114034=>"111110011",
114035=>"100000010",
114036=>"000000101",
114037=>"100100000",
114038=>"111011111",
114039=>"110100111",
114040=>"110000000",
114041=>"010110110",
114042=>"000111111",
114043=>"100100101",
114044=>"010001001",
114045=>"100000011",
114046=>"110011000",
114047=>"101100100",
114048=>"011010000",
114049=>"111000000",
114050=>"100011111",
114051=>"000000100",
114052=>"111100111",
114053=>"010100000",
114054=>"111110111",
114055=>"011010010",
114056=>"111001011",
114057=>"001000000",
114058=>"111100101",
114059=>"100100101",
114060=>"011011000",
114061=>"000000010",
114062=>"101000000",
114063=>"100000001",
114064=>"110111110",
114065=>"001011111",
114066=>"011011000",
114067=>"011101010",
114068=>"111001100",
114069=>"100000100",
114070=>"000010011",
114071=>"100000000",
114072=>"000010000",
114073=>"111001001",
114074=>"100110000",
114075=>"100100100",
114076=>"111011011",
114077=>"111101000",
114078=>"111011111",
114079=>"100100001",
114080=>"100111011",
114081=>"000111010",
114082=>"010111111",
114083=>"110100100",
114084=>"000000100",
114085=>"111010000",
114086=>"001111011",
114087=>"000000011",
114088=>"010011111",
114089=>"000000000",
114090=>"100000100",
114091=>"100000111",
114092=>"000011000",
114093=>"101000110",
114094=>"100110010",
114095=>"111110100",
114096=>"001010000",
114097=>"100111100",
114098=>"000100000",
114099=>"000010001",
114100=>"000000000",
114101=>"011111000",
114102=>"011011000",
114103=>"011000110",
114104=>"011010110",
114105=>"110111001",
114106=>"111111010",
114107=>"010111111",
114108=>"111101000",
114109=>"111111110",
114110=>"001001101",
114111=>"010000001",
114112=>"000000000",
114113=>"000000000",
114114=>"011001000",
114115=>"000111111",
114116=>"000100100",
114117=>"010110111",
114118=>"010111011",
114119=>"000000011",
114120=>"101000000",
114121=>"000000000",
114122=>"111011000",
114123=>"011011111",
114124=>"000000101",
114125=>"000010011",
114126=>"000011011",
114127=>"000100111",
114128=>"110000010",
114129=>"100010110",
114130=>"111100111",
114131=>"011000000",
114132=>"111101110",
114133=>"000100000",
114134=>"000100110",
114135=>"100000111",
114136=>"000000000",
114137=>"000000000",
114138=>"000010111",
114139=>"100000000",
114140=>"100110111",
114141=>"100010111",
114142=>"111011000",
114143=>"111010010",
114144=>"011011011",
114145=>"101100011",
114146=>"111110110",
114147=>"101111111",
114148=>"100100100",
114149=>"000101110",
114150=>"111000011",
114151=>"000110110",
114152=>"011000000",
114153=>"000001111",
114154=>"001000000",
114155=>"010010100",
114156=>"000111101",
114157=>"111011001",
114158=>"000100111",
114159=>"000000000",
114160=>"100100100",
114161=>"000101111",
114162=>"000101111",
114163=>"110000011",
114164=>"110111001",
114165=>"111100111",
114166=>"010000100",
114167=>"000100001",
114168=>"011111110",
114169=>"111100000",
114170=>"010000000",
114171=>"000000001",
114172=>"001000010",
114173=>"000100000",
114174=>"000111001",
114175=>"101000000",
114176=>"110110000",
114177=>"000000001",
114178=>"000000000",
114179=>"010000000",
114180=>"000111101",
114181=>"011001001",
114182=>"111000000",
114183=>"110101001",
114184=>"101111000",
114185=>"011000000",
114186=>"110011011",
114187=>"000001111",
114188=>"000000000",
114189=>"110111101",
114190=>"011100100",
114191=>"000010000",
114192=>"111000001",
114193=>"000000000",
114194=>"100111000",
114195=>"010000001",
114196=>"000110010",
114197=>"011000111",
114198=>"000000111",
114199=>"011111101",
114200=>"010000000",
114201=>"000001111",
114202=>"111111100",
114203=>"000000000",
114204=>"010000000",
114205=>"111111101",
114206=>"001011100",
114207=>"011111000",
114208=>"000010000",
114209=>"000000000",
114210=>"101010101",
114211=>"101000010",
114212=>"111110111",
114213=>"011011011",
114214=>"011111110",
114215=>"000110000",
114216=>"000000001",
114217=>"000111101",
114218=>"100111001",
114219=>"000000000",
114220=>"111110000",
114221=>"010000000",
114222=>"111101101",
114223=>"000000000",
114224=>"010111100",
114225=>"110110111",
114226=>"100111101",
114227=>"111111101",
114228=>"111111000",
114229=>"010110000",
114230=>"000100100",
114231=>"111000001",
114232=>"101011100",
114233=>"110000110",
114234=>"000111010",
114235=>"000100111",
114236=>"111010000",
114237=>"111010001",
114238=>"000000000",
114239=>"000101110",
114240=>"101000000",
114241=>"001111101",
114242=>"110001001",
114243=>"000000001",
114244=>"000110110",
114245=>"000000000",
114246=>"010111000",
114247=>"000111111",
114248=>"010110110",
114249=>"000000010",
114250=>"000001000",
114251=>"000000000",
114252=>"101111000",
114253=>"100101111",
114254=>"001111111",
114255=>"101101101",
114256=>"111000000",
114257=>"001000111",
114258=>"000100101",
114259=>"000100000",
114260=>"010111111",
114261=>"011011011",
114262=>"100100010",
114263=>"000010111",
114264=>"000111011",
114265=>"011011110",
114266=>"100000000",
114267=>"010011001",
114268=>"111110111",
114269=>"000110100",
114270=>"000010010",
114271=>"000000000",
114272=>"111111111",
114273=>"110010000",
114274=>"111001111",
114275=>"001000011",
114276=>"000000110",
114277=>"111011000",
114278=>"110000000",
114279=>"111111000",
114280=>"010110111",
114281=>"011110111",
114282=>"111110000",
114283=>"110111111",
114284=>"000000011",
114285=>"111111001",
114286=>"000000000",
114287=>"000000000",
114288=>"100110110",
114289=>"000111100",
114290=>"100000001",
114291=>"110000000",
114292=>"011000001",
114293=>"111111110",
114294=>"000110100",
114295=>"111100000",
114296=>"000111111",
114297=>"000010110",
114298=>"001010001",
114299=>"010110110",
114300=>"001000100",
114301=>"111011111",
114302=>"000011101",
114303=>"000000000",
114304=>"101001010",
114305=>"000000001",
114306=>"111111110",
114307=>"111000110",
114308=>"101001000",
114309=>"100000000",
114310=>"100100110",
114311=>"110000000",
114312=>"000000111",
114313=>"011000000",
114314=>"111011011",
114315=>"000101110",
114316=>"000101001",
114317=>"111111111",
114318=>"000001110",
114319=>"110000110",
114320=>"111110000",
114321=>"010000000",
114322=>"111110000",
114323=>"001001000",
114324=>"010100000",
114325=>"101000000",
114326=>"111111111",
114327=>"010010000",
114328=>"010111111",
114329=>"011111101",
114330=>"011010111",
114331=>"101101000",
114332=>"111010000",
114333=>"000000100",
114334=>"101111111",
114335=>"101001000",
114336=>"010110110",
114337=>"000111101",
114338=>"110111000",
114339=>"101000000",
114340=>"111001111",
114341=>"100000110",
114342=>"000000000",
114343=>"000111000",
114344=>"000000000",
114345=>"000111111",
114346=>"111001011",
114347=>"101000000",
114348=>"101001000",
114349=>"111000011",
114350=>"101110010",
114351=>"111000000",
114352=>"000000000",
114353=>"111100000",
114354=>"000010111",
114355=>"101101011",
114356=>"010111111",
114357=>"010010000",
114358=>"010111111",
114359=>"111111000",
114360=>"110001110",
114361=>"001001000",
114362=>"010000101",
114363=>"101111111",
114364=>"111010110",
114365=>"001001111",
114366=>"100110011",
114367=>"110111010",
114368=>"000001111",
114369=>"111000001",
114370=>"001000110",
114371=>"111000101",
114372=>"000110111",
114373=>"111001011",
114374=>"000010001",
114375=>"000111111",
114376=>"000100101",
114377=>"000000010",
114378=>"000000111",
114379=>"000110110",
114380=>"110111001",
114381=>"100000011",
114382=>"000011011",
114383=>"111110010",
114384=>"111111001",
114385=>"111011110",
114386=>"000000010",
114387=>"111111011",
114388=>"000000000",
114389=>"011011001",
114390=>"000000110",
114391=>"110011111",
114392=>"110111000",
114393=>"111110000",
114394=>"000001111",
114395=>"000011000",
114396=>"000100010",
114397=>"111111101",
114398=>"000111111",
114399=>"111000000",
114400=>"101010010",
114401=>"100000000",
114402=>"111110000",
114403=>"000111011",
114404=>"110110101",
114405=>"010011000",
114406=>"111111001",
114407=>"101001111",
114408=>"111000111",
114409=>"001111110",
114410=>"011111100",
114411=>"001001111",
114412=>"111101111",
114413=>"011111101",
114414=>"011000011",
114415=>"000000000",
114416=>"000000000",
114417=>"011110100",
114418=>"101101000",
114419=>"100110000",
114420=>"111001000",
114421=>"010000000",
114422=>"010111111",
114423=>"111000101",
114424=>"000110110",
114425=>"000000001",
114426=>"000000100",
114427=>"010010010",
114428=>"111000111",
114429=>"011111000",
114430=>"011011111",
114431=>"111101001",
114432=>"000001000",
114433=>"011011010",
114434=>"100001110",
114435=>"111100110",
114436=>"111100100",
114437=>"111111011",
114438=>"000000110",
114439=>"001110110",
114440=>"111110111",
114441=>"011011000",
114442=>"000000110",
114443=>"110110100",
114444=>"011111111",
114445=>"111011000",
114446=>"111100000",
114447=>"100111101",
114448=>"001010010",
114449=>"100011111",
114450=>"110100001",
114451=>"100011011",
114452=>"100100001",
114453=>"000011011",
114454=>"010011011",
114455=>"111100100",
114456=>"000001100",
114457=>"011001111",
114458=>"011011010",
114459=>"011001011",
114460=>"001110011",
114461=>"000000010",
114462=>"011011000",
114463=>"000000100",
114464=>"100100001",
114465=>"000010100",
114466=>"110010001",
114467=>"000011011",
114468=>"110110100",
114469=>"100101101",
114470=>"011011010",
114471=>"111010111",
114472=>"100111100",
114473=>"100100100",
114474=>"011111011",
114475=>"011000001",
114476=>"001000001",
114477=>"111010111",
114478=>"011010101",
114479=>"100000100",
114480=>"011010001",
114481=>"100100100",
114482=>"001111101",
114483=>"011111001",
114484=>"000101001",
114485=>"001011000",
114486=>"011011010",
114487=>"011010011",
114488=>"011001000",
114489=>"001011000",
114490=>"100100100",
114491=>"011011111",
114492=>"100001101",
114493=>"100100101",
114494=>"001011011",
114495=>"111111101",
114496=>"001000011",
114497=>"111011011",
114498=>"110111011",
114499=>"000011110",
114500=>"101011011",
114501=>"110000000",
114502=>"000111111",
114503=>"110000111",
114504=>"110111111",
114505=>"100110111",
114506=>"101100011",
114507=>"001000111",
114508=>"111011011",
114509=>"101100100",
114510=>"100100101",
114511=>"100100111",
114512=>"110000110",
114513=>"000100100",
114514=>"010111111",
114515=>"001000011",
114516=>"110000000",
114517=>"001111101",
114518=>"100100100",
114519=>"000011000",
114520=>"111001000",
114521=>"111110011",
114522=>"101101101",
114523=>"000000111",
114524=>"011011011",
114525=>"001000000",
114526=>"011010011",
114527=>"011010011",
114528=>"011011011",
114529=>"011011011",
114530=>"100001011",
114531=>"111111000",
114532=>"100100101",
114533=>"001100101",
114534=>"000111000",
114535=>"101000000",
114536=>"011011000",
114537=>"010011001",
114538=>"110110111",
114539=>"110010101",
114540=>"111111101",
114541=>"100100101",
114542=>"000000001",
114543=>"000000011",
114544=>"001111110",
114545=>"011011111",
114546=>"000011011",
114547=>"110100111",
114548=>"011010111",
114549=>"000000011",
114550=>"011011010",
114551=>"011111011",
114552=>"111011000",
114553=>"110001111",
114554=>"100100100",
114555=>"001100100",
114556=>"111111101",
114557=>"110100000",
114558=>"000000101",
114559=>"011011110",
114560=>"110000000",
114561=>"111100100",
114562=>"011011011",
114563=>"011001101",
114564=>"111100110",
114565=>"111010101",
114566=>"101100101",
114567=>"101011000",
114568=>"101100100",
114569=>"101100111",
114570=>"111101111",
114571=>"111000011",
114572=>"110111110",
114573=>"001100100",
114574=>"111100101",
114575=>"001001010",
114576=>"110000100",
114577=>"110110011",
114578=>"000011110",
114579=>"011011000",
114580=>"110110110",
114581=>"001011011",
114582=>"111001011",
114583=>"111100100",
114584=>"000111100",
114585=>"110000000",
114586=>"100101100",
114587=>"000001001",
114588=>"011101011",
114589=>"000001001",
114590=>"011011011",
114591=>"100100001",
114592=>"100000000",
114593=>"011000000",
114594=>"100111100",
114595=>"100101011",
114596=>"101100101",
114597=>"100000001",
114598=>"100100100",
114599=>"011011011",
114600=>"011011011",
114601=>"001011111",
114602=>"100100100",
114603=>"000011001",
114604=>"100100001",
114605=>"010110110",
114606=>"110111101",
114607=>"000010111",
114608=>"010010000",
114609=>"000011011",
114610=>"100100100",
114611=>"100101101",
114612=>"100110101",
114613=>"111110110",
114614=>"011010111",
114615=>"100100000",
114616=>"001011011",
114617=>"001101101",
114618=>"111011101",
114619=>"101100110",
114620=>"100000001",
114621=>"100110111",
114622=>"001011000",
114623=>"011010110",
114624=>"110111010",
114625=>"011011011",
114626=>"011011111",
114627=>"111101111",
114628=>"000000100",
114629=>"111100000",
114630=>"011000000",
114631=>"100000111",
114632=>"101001000",
114633=>"011011100",
114634=>"111011000",
114635=>"001001011",
114636=>"011011010",
114637=>"000011001",
114638=>"011010000",
114639=>"110111100",
114640=>"100100100",
114641=>"100100111",
114642=>"011111100",
114643=>"100111101",
114644=>"000111000",
114645=>"101101111",
114646=>"110011001",
114647=>"111111001",
114648=>"010110111",
114649=>"000011011",
114650=>"101100111",
114651=>"100101111",
114652=>"111100111",
114653=>"001000110",
114654=>"011011111",
114655=>"110000110",
114656=>"100010011",
114657=>"110100111",
114658=>"000000100",
114659=>"110100111",
114660=>"010010011",
114661=>"110111110",
114662=>"110100011",
114663=>"000001010",
114664=>"001001111",
114665=>"011011111",
114666=>"001001001",
114667=>"101101000",
114668=>"000011010",
114669=>"000000111",
114670=>"000000000",
114671=>"100100001",
114672=>"111001001",
114673=>"000000011",
114674=>"011010000",
114675=>"100100111",
114676=>"111110000",
114677=>"001001001",
114678=>"101001001",
114679=>"001001001",
114680=>"001011010",
114681=>"110100100",
114682=>"011100100",
114683=>"111011011",
114684=>"001001101",
114685=>"110111111",
114686=>"011100001",
114687=>"111100101",
114688=>"100010111",
114689=>"000000001",
114690=>"111001001",
114691=>"001000110",
114692=>"101000011",
114693=>"100110111",
114694=>"111101000",
114695=>"000101000",
114696=>"000010111",
114697=>"111001110",
114698=>"001000100",
114699=>"110100000",
114700=>"110000000",
114701=>"010101001",
114702=>"001000010",
114703=>"000110111",
114704=>"110110000",
114705=>"111101000",
114706=>"111111000",
114707=>"111111100",
114708=>"111111111",
114709=>"101000000",
114710=>"000110111",
114711=>"111111000",
114712=>"111001000",
114713=>"001110100",
114714=>"000110111",
114715=>"010000011",
114716=>"111001101",
114717=>"101111001",
114718=>"111111111",
114719=>"101110110",
114720=>"000011111",
114721=>"100110111",
114722=>"000101100",
114723=>"000100110",
114724=>"100011001",
114725=>"011111110",
114726=>"110000000",
114727=>"101000111",
114728=>"001110110",
114729=>"000010110",
114730=>"011101000",
114731=>"000111110",
114732=>"000110101",
114733=>"101010000",
114734=>"000110001",
114735=>"001111001",
114736=>"111001010",
114737=>"000011011",
114738=>"101111000",
114739=>"010111001",
114740=>"111011101",
114741=>"111001100",
114742=>"000000110",
114743=>"011001001",
114744=>"011111111",
114745=>"111001001",
114746=>"111101100",
114747=>"000001101",
114748=>"000100010",
114749=>"111111011",
114750=>"100000000",
114751=>"000001111",
114752=>"000101000",
114753=>"000011100",
114754=>"000001001",
114755=>"100110111",
114756=>"010111111",
114757=>"100000001",
114758=>"111001000",
114759=>"000010110",
114760=>"100001110",
114761=>"000111111",
114762=>"111001001",
114763=>"110101000",
114764=>"000110010",
114765=>"000100100",
114766=>"000000100",
114767=>"001011101",
114768=>"111001010",
114769=>"010111101",
114770=>"111101001",
114771=>"000000001",
114772=>"111001000",
114773=>"101111110",
114774=>"111000001",
114775=>"111111000",
114776=>"111011100",
114777=>"100100100",
114778=>"111000000",
114779=>"100000011",
114780=>"001011000",
114781=>"001001011",
114782=>"101110111",
114783=>"001111111",
114784=>"000111111",
114785=>"000000111",
114786=>"110101001",
114787=>"111000000",
114788=>"000000101",
114789=>"011101110",
114790=>"100000001",
114791=>"111110010",
114792=>"000010011",
114793=>"111111000",
114794=>"011111101",
114795=>"000111111",
114796=>"000000010",
114797=>"111101000",
114798=>"111000000",
114799=>"101000101",
114800=>"000000010",
114801=>"001111001",
114802=>"000010011",
114803=>"110111000",
114804=>"010110101",
114805=>"111101100",
114806=>"000000000",
114807=>"000101111",
114808=>"111111000",
114809=>"111101000",
114810=>"100000110",
114811=>"101101111",
114812=>"100111110",
114813=>"000100100",
114814=>"100110111",
114815=>"100000110",
114816=>"100000000",
114817=>"010111100",
114818=>"000110000",
114819=>"000000000",
114820=>"000111111",
114821=>"111001001",
114822=>"100110110",
114823=>"100000100",
114824=>"000000001",
114825=>"111001001",
114826=>"110000100",
114827=>"110110110",
114828=>"000000110",
114829=>"101000100",
114830=>"110000000",
114831=>"111001001",
114832=>"010010011",
114833=>"000000111",
114834=>"000011110",
114835=>"000000000",
114836=>"011001011",
114837=>"101111000",
114838=>"111111111",
114839=>"000011011",
114840=>"101110010",
114841=>"000010010",
114842=>"111001001",
114843=>"101001001",
114844=>"110111101",
114845=>"111101000",
114846=>"111000001",
114847=>"111101000",
114848=>"011000100",
114849=>"010111000",
114850=>"000010110",
114851=>"101111010",
114852=>"111010010",
114853=>"010001000",
114854=>"000110110",
114855=>"000000111",
114856=>"000110111",
114857=>"000111101",
114858=>"111101000",
114859=>"111101001",
114860=>"000000000",
114861=>"000110111",
114862=>"111100100",
114863=>"111101001",
114864=>"010111111",
114865=>"010011101",
114866=>"110110110",
114867=>"001100110",
114868=>"000011111",
114869=>"110100000",
114870=>"000000100",
114871=>"111000111",
114872=>"000010111",
114873=>"000000111",
114874=>"000010000",
114875=>"000001000",
114876=>"110111101",
114877=>"111111111",
114878=>"000110110",
114879=>"000000000",
114880=>"111101101",
114881=>"010111000",
114882=>"000111011",
114883=>"111000011",
114884=>"111111101",
114885=>"000000001",
114886=>"000000111",
114887=>"111001000",
114888=>"010010000",
114889=>"011000010",
114890=>"001111110",
114891=>"111001000",
114892=>"000011011",
114893=>"100111111",
114894=>"111101101",
114895=>"000000011",
114896=>"111000000",
114897=>"000000110",
114898=>"001100110",
114899=>"010110111",
114900=>"111000000",
114901=>"110100110",
114902=>"110110111",
114903=>"010000001",
114904=>"000111101",
114905=>"000000110",
114906=>"100110000",
114907=>"111001000",
114908=>"000011101",
114909=>"001011111",
114910=>"110000000",
114911=>"111101001",
114912=>"001111111",
114913=>"111001100",
114914=>"001010000",
114915=>"011011011",
114916=>"111111000",
114917=>"000010110",
114918=>"000001001",
114919=>"010101100",
114920=>"000010000",
114921=>"000101010",
114922=>"000001001",
114923=>"010111100",
114924=>"000110111",
114925=>"000000000",
114926=>"000001001",
114927=>"111011110",
114928=>"110110111",
114929=>"000000100",
114930=>"111010011",
114931=>"000100100",
114932=>"000010110",
114933=>"111001000",
114934=>"000000100",
114935=>"000100000",
114936=>"000111111",
114937=>"000111001",
114938=>"010110000",
114939=>"100010111",
114940=>"111001000",
114941=>"000110111",
114942=>"101110110",
114943=>"111001000",
114944=>"110100110",
114945=>"000100100",
114946=>"010010000",
114947=>"000000000",
114948=>"110110100",
114949=>"000000000",
114950=>"111001101",
114951=>"010110100",
114952=>"000000000",
114953=>"000000101",
114954=>"101111010",
114955=>"101100111",
114956=>"000100100",
114957=>"011101000",
114958=>"100000000",
114959=>"000000000",
114960=>"010000000",
114961=>"111000011",
114962=>"011010111",
114963=>"001000000",
114964=>"000011000",
114965=>"111111011",
114966=>"010001000",
114967=>"110110111",
114968=>"111000100",
114969=>"111011110",
114970=>"111111111",
114971=>"000000000",
114972=>"000111011",
114973=>"000101111",
114974=>"001001011",
114975=>"010000000",
114976=>"001000000",
114977=>"110111111",
114978=>"000000101",
114979=>"000000000",
114980=>"010111110",
114981=>"001011011",
114982=>"111001000",
114983=>"101101111",
114984=>"111111111",
114985=>"000101100",
114986=>"000000000",
114987=>"000000100",
114988=>"110110110",
114989=>"110100001",
114990=>"111100010",
114991=>"110111111",
114992=>"110111111",
114993=>"010110000",
114994=>"000100111",
114995=>"011111011",
114996=>"111111111",
114997=>"000000000",
114998=>"111011001",
114999=>"101001000",
115000=>"010111100",
115001=>"001101101",
115002=>"000000100",
115003=>"110111010",
115004=>"111001001",
115005=>"111111111",
115006=>"010100000",
115007=>"000100001",
115008=>"000000100",
115009=>"001001111",
115010=>"111111000",
115011=>"100100000",
115012=>"101101000",
115013=>"000000111",
115014=>"000000000",
115015=>"000000100",
115016=>"000000100",
115017=>"000000000",
115018=>"010111111",
115019=>"110111011",
115020=>"000000000",
115021=>"000100010",
115022=>"110010010",
115023=>"010000010",
115024=>"101011010",
115025=>"010111111",
115026=>"001101010",
115027=>"001000000",
115028=>"000000000",
115029=>"010100111",
115030=>"011111101",
115031=>"001001111",
115032=>"001000000",
115033=>"111111110",
115034=>"011010000",
115035=>"111111110",
115036=>"111111111",
115037=>"011000000",
115038=>"111011010",
115039=>"111000000",
115040=>"000000000",
115041=>"001101011",
115042=>"000000000",
115043=>"110111000",
115044=>"000111010",
115045=>"000000000",
115046=>"101110000",
115047=>"000011000",
115048=>"000111000",
115049=>"000011111",
115050=>"001000100",
115051=>"110111011",
115052=>"110010011",
115053=>"010111111",
115054=>"000111000",
115055=>"000100100",
115056=>"111111111",
115057=>"000010001",
115058=>"110110100",
115059=>"000101010",
115060=>"000100011",
115061=>"000000100",
115062=>"111111000",
115063=>"000101101",
115064=>"000000000",
115065=>"100000000",
115066=>"100110111",
115067=>"111000111",
115068=>"010111001",
115069=>"100000001",
115070=>"111110011",
115071=>"000000000",
115072=>"000100000",
115073=>"001111010",
115074=>"000000111",
115075=>"110111111",
115076=>"011000000",
115077=>"000000000",
115078=>"110110110",
115079=>"110000000",
115080=>"000011011",
115081=>"111111111",
115082=>"100001001",
115083=>"000111111",
115084=>"010011001",
115085=>"100111001",
115086=>"110010011",
115087=>"000000000",
115088=>"000111101",
115089=>"111111011",
115090=>"000000100",
115091=>"011000001",
115092=>"110100100",
115093=>"000000000",
115094=>"101100100",
115095=>"000000010",
115096=>"100100101",
115097=>"010110001",
115098=>"000000000",
115099=>"000000000",
115100=>"001111111",
115101=>"110000000",
115102=>"000000111",
115103=>"101000000",
115104=>"100110111",
115105=>"010000110",
115106=>"001000000",
115107=>"000000000",
115108=>"111101001",
115109=>"100100010",
115110=>"111011100",
115111=>"010011011",
115112=>"110111110",
115113=>"100010100",
115114=>"000000010",
115115=>"000001100",
115116=>"111001111",
115117=>"100000000",
115118=>"001111111",
115119=>"001111001",
115120=>"111100000",
115121=>"000110011",
115122=>"101100101",
115123=>"000100000",
115124=>"001011110",
115125=>"001000000",
115126=>"100000100",
115127=>"111101100",
115128=>"110000100",
115129=>"010000000",
115130=>"111001111",
115131=>"100000010",
115132=>"000111011",
115133=>"100010110",
115134=>"000000000",
115135=>"011011111",
115136=>"011111011",
115137=>"111111111",
115138=>"101111111",
115139=>"000111110",
115140=>"000111111",
115141=>"111010010",
115142=>"000000100",
115143=>"111011011",
115144=>"100001111",
115145=>"100101101",
115146=>"111100100",
115147=>"101000001",
115148=>"000010000",
115149=>"001111100",
115150=>"111111010",
115151=>"110010011",
115152=>"011000100",
115153=>"100000000",
115154=>"001110000",
115155=>"000000000",
115156=>"111111111",
115157=>"001101110",
115158=>"101000000",
115159=>"000000111",
115160=>"011011011",
115161=>"000101011",
115162=>"100110111",
115163=>"000000101",
115164=>"010010011",
115165=>"000000101",
115166=>"111110011",
115167=>"101001000",
115168=>"110111111",
115169=>"000011011",
115170=>"000000001",
115171=>"011010000",
115172=>"101000011",
115173=>"000000000",
115174=>"100000000",
115175=>"110110110",
115176=>"000101000",
115177=>"000111011",
115178=>"011011011",
115179=>"111100110",
115180=>"000000000",
115181=>"000000110",
115182=>"001001111",
115183=>"110000000",
115184=>"101000110",
115185=>"100100010",
115186=>"101100100",
115187=>"110000000",
115188=>"001001011",
115189=>"010111011",
115190=>"000000000",
115191=>"110111011",
115192=>"010010010",
115193=>"011111101",
115194=>"000011000",
115195=>"000000000",
115196=>"000000000",
115197=>"101000101",
115198=>"010010000",
115199=>"111110000",
115200=>"010000001",
115201=>"011010001",
115202=>"111100111",
115203=>"000000000",
115204=>"000000000",
115205=>"100100001",
115206=>"001110111",
115207=>"000101000",
115208=>"000001110",
115209=>"111111111",
115210=>"111110100",
115211=>"000000001",
115212=>"000000000",
115213=>"010010000",
115214=>"110110000",
115215=>"111101000",
115216=>"001111111",
115217=>"000111000",
115218=>"111111111",
115219=>"000000100",
115220=>"000011011",
115221=>"000000000",
115222=>"000010000",
115223=>"111111000",
115224=>"000001000",
115225=>"011010110",
115226=>"001001101",
115227=>"111111101",
115228=>"111110011",
115229=>"000011000",
115230=>"000111000",
115231=>"010000000",
115232=>"000100101",
115233=>"000000000",
115234=>"101000000",
115235=>"111000110",
115236=>"011110101",
115237=>"010110100",
115238=>"100000000",
115239=>"101110111",
115240=>"001010000",
115241=>"000011010",
115242=>"111111111",
115243=>"100111101",
115244=>"000011011",
115245=>"010010000",
115246=>"110111001",
115247=>"111111111",
115248=>"000111010",
115249=>"111110110",
115250=>"011001001",
115251=>"111111101",
115252=>"010000100",
115253=>"000000110",
115254=>"111010000",
115255=>"111110111",
115256=>"111111111",
115257=>"111111010",
115258=>"111111011",
115259=>"111100101",
115260=>"010011011",
115261=>"111111111",
115262=>"000000000",
115263=>"010100000",
115264=>"111010000",
115265=>"101111001",
115266=>"011000000",
115267=>"000000000",
115268=>"101111000",
115269=>"101000000",
115270=>"111100001",
115271=>"111111111",
115272=>"011111110",
115273=>"101111111",
115274=>"111001111",
115275=>"010000000",
115276=>"111110101",
115277=>"111111011",
115278=>"101000110",
115279=>"001100011",
115280=>"000000000",
115281=>"111111111",
115282=>"000000010",
115283=>"010111000",
115284=>"010010110",
115285=>"111111000",
115286=>"111111111",
115287=>"101000101",
115288=>"111011001",
115289=>"111000000",
115290=>"110110010",
115291=>"000111110",
115292=>"111111100",
115293=>"111100100",
115294=>"011111111",
115295=>"000000000",
115296=>"110111111",
115297=>"111000000",
115298=>"111101100",
115299=>"011111010",
115300=>"000110010",
115301=>"010000000",
115302=>"111011111",
115303=>"000100101",
115304=>"000010010",
115305=>"110010000",
115306=>"011110000",
115307=>"110100001",
115308=>"010111010",
115309=>"111110010",
115310=>"000010100",
115311=>"000111001",
115312=>"110110001",
115313=>"000110110",
115314=>"100111000",
115315=>"010011011",
115316=>"100111111",
115317=>"000000011",
115318=>"111000000",
115319=>"111011111",
115320=>"101100011",
115321=>"111111010",
115322=>"010111111",
115323=>"001101001",
115324=>"101100111",
115325=>"111011000",
115326=>"100101111",
115327=>"111011010",
115328=>"010101001",
115329=>"000000000",
115330=>"011111000",
115331=>"000001011",
115332=>"000000000",
115333=>"010011011",
115334=>"100111000",
115335=>"000010110",
115336=>"011011000",
115337=>"101111001",
115338=>"100110011",
115339=>"111000001",
115340=>"000010111",
115341=>"000001001",
115342=>"101101111",
115343=>"000011011",
115344=>"010111100",
115345=>"110100000",
115346=>"001110111",
115347=>"110010000",
115348=>"000101100",
115349=>"100000000",
115350=>"000000000",
115351=>"101100100",
115352=>"110110011",
115353=>"010111101",
115354=>"111110000",
115355=>"111001000",
115356=>"000110100",
115357=>"111111111",
115358=>"101010111",
115359=>"000010000",
115360=>"011111011",
115361=>"000111000",
115362=>"111111001",
115363=>"000100010",
115364=>"110110000",
115365=>"000010000",
115366=>"101011001",
115367=>"000111000",
115368=>"011010111",
115369=>"010000001",
115370=>"111011101",
115371=>"100111100",
115372=>"011111101",
115373=>"111100111",
115374=>"110111100",
115375=>"000010000",
115376=>"111101111",
115377=>"000010001",
115378=>"111111111",
115379=>"111001011",
115380=>"000100100",
115381=>"111111010",
115382=>"000000010",
115383=>"111110101",
115384=>"011011110",
115385=>"000110100",
115386=>"111111110",
115387=>"000000111",
115388=>"000110001",
115389=>"111111111",
115390=>"000010011",
115391=>"010110111",
115392=>"011111010",
115393=>"000100111",
115394=>"111011001",
115395=>"111100000",
115396=>"101000111",
115397=>"111001001",
115398=>"111101001",
115399=>"111111111",
115400=>"011011000",
115401=>"000000000",
115402=>"001000111",
115403=>"010001110",
115404=>"000000000",
115405=>"001011110",
115406=>"010100111",
115407=>"000000101",
115408=>"111111110",
115409=>"000010010",
115410=>"000000000",
115411=>"110101011",
115412=>"011011100",
115413=>"101000000",
115414=>"111111000",
115415=>"000000111",
115416=>"000000010",
115417=>"110011110",
115418=>"110110111",
115419=>"110111110",
115420=>"000111100",
115421=>"110111111",
115422=>"000111111",
115423=>"110111110",
115424=>"110000011",
115425=>"110010000",
115426=>"111010100",
115427=>"100010000",
115428=>"000000000",
115429=>"000000000",
115430=>"101100000",
115431=>"010011000",
115432=>"000000000",
115433=>"000110010",
115434=>"111011000",
115435=>"010001000",
115436=>"111000100",
115437=>"010001100",
115438=>"111111111",
115439=>"011111111",
115440=>"000000000",
115441=>"101100001",
115442=>"100111101",
115443=>"011011110",
115444=>"011011000",
115445=>"111110000",
115446=>"111111111",
115447=>"001000101",
115448=>"000111111",
115449=>"011110011",
115450=>"111111111",
115451=>"100000000",
115452=>"111111111",
115453=>"011001000",
115454=>"111111100",
115455=>"001110110",
115456=>"011010000",
115457=>"000000010",
115458=>"110111111",
115459=>"010010000",
115460=>"100110110",
115461=>"000110111",
115462=>"010111000",
115463=>"111000000",
115464=>"000000000",
115465=>"000000000",
115466=>"000000000",
115467=>"010010000",
115468=>"000111000",
115469=>"000010000",
115470=>"101101101",
115471=>"111111111",
115472=>"000000000",
115473=>"011110000",
115474=>"010100100",
115475=>"000000000",
115476=>"100001000",
115477=>"011111011",
115478=>"111111111",
115479=>"111000000",
115480=>"000100000",
115481=>"001111111",
115482=>"101000000",
115483=>"111110111",
115484=>"011111101",
115485=>"010011011",
115486=>"111110100",
115487=>"010100000",
115488=>"011110000",
115489=>"000110000",
115490=>"111100100",
115491=>"111000000",
115492=>"011001011",
115493=>"111111001",
115494=>"011011000",
115495=>"101000110",
115496=>"000000000",
115497=>"000000001",
115498=>"000010110",
115499=>"111100111",
115500=>"100011000",
115501=>"100010000",
115502=>"111101111",
115503=>"111110111",
115504=>"000000000",
115505=>"100100100",
115506=>"011000011",
115507=>"111111101",
115508=>"000000110",
115509=>"000111000",
115510=>"001011011",
115511=>"010000101",
115512=>"111111000",
115513=>"111001101",
115514=>"000001000",
115515=>"000000000",
115516=>"111110101",
115517=>"101111111",
115518=>"010000000",
115519=>"000100000",
115520=>"110000100",
115521=>"110010110",
115522=>"011100000",
115523=>"001100110",
115524=>"010111111",
115525=>"000001111",
115526=>"010010010",
115527=>"000101111",
115528=>"010000000",
115529=>"101000001",
115530=>"000000111",
115531=>"000000000",
115532=>"101000101",
115533=>"110111111",
115534=>"101111001",
115535=>"111111111",
115536=>"111111011",
115537=>"000110111",
115538=>"010111010",
115539=>"001111001",
115540=>"000100100",
115541=>"001010010",
115542=>"110100111",
115543=>"100000000",
115544=>"000000000",
115545=>"110110100",
115546=>"001011001",
115547=>"100100000",
115548=>"010011000",
115549=>"011001001",
115550=>"111111111",
115551=>"100001011",
115552=>"000000110",
115553=>"111000111",
115554=>"000000000",
115555=>"011011110",
115556=>"010111101",
115557=>"100100000",
115558=>"000110000",
115559=>"110110000",
115560=>"010111000",
115561=>"111101100",
115562=>"111100000",
115563=>"000000000",
115564=>"111100101",
115565=>"000000000",
115566=>"010111011",
115567=>"111111111",
115568=>"000110110",
115569=>"111011000",
115570=>"100110000",
115571=>"111000111",
115572=>"000000111",
115573=>"111010101",
115574=>"111111000",
115575=>"000100110",
115576=>"110110100",
115577=>"111011000",
115578=>"000100001",
115579=>"111111111",
115580=>"110110111",
115581=>"100100000",
115582=>"000000001",
115583=>"001011011",
115584=>"100111111",
115585=>"111110100",
115586=>"000000001",
115587=>"100111111",
115588=>"111111100",
115589=>"000000000",
115590=>"110100100",
115591=>"110010111",
115592=>"001011111",
115593=>"000101111",
115594=>"000000000",
115595=>"111111111",
115596=>"000011111",
115597=>"000111010",
115598=>"111111111",
115599=>"111000001",
115600=>"010100100",
115601=>"110110110",
115602=>"100000000",
115603=>"111100011",
115604=>"111001100",
115605=>"010111111",
115606=>"000111110",
115607=>"000000001",
115608=>"011011011",
115609=>"111011101",
115610=>"110111011",
115611=>"000000000",
115612=>"000011001",
115613=>"010111111",
115614=>"000000000",
115615=>"101000111",
115616=>"110110100",
115617=>"111110011",
115618=>"111111010",
115619=>"100101111",
115620=>"000000000",
115621=>"101011000",
115622=>"101001001",
115623=>"000011011",
115624=>"110100111",
115625=>"111111000",
115626=>"000000000",
115627=>"011101111",
115628=>"110100000",
115629=>"111111111",
115630=>"111111011",
115631=>"000001101",
115632=>"111100111",
115633=>"001000100",
115634=>"111001111",
115635=>"110110010",
115636=>"000101000",
115637=>"011100000",
115638=>"111110110",
115639=>"010111110",
115640=>"000011100",
115641=>"101101001",
115642=>"000000010",
115643=>"010110111",
115644=>"111111111",
115645=>"111111111",
115646=>"000000000",
115647=>"111111111",
115648=>"010010000",
115649=>"000000110",
115650=>"111000001",
115651=>"001001001",
115652=>"000000001",
115653=>"000111011",
115654=>"110100001",
115655=>"000000100",
115656=>"111001111",
115657=>"001000000",
115658=>"011111010",
115659=>"010111110",
115660=>"100110111",
115661=>"001011011",
115662=>"110000000",
115663=>"100000000",
115664=>"111100100",
115665=>"000100100",
115666=>"101101111",
115667=>"000101111",
115668=>"101000101",
115669=>"110110000",
115670=>"110110000",
115671=>"100000000",
115672=>"100000000",
115673=>"011111011",
115674=>"101000001",
115675=>"101100100",
115676=>"101110101",
115677=>"000001000",
115678=>"000011111",
115679=>"110011000",
115680=>"000000001",
115681=>"011111101",
115682=>"000000000",
115683=>"001101101",
115684=>"101000000",
115685=>"010110110",
115686=>"000110010",
115687=>"100110010",
115688=>"000100000",
115689=>"011100110",
115690=>"111111000",
115691=>"111000000",
115692=>"000010000",
115693=>"101000001",
115694=>"111111111",
115695=>"101000000",
115696=>"000000000",
115697=>"110011111",
115698=>"111000000",
115699=>"110111010",
115700=>"111000001",
115701=>"001111101",
115702=>"000000010",
115703=>"111101100",
115704=>"111111110",
115705=>"001111000",
115706=>"000111111",
115707=>"111100001",
115708=>"111111111",
115709=>"010111010",
115710=>"010100000",
115711=>"110100110",
115712=>"000000111",
115713=>"000000100",
115714=>"101000100",
115715=>"000000000",
115716=>"100100100",
115717=>"111000000",
115718=>"101001111",
115719=>"100100000",
115720=>"000000111",
115721=>"110000101",
115722=>"000001001",
115723=>"010011000",
115724=>"001010010",
115725=>"111101000",
115726=>"100100010",
115727=>"101011111",
115728=>"101000100",
115729=>"111000101",
115730=>"010101100",
115731=>"000100000",
115732=>"001110111",
115733=>"111011101",
115734=>"000000110",
115735=>"101101001",
115736=>"111100000",
115737=>"000000000",
115738=>"001101111",
115739=>"111111111",
115740=>"111011100",
115741=>"000100101",
115742=>"100101101",
115743=>"000111111",
115744=>"100101111",
115745=>"011111000",
115746=>"100010111",
115747=>"000011110",
115748=>"010111011",
115749=>"001100001",
115750=>"101000111",
115751=>"000000011",
115752=>"000011111",
115753=>"001110111",
115754=>"100101101",
115755=>"110011110",
115756=>"011000110",
115757=>"111010010",
115758=>"011101101",
115759=>"010111101",
115760=>"011110111",
115761=>"000011010",
115762=>"010000010",
115763=>"110111111",
115764=>"111000000",
115765=>"101010111",
115766=>"110100000",
115767=>"011000100",
115768=>"111111100",
115769=>"101000000",
115770=>"011010011",
115771=>"100011011",
115772=>"100000100",
115773=>"111111111",
115774=>"000100000",
115775=>"000011001",
115776=>"000000111",
115777=>"001001011",
115778=>"101111111",
115779=>"000100101",
115780=>"000011011",
115781=>"101000000",
115782=>"101101101",
115783=>"111111000",
115784=>"111100000",
115785=>"110101101",
115786=>"000000000",
115787=>"111111101",
115788=>"011100101",
115789=>"000101110",
115790=>"000100011",
115791=>"111111100",
115792=>"111000000",
115793=>"011010000",
115794=>"011010000",
115795=>"010011001",
115796=>"111000001",
115797=>"001111100",
115798=>"101000010",
115799=>"111000100",
115800=>"011111011",
115801=>"011001000",
115802=>"100100110",
115803=>"000011011",
115804=>"000101010",
115805=>"100001001",
115806=>"111011111",
115807=>"100000111",
115808=>"000010101",
115809=>"010101000",
115810=>"111000100",
115811=>"001001001",
115812=>"000011010",
115813=>"011000000",
115814=>"010101011",
115815=>"100010011",
115816=>"000010010",
115817=>"111000000",
115818=>"010111101",
115819=>"111000010",
115820=>"000100111",
115821=>"111101111",
115822=>"010000101",
115823=>"111010000",
115824=>"001000110",
115825=>"111000000",
115826=>"011001000",
115827=>"100001011",
115828=>"111001000",
115829=>"011000100",
115830=>"111000000",
115831=>"000000111",
115832=>"011000101",
115833=>"111010100",
115834=>"000111111",
115835=>"000110001",
115836=>"000110000",
115837=>"000000100",
115838=>"000010000",
115839=>"101101000",
115840=>"001101101",
115841=>"111101101",
115842=>"001000110",
115843=>"000000000",
115844=>"010011001",
115845=>"000001111",
115846=>"100111100",
115847=>"100000001",
115848=>"110111011",
115849=>"000000010",
115850=>"000100100",
115851=>"100010000",
115852=>"000110111",
115853=>"000100010",
115854=>"000101010",
115855=>"001000000",
115856=>"010100010",
115857=>"000110011",
115858=>"011001000",
115859=>"111101000",
115860=>"000100111",
115861=>"111000000",
115862=>"111110111",
115863=>"000001011",
115864=>"111110010",
115865=>"000000000",
115866=>"000000000",
115867=>"001011100",
115868=>"100100111",
115869=>"010101111",
115870=>"101111000",
115871=>"110110100",
115872=>"001101010",
115873=>"011000101",
115874=>"000000101",
115875=>"001000111",
115876=>"010000101",
115877=>"100000011",
115878=>"000110110",
115879=>"110101111",
115880=>"111100000",
115881=>"100000110",
115882=>"101111101",
115883=>"111100000",
115884=>"000001010",
115885=>"001101000",
115886=>"110001001",
115887=>"000010010",
115888=>"000011100",
115889=>"010011101",
115890=>"000000010",
115891=>"010010110",
115892=>"101011011",
115893=>"011111010",
115894=>"001000001",
115895=>"000000000",
115896=>"001000001",
115897=>"000001001",
115898=>"000000001",
115899=>"010111011",
115900=>"010010011",
115901=>"101000110",
115902=>"001100010",
115903=>"011010111",
115904=>"111000001",
115905=>"100000100",
115906=>"111000100",
115907=>"101101111",
115908=>"100000100",
115909=>"110110011",
115910=>"110110110",
115911=>"010000111",
115912=>"110000000",
115913=>"101010111",
115914=>"100100111",
115915=>"111011111",
115916=>"000100100",
115917=>"000001000",
115918=>"000000000",
115919=>"100010011",
115920=>"111010000",
115921=>"100100111",
115922=>"000000010",
115923=>"000101111",
115924=>"101111111",
115925=>"110110000",
115926=>"111111100",
115927=>"101100100",
115928=>"010010000",
115929=>"010010111",
115930=>"000100001",
115931=>"111100101",
115932=>"000010001",
115933=>"101001101",
115934=>"000011111",
115935=>"111101101",
115936=>"011110110",
115937=>"111101000",
115938=>"101011011",
115939=>"000001011",
115940=>"100000101",
115941=>"000111010",
115942=>"000010011",
115943=>"011100100",
115944=>"110101101",
115945=>"000000111",
115946=>"000100100",
115947=>"011100000",
115948=>"000010010",
115949=>"010010001",
115950=>"100000000",
115951=>"100100101",
115952=>"010111010",
115953=>"011011100",
115954=>"000000101",
115955=>"000110110",
115956=>"001101100",
115957=>"001001000",
115958=>"100101101",
115959=>"100001111",
115960=>"111000000",
115961=>"111110101",
115962=>"011111101",
115963=>"101111111",
115964=>"111101111",
115965=>"000011011",
115966=>"000100011",
115967=>"111100100",
115968=>"001100010",
115969=>"001011000",
115970=>"100000110",
115971=>"001010111",
115972=>"000000010",
115973=>"100000000",
115974=>"001001010",
115975=>"111000001",
115976=>"010100110",
115977=>"110010100",
115978=>"001011001",
115979=>"100110100",
115980=>"110100100",
115981=>"000000000",
115982=>"100001101",
115983=>"001010000",
115984=>"010000000",
115985=>"111111000",
115986=>"000100001",
115987=>"100100110",
115988=>"011001001",
115989=>"011110110",
115990=>"011101000",
115991=>"100111000",
115992=>"001000000",
115993=>"000000011",
115994=>"100001001",
115995=>"110111111",
115996=>"111011011",
115997=>"011000000",
115998=>"110110111",
115999=>"100111011",
116000=>"100100110",
116001=>"111101001",
116002=>"001001000",
116003=>"011111101",
116004=>"010001000",
116005=>"001000100",
116006=>"000100000",
116007=>"111010011",
116008=>"111110100",
116009=>"011011001",
116010=>"000000010",
116011=>"000111011",
116012=>"000001011",
116013=>"011111100",
116014=>"111001101",
116015=>"100101000",
116016=>"111110100",
116017=>"011001011",
116018=>"111000111",
116019=>"100001010",
116020=>"010001000",
116021=>"010010000",
116022=>"010011010",
116023=>"110001100",
116024=>"100100111",
116025=>"110100000",
116026=>"000110111",
116027=>"111110111",
116028=>"010110100",
116029=>"111011001",
116030=>"001000000",
116031=>"000111110",
116032=>"110110111",
116033=>"001001011",
116034=>"100100100",
116035=>"100110010",
116036=>"000011000",
116037=>"100110101",
116038=>"011111110",
116039=>"011100100",
116040=>"011101010",
116041=>"011010110",
116042=>"111110110",
116043=>"011100110",
116044=>"111101110",
116045=>"111011000",
116046=>"000110111",
116047=>"000101000",
116048=>"100011011",
116049=>"011101011",
116050=>"001100000",
116051=>"111010000",
116052=>"010011001",
116053=>"011000011",
116054=>"001001001",
116055=>"110110101",
116056=>"000111011",
116057=>"011011111",
116058=>"010001001",
116059=>"001011111",
116060=>"010000100",
116061=>"000001000",
116062=>"111110111",
116063=>"111111010",
116064=>"111011010",
116065=>"001001100",
116066=>"000100111",
116067=>"001011011",
116068=>"100100111",
116069=>"111111111",
116070=>"110100111",
116071=>"100000000",
116072=>"000110111",
116073=>"110000101",
116074=>"011110100",
116075=>"010010000",
116076=>"111101001",
116077=>"001001000",
116078=>"000001000",
116079=>"011111000",
116080=>"010001001",
116081=>"111110001",
116082=>"110000001",
116083=>"011010000",
116084=>"000001000",
116085=>"110100110",
116086=>"000011010",
116087=>"000000111",
116088=>"100100100",
116089=>"011011001",
116090=>"100101011",
116091=>"010100110",
116092=>"001001000",
116093=>"110100110",
116094=>"100110110",
116095=>"110110110",
116096=>"111110000",
116097=>"100100011",
116098=>"011011111",
116099=>"001001011",
116100=>"011100001",
116101=>"001000000",
116102=>"011111000",
116103=>"100000011",
116104=>"000001111",
116105=>"100110001",
116106=>"000010000",
116107=>"100111001",
116108=>"010110010",
116109=>"110110010",
116110=>"000010111",
116111=>"000000000",
116112=>"001001000",
116113=>"000110100",
116114=>"000110110",
116115=>"000110000",
116116=>"001101101",
116117=>"010100100",
116118=>"011011111",
116119=>"100110010",
116120=>"110111111",
116121=>"010100000",
116122=>"000100110",
116123=>"000110100",
116124=>"111100000",
116125=>"000111010",
116126=>"001101111",
116127=>"111100110",
116128=>"011100011",
116129=>"010000011",
116130=>"100100111",
116131=>"000100101",
116132=>"001010011",
116133=>"110011110",
116134=>"000100001",
116135=>"010000000",
116136=>"001011000",
116137=>"000110110",
116138=>"000100110",
116139=>"110111011",
116140=>"111000011",
116141=>"110000101",
116142=>"000011011",
116143=>"000100110",
116144=>"100110100",
116145=>"110110001",
116146=>"001111011",
116147=>"110100000",
116148=>"101001000",
116149=>"000001000",
116150=>"001001001",
116151=>"110001000",
116152=>"011000000",
116153=>"001100010",
116154=>"011100100",
116155=>"100100100",
116156=>"000000111",
116157=>"011111001",
116158=>"100100111",
116159=>"111110000",
116160=>"100000100",
116161=>"001011000",
116162=>"001110000",
116163=>"111001001",
116164=>"000000101",
116165=>"001001110",
116166=>"111100000",
116167=>"000100110",
116168=>"110100110",
116169=>"100001001",
116170=>"100111011",
116171=>"000110010",
116172=>"110110111",
116173=>"111101100",
116174=>"000011001",
116175=>"000100110",
116176=>"100011001",
116177=>"010011001",
116178=>"000100000",
116179=>"111011000",
116180=>"010001001",
116181=>"000011101",
116182=>"001001001",
116183=>"100011000",
116184=>"111000011",
116185=>"000000000",
116186=>"000110101",
116187=>"110100100",
116188=>"011010111",
116189=>"100100100",
116190=>"011001000",
116191=>"000100010",
116192=>"100100100",
116193=>"111011001",
116194=>"010110110",
116195=>"010010110",
116196=>"110000000",
116197=>"011010011",
116198=>"000000000",
116199=>"000011011",
116200=>"110010000",
116201=>"000001001",
116202=>"111011011",
116203=>"010110110",
116204=>"100100100",
116205=>"111001001",
116206=>"110100100",
116207=>"011100100",
116208=>"100100110",
116209=>"011011000",
116210=>"111110110",
116211=>"011011001",
116212=>"101111100",
116213=>"100011001",
116214=>"000000100",
116215=>"000000000",
116216=>"000100010",
116217=>"111100110",
116218=>"111111110",
116219=>"111111001",
116220=>"010110000",
116221=>"011000010",
116222=>"001011111",
116223=>"011011110",
116224=>"101111110",
116225=>"000000000",
116226=>"101001000",
116227=>"000000001",
116228=>"000100110",
116229=>"111101111",
116230=>"101110110",
116231=>"100100000",
116232=>"101001000",
116233=>"001000000",
116234=>"011111011",
116235=>"001011111",
116236=>"001100111",
116237=>"111100101",
116238=>"110000110",
116239=>"111111010",
116240=>"000000010",
116241=>"000000000",
116242=>"001101101",
116243=>"010110111",
116244=>"010110101",
116245=>"111000111",
116246=>"001101000",
116247=>"111111000",
116248=>"010000010",
116249=>"000000000",
116250=>"100101111",
116251=>"000000101",
116252=>"100010000",
116253=>"011110101",
116254=>"111101000",
116255=>"000000111",
116256=>"110001000",
116257=>"000010000",
116258=>"000101111",
116259=>"000000111",
116260=>"011100111",
116261=>"111001111",
116262=>"000000011",
116263=>"000110000",
116264=>"011010011",
116265=>"100111111",
116266=>"110010010",
116267=>"000010000",
116268=>"011100001",
116269=>"111100111",
116270=>"111111111",
116271=>"110000111",
116272=>"111101001",
116273=>"100111010",
116274=>"000001000",
116275=>"111111111",
116276=>"000011111",
116277=>"001000011",
116278=>"000000011",
116279=>"000110100",
116280=>"111101001",
116281=>"001001111",
116282=>"001111101",
116283=>"010000110",
116284=>"000011111",
116285=>"011110110",
116286=>"101000000",
116287=>"101001100",
116288=>"100000000",
116289=>"000010101",
116290=>"101101000",
116291=>"001101101",
116292=>"100111111",
116293=>"101101001",
116294=>"111010010",
116295=>"111101111",
116296=>"110001100",
116297=>"000100000",
116298=>"000101101",
116299=>"111010110",
116300=>"101101111",
116301=>"111111111",
116302=>"000011010",
116303=>"100100001",
116304=>"000000010",
116305=>"111010000",
116306=>"010010111",
116307=>"011001000",
116308=>"000000110",
116309=>"001001000",
116310=>"010010111",
116311=>"000000000",
116312=>"101111011",
116313=>"000101111",
116314=>"100001011",
116315=>"000001111",
116316=>"110111010",
116317=>"100000001",
116318=>"110010111",
116319=>"100100111",
116320=>"100101111",
116321=>"001000100",
116322=>"111000111",
116323=>"011100100",
116324=>"011111110",
116325=>"111010010",
116326=>"001001111",
116327=>"101111111",
116328=>"000101111",
116329=>"111110001",
116330=>"101110010",
116331=>"001111010",
116332=>"010000101",
116333=>"111111100",
116334=>"001100100",
116335=>"111111100",
116336=>"100100100",
116337=>"000110010",
116338=>"100000000",
116339=>"111100000",
116340=>"110111110",
116341=>"101000101",
116342=>"111011000",
116343=>"000001111",
116344=>"000000101",
116345=>"000111111",
116346=>"111111111",
116347=>"111101000",
116348=>"000001000",
116349=>"111101000",
116350=>"101111111",
116351=>"001001101",
116352=>"010010001",
116353=>"100100101",
116354=>"000110111",
116355=>"000010010",
116356=>"111000110",
116357=>"010110111",
116358=>"110110101",
116359=>"000100000",
116360=>"001001001",
116361=>"000010110",
116362=>"111010000",
116363=>"000011000",
116364=>"000001000",
116365=>"101101111",
116366=>"000010000",
116367=>"000000011",
116368=>"001111111",
116369=>"111101110",
116370=>"111010000",
116371=>"100000001",
116372=>"000000010",
116373=>"000111111",
116374=>"110110010",
116375=>"100100110",
116376=>"001001001",
116377=>"000000000",
116378=>"110111011",
116379=>"100000000",
116380=>"101111000",
116381=>"000000000",
116382=>"010111000",
116383=>"001101000",
116384=>"001000000",
116385=>"010001000",
116386=>"000000000",
116387=>"000000000",
116388=>"111111011",
116389=>"111111111",
116390=>"001111001",
116391=>"000100001",
116392=>"011011011",
116393=>"111001000",
116394=>"111000000",
116395=>"000000100",
116396=>"000001000",
116397=>"001001111",
116398=>"011011010",
116399=>"001000110",
116400=>"000100101",
116401=>"000001011",
116402=>"000001100",
116403=>"000101011",
116404=>"111111011",
116405=>"011011011",
116406=>"011100111",
116407=>"111011000",
116408=>"000110111",
116409=>"000001000",
116410=>"110111111",
116411=>"110100111",
116412=>"010000111",
116413=>"100001000",
116414=>"100000000",
116415=>"000000000",
116416=>"111000100",
116417=>"000011010",
116418=>"110111111",
116419=>"001100110",
116420=>"111111111",
116421=>"111110001",
116422=>"111111000",
116423=>"111111000",
116424=>"000110011",
116425=>"000000101",
116426=>"000111011",
116427=>"000010000",
116428=>"000110111",
116429=>"000100000",
116430=>"000000010",
116431=>"100100000",
116432=>"000011111",
116433=>"011001001",
116434=>"100000010",
116435=>"111111111",
116436=>"000000111",
116437=>"000000100",
116438=>"101100101",
116439=>"010110000",
116440=>"011011001",
116441=>"000111111",
116442=>"000001000",
116443=>"111011000",
116444=>"001000000",
116445=>"000101110",
116446=>"100101011",
116447=>"110110000",
116448=>"000000101",
116449=>"111000000",
116450=>"111110111",
116451=>"100100100",
116452=>"000000000",
116453=>"010111110",
116454=>"101011010",
116455=>"010010110",
116456=>"000111111",
116457=>"010111110",
116458=>"110011000",
116459=>"100000010",
116460=>"000101111",
116461=>"111011011",
116462=>"101001000",
116463=>"100001111",
116464=>"000000011",
116465=>"111011101",
116466=>"001100101",
116467=>"101101101",
116468=>"011011111",
116469=>"000101111",
116470=>"101011111",
116471=>"001001101",
116472=>"010000000",
116473=>"110111101",
116474=>"101101111",
116475=>"010111111",
116476=>"111111011",
116477=>"001111110",
116478=>"100011110",
116479=>"000000000",
116480=>"100000110",
116481=>"000000000",
116482=>"100111111",
116483=>"100000000",
116484=>"001100100",
116485=>"011000011",
116486=>"111111111",
116487=>"001101101",
116488=>"000100100",
116489=>"000111000",
116490=>"001001011",
116491=>"001101111",
116492=>"010000000",
116493=>"110000000",
116494=>"110100100",
116495=>"111111111",
116496=>"011000111",
116497=>"101111111",
116498=>"011011011",
116499=>"000000000",
116500=>"000000000",
116501=>"001010111",
116502=>"110011111",
116503=>"111111000",
116504=>"001000000",
116505=>"010000010",
116506=>"100100101",
116507=>"111111111",
116508=>"000001100",
116509=>"101111011",
116510=>"000010011",
116511=>"101101000",
116512=>"000011010",
116513=>"111000111",
116514=>"110111101",
116515=>"001111111",
116516=>"011011010",
116517=>"001000010",
116518=>"000010010",
116519=>"111111011",
116520=>"011000000",
116521=>"100100100",
116522=>"010000110",
116523=>"000011010",
116524=>"111011011",
116525=>"000000001",
116526=>"000111111",
116527=>"110111111",
116528=>"111111000",
116529=>"110110111",
116530=>"010001101",
116531=>"010011011",
116532=>"111111111",
116533=>"111100110",
116534=>"011111111",
116535=>"111101101",
116536=>"000000000",
116537=>"001111100",
116538=>"111111111",
116539=>"111111111",
116540=>"001011101",
116541=>"111111000",
116542=>"000000000",
116543=>"010100101",
116544=>"111100111",
116545=>"010010010",
116546=>"001010000",
116547=>"000000100",
116548=>"111000011",
116549=>"000000100",
116550=>"110000000",
116551=>"100111111",
116552=>"000000000",
116553=>"101000111",
116554=>"100101001",
116555=>"110000000",
116556=>"000111111",
116557=>"100100100",
116558=>"001001011",
116559=>"000000101",
116560=>"000111011",
116561=>"111111111",
116562=>"101000100",
116563=>"001100111",
116564=>"000100000",
116565=>"111101111",
116566=>"111011001",
116567=>"000100110",
116568=>"001111111",
116569=>"110110110",
116570=>"111101100",
116571=>"011011111",
116572=>"001111100",
116573=>"000110110",
116574=>"011000111",
116575=>"000100011",
116576=>"000000000",
116577=>"000000000",
116578=>"010000010",
116579=>"111011000",
116580=>"101011111",
116581=>"111000100",
116582=>"000000000",
116583=>"101100000",
116584=>"111000000",
116585=>"010010111",
116586=>"000000010",
116587=>"000100001",
116588=>"001000000",
116589=>"011111111",
116590=>"101000100",
116591=>"111000101",
116592=>"100100100",
116593=>"010010000",
116594=>"110011011",
116595=>"111111001",
116596=>"000100000",
116597=>"001111001",
116598=>"001000100",
116599=>"111111111",
116600=>"001000111",
116601=>"000111010",
116602=>"110100001",
116603=>"111111111",
116604=>"100011111",
116605=>"010001111",
116606=>"110001111",
116607=>"000000000",
116608=>"010000001",
116609=>"100100000",
116610=>"010110111",
116611=>"111111101",
116612=>"101000000",
116613=>"111000100",
116614=>"110010000",
116615=>"101110110",
116616=>"001000001",
116617=>"001100010",
116618=>"111000010",
116619=>"100010010",
116620=>"000000000",
116621=>"010001011",
116622=>"000111111",
116623=>"001001101",
116624=>"111011000",
116625=>"111000000",
116626=>"011000100",
116627=>"111000000",
116628=>"000000000",
116629=>"111001101",
116630=>"011111111",
116631=>"001001000",
116632=>"110101100",
116633=>"100001111",
116634=>"111111101",
116635=>"101000000",
116636=>"000110100",
116637=>"010000111",
116638=>"001000111",
116639=>"000011000",
116640=>"100111111",
116641=>"011111011",
116642=>"111000000",
116643=>"110111101",
116644=>"111000000",
116645=>"110110110",
116646=>"000001001",
116647=>"011001100",
116648=>"000000010",
116649=>"111111001",
116650=>"010001100",
116651=>"001101111",
116652=>"111000001",
116653=>"000000000",
116654=>"001101111",
116655=>"001000000",
116656=>"001101101",
116657=>"000001100",
116658=>"010011011",
116659=>"000011011",
116660=>"111000001",
116661=>"000100001",
116662=>"011011010",
116663=>"111000000",
116664=>"110110110",
116665=>"001000100",
116666=>"000000000",
116667=>"000101100",
116668=>"000110111",
116669=>"001011011",
116670=>"110010101",
116671=>"000111000",
116672=>"000000111",
116673=>"000011000",
116674=>"000000000",
116675=>"100110110",
116676=>"111111110",
116677=>"000000001",
116678=>"111111000",
116679=>"000100111",
116680=>"101111111",
116681=>"000101100",
116682=>"000000000",
116683=>"010010111",
116684=>"000000111",
116685=>"011110110",
116686=>"111111000",
116687=>"010011111",
116688=>"011000000",
116689=>"011000000",
116690=>"111000100",
116691=>"111101110",
116692=>"000111111",
116693=>"010000000",
116694=>"001111111",
116695=>"000000000",
116696=>"011000000",
116697=>"111000000",
116698=>"000010111",
116699=>"011100000",
116700=>"111111001",
116701=>"111011000",
116702=>"111100000",
116703=>"101000000",
116704=>"000000000",
116705=>"111000011",
116706=>"111001011",
116707=>"000111111",
116708=>"000101100",
116709=>"100100111",
116710=>"000000000",
116711=>"100111111",
116712=>"011000111",
116713=>"000001101",
116714=>"100111011",
116715=>"000000000",
116716=>"000100100",
116717=>"011001101",
116718=>"001000000",
116719=>"010000111",
116720=>"000111100",
116721=>"000100000",
116722=>"111000000",
116723=>"111010000",
116724=>"011000001",
116725=>"111111110",
116726=>"000010101",
116727=>"111110011",
116728=>"000000000",
116729=>"111101101",
116730=>"000101100",
116731=>"111010010",
116732=>"000011111",
116733=>"100100010",
116734=>"101001111",
116735=>"000000001",
116736=>"011001011",
116737=>"000101101",
116738=>"001001000",
116739=>"000001000",
116740=>"001000101",
116741=>"111110000",
116742=>"010111111",
116743=>"001110110",
116744=>"110111110",
116745=>"111111111",
116746=>"001000000",
116747=>"010000000",
116748=>"000010111",
116749=>"110111101",
116750=>"010101001",
116751=>"000001100",
116752=>"000000001",
116753=>"111111110",
116754=>"100111001",
116755=>"010100000",
116756=>"110010101",
116757=>"111101111",
116758=>"000001001",
116759=>"000001001",
116760=>"100111111",
116761=>"001000101",
116762=>"010000000",
116763=>"000111111",
116764=>"111000000",
116765=>"000101010",
116766=>"010100010",
116767=>"000111111",
116768=>"111000000",
116769=>"110000111",
116770=>"001001110",
116771=>"000110000",
116772=>"000010011",
116773=>"111000100",
116774=>"000000000",
116775=>"011100110",
116776=>"011001000",
116777=>"110110000",
116778=>"110000000",
116779=>"000000000",
116780=>"111001001",
116781=>"001001100",
116782=>"111000111",
116783=>"100111100",
116784=>"000000001",
116785=>"011111100",
116786=>"000000111",
116787=>"000000000",
116788=>"000010110",
116789=>"100011010",
116790=>"000000000",
116791=>"000101101",
116792=>"000010011",
116793=>"001101111",
116794=>"001101101",
116795=>"010110100",
116796=>"110111011",
116797=>"111111111",
116798=>"000000100",
116799=>"011111010",
116800=>"000010111",
116801=>"000101111",
116802=>"101101101",
116803=>"011001001",
116804=>"111101000",
116805=>"110110110",
116806=>"000000011",
116807=>"111010000",
116808=>"000111101",
116809=>"111000101",
116810=>"001000111",
116811=>"111110010",
116812=>"111111100",
116813=>"110110111",
116814=>"110110011",
116815=>"011111111",
116816=>"000000010",
116817=>"000111111",
116818=>"010111001",
116819=>"011011111",
116820=>"101101001",
116821=>"110111110",
116822=>"011111001",
116823=>"001000000",
116824=>"111111001",
116825=>"100000100",
116826=>"100111100",
116827=>"111010011",
116828=>"000101101",
116829=>"010010000",
116830=>"101111011",
116831=>"100001111",
116832=>"110111101",
116833=>"000001001",
116834=>"001000000",
116835=>"011011001",
116836=>"001010111",
116837=>"100000111",
116838=>"000000000",
116839=>"110111100",
116840=>"111001000",
116841=>"111000000",
116842=>"101001101",
116843=>"100000110",
116844=>"110111111",
116845=>"000000000",
116846=>"110010000",
116847=>"111010000",
116848=>"110000101",
116849=>"000000000",
116850=>"001001000",
116851=>"101010000",
116852=>"110011000",
116853=>"111000001",
116854=>"011111111",
116855=>"111110110",
116856=>"000001000",
116857=>"101000111",
116858=>"000100000",
116859=>"001101001",
116860=>"110000001",
116861=>"100100100",
116862=>"001000111",
116863=>"110000000",
116864=>"101111110",
116865=>"000000000",
116866=>"111111111",
116867=>"000101111",
116868=>"110111111",
116869=>"000100111",
116870=>"111001011",
116871=>"000000100",
116872=>"100000000",
116873=>"001101111",
116874=>"101001110",
116875=>"010000000",
116876=>"110000000",
116877=>"010001000",
116878=>"000010010",
116879=>"001000001",
116880=>"101000100",
116881=>"000000111",
116882=>"010100010",
116883=>"000000110",
116884=>"000010010",
116885=>"111000000",
116886=>"010000101",
116887=>"010011011",
116888=>"111010000",
116889=>"101001110",
116890=>"001101001",
116891=>"000000011",
116892=>"000100000",
116893=>"000000110",
116894=>"100101101",
116895=>"010000000",
116896=>"001100101",
116897=>"001000000",
116898=>"011101111",
116899=>"000000000",
116900=>"111000000",
116901=>"001111111",
116902=>"110110000",
116903=>"110000001",
116904=>"010000001",
116905=>"000101010",
116906=>"110111000",
116907=>"011000000",
116908=>"111111110",
116909=>"001001000",
116910=>"100000100",
116911=>"001001111",
116912=>"111001110",
116913=>"100011011",
116914=>"111111000",
116915=>"001010000",
116916=>"001100111",
116917=>"110010000",
116918=>"000100111",
116919=>"110110000",
116920=>"011011110",
116921=>"000000110",
116922=>"111000000",
116923=>"001111111",
116924=>"100110111",
116925=>"111110000",
116926=>"110110011",
116927=>"000000000",
116928=>"001001111",
116929=>"000111000",
116930=>"100101111",
116931=>"000010001",
116932=>"101101000",
116933=>"001001001",
116934=>"001010010",
116935=>"110101001",
116936=>"111101011",
116937=>"000111111",
116938=>"001100110",
116939=>"111110110",
116940=>"011100110",
116941=>"011000000",
116942=>"000000000",
116943=>"110110111",
116944=>"000000000",
116945=>"110100001",
116946=>"011010000",
116947=>"001111100",
116948=>"000010000",
116949=>"001100100",
116950=>"110000000",
116951=>"101111111",
116952=>"100111101",
116953=>"000000000",
116954=>"000100111",
116955=>"101000000",
116956=>"100010001",
116957=>"010111110",
116958=>"110111010",
116959=>"001001000",
116960=>"101110010",
116961=>"101001111",
116962=>"000000000",
116963=>"001110110",
116964=>"111001000",
116965=>"110010000",
116966=>"110010101",
116967=>"111111111",
116968=>"000000000",
116969=>"000000000",
116970=>"111100000",
116971=>"000000000",
116972=>"000000000",
116973=>"010001010",
116974=>"001000001",
116975=>"011110000",
116976=>"111110000",
116977=>"000000000",
116978=>"101000011",
116979=>"100111011",
116980=>"110100110",
116981=>"100100000",
116982=>"000001000",
116983=>"001001010",
116984=>"000000000",
116985=>"101101001",
116986=>"111111111",
116987=>"000111111",
116988=>"001101111",
116989=>"011000000",
116990=>"010100100",
116991=>"000001111",
116992=>"011010100",
116993=>"110110110",
116994=>"111000000",
116995=>"110110001",
116996=>"000111111",
116997=>"100000100",
116998=>"111111000",
116999=>"110100110",
117000=>"111001111",
117001=>"110000000",
117002=>"000000100",
117003=>"100111111",
117004=>"100000000",
117005=>"000111111",
117006=>"000000000",
117007=>"110100000",
117008=>"110110110",
117009=>"111111110",
117010=>"111011011",
117011=>"000110101",
117012=>"111110111",
117013=>"110111000",
117014=>"010001001",
117015=>"110010110",
117016=>"001110101",
117017=>"110100111",
117018=>"010111000",
117019=>"111011010",
117020=>"101110111",
117021=>"010010111",
117022=>"111000010",
117023=>"100101001",
117024=>"100000100",
117025=>"010110111",
117026=>"101001000",
117027=>"101111010",
117028=>"001000001",
117029=>"000010010",
117030=>"111001001",
117031=>"110110110",
117032=>"100000000",
117033=>"001111110",
117034=>"110100000",
117035=>"101111111",
117036=>"000011001",
117037=>"111001000",
117038=>"101111000",
117039=>"111110110",
117040=>"110000001",
117041=>"000011111",
117042=>"011110010",
117043=>"011010001",
117044=>"111010000",
117045=>"000000110",
117046=>"000100110",
117047=>"000000110",
117048=>"110000110",
117049=>"010110100",
117050=>"101000000",
117051=>"000000000",
117052=>"100000011",
117053=>"000101001",
117054=>"000000000",
117055=>"111001001",
117056=>"111010110",
117057=>"111111110",
117058=>"111111001",
117059=>"011011000",
117060=>"000110000",
117061=>"110000011",
117062=>"000001111",
117063=>"111011000",
117064=>"100100100",
117065=>"111001110",
117066=>"000000001",
117067=>"001000000",
117068=>"111000000",
117069=>"000000000",
117070=>"001111101",
117071=>"000000110",
117072=>"000001101",
117073=>"110010000",
117074=>"110101010",
117075=>"011001101",
117076=>"111100000",
117077=>"111000000",
117078=>"011011111",
117079=>"110111000",
117080=>"000010010",
117081=>"000001001",
117082=>"000110111",
117083=>"011000001",
117084=>"011111111",
117085=>"011011001",
117086=>"111110010",
117087=>"100100000",
117088=>"100110111",
117089=>"111110000",
117090=>"111000000",
117091=>"000011011",
117092=>"000001101",
117093=>"111111111",
117094=>"100100110",
117095=>"110001001",
117096=>"100000001",
117097=>"110000000",
117098=>"101000000",
117099=>"000011110",
117100=>"000000010",
117101=>"000110110",
117102=>"000111001",
117103=>"110000100",
117104=>"101100101",
117105=>"000111000",
117106=>"000001111",
117107=>"111010011",
117108=>"110110000",
117109=>"001000001",
117110=>"001101000",
117111=>"111000000",
117112=>"111110100",
117113=>"111110110",
117114=>"011110101",
117115=>"111000000",
117116=>"100000011",
117117=>"100000000",
117118=>"110110011",
117119=>"001001000",
117120=>"000110110",
117121=>"111000000",
117122=>"111000010",
117123=>"010010000",
117124=>"000000111",
117125=>"111001011",
117126=>"000111001",
117127=>"000110110",
117128=>"001100001",
117129=>"000010110",
117130=>"000000001",
117131=>"010000010",
117132=>"101110000",
117133=>"110000000",
117134=>"011111000",
117135=>"000000000",
117136=>"111001001",
117137=>"001011000",
117138=>"001010000",
117139=>"000000111",
117140=>"001000110",
117141=>"110111110",
117142=>"000000010",
117143=>"100001010",
117144=>"110100000",
117145=>"110000000",
117146=>"111000000",
117147=>"110111000",
117148=>"000001001",
117149=>"111000000",
117150=>"011101000",
117151=>"010111010",
117152=>"000110001",
117153=>"111111110",
117154=>"101101000",
117155=>"110011001",
117156=>"111110110",
117157=>"000100111",
117158=>"111111001",
117159=>"111111000",
117160=>"000010000",
117161=>"010000001",
117162=>"111111001",
117163=>"000110010",
117164=>"001000111",
117165=>"101001000",
117166=>"100110111",
117167=>"010001111",
117168=>"101110110",
117169=>"000100111",
117170=>"110000000",
117171=>"001001000",
117172=>"101001000",
117173=>"000000001",
117174=>"010000111",
117175=>"000000000",
117176=>"001010000",
117177=>"000001100",
117178=>"101111000",
117179=>"010010011",
117180=>"111111001",
117181=>"110111101",
117182=>"111000000",
117183=>"010010110",
117184=>"001001111",
117185=>"000001111",
117186=>"110111111",
117187=>"111001000",
117188=>"000000010",
117189=>"000001101",
117190=>"010000000",
117191=>"101001000",
117192=>"110000000",
117193=>"001100111",
117194=>"000111111",
117195=>"000110110",
117196=>"111111000",
117197=>"011100100",
117198=>"000010111",
117199=>"110010111",
117200=>"000000000",
117201=>"000101111",
117202=>"000111101",
117203=>"001111011",
117204=>"101001000",
117205=>"000111111",
117206=>"011111000",
117207=>"110110110",
117208=>"000100110",
117209=>"000110111",
117210=>"011010000",
117211=>"000000011",
117212=>"010000001",
117213=>"111000000",
117214=>"010010111",
117215=>"010110110",
117216=>"111011111",
117217=>"110001111",
117218=>"111000000",
117219=>"001100010",
117220=>"111010000",
117221=>"001001100",
117222=>"100110100",
117223=>"011111111",
117224=>"111110000",
117225=>"000010100",
117226=>"001001100",
117227=>"111111000",
117228=>"000100000",
117229=>"000110111",
117230=>"010010010",
117231=>"001101100",
117232=>"111000110",
117233=>"000111011",
117234=>"111011001",
117235=>"000001011",
117236=>"100110010",
117237=>"000000111",
117238=>"000000000",
117239=>"111111110",
117240=>"000110110",
117241=>"110001011",
117242=>"111000111",
117243=>"001001111",
117244=>"111001000",
117245=>"000010000",
117246=>"000000000",
117247=>"101001001",
117248=>"010011001",
117249=>"110111111",
117250=>"111000101",
117251=>"000010000",
117252=>"001100110",
117253=>"111010000",
117254=>"101111111",
117255=>"000100000",
117256=>"000100110",
117257=>"000101100",
117258=>"000000011",
117259=>"110111000",
117260=>"000000100",
117261=>"011000100",
117262=>"001011010",
117263=>"111011001",
117264=>"111111000",
117265=>"100101101",
117266=>"010111100",
117267=>"111111000",
117268=>"101110110",
117269=>"000001011",
117270=>"111011011",
117271=>"011111000",
117272=>"010011000",
117273=>"010010000",
117274=>"000111011",
117275=>"000111111",
117276=>"111000010",
117277=>"000111111",
117278=>"111000000",
117279=>"000010010",
117280=>"010010110",
117281=>"000010000",
117282=>"000000001",
117283=>"000011111",
117284=>"000010010",
117285=>"011111010",
117286=>"000100000",
117287=>"111011111",
117288=>"001011111",
117289=>"000000000",
117290=>"110111110",
117291=>"111100100",
117292=>"100111100",
117293=>"101010000",
117294=>"011010000",
117295=>"111111100",
117296=>"111101100",
117297=>"101011001",
117298=>"101110001",
117299=>"111111000",
117300=>"111000111",
117301=>"000101010",
117302=>"001110100",
117303=>"010111010",
117304=>"111101001",
117305=>"000000000",
117306=>"010011010",
117307=>"101111101",
117308=>"110110100",
117309=>"101011011",
117310=>"111111101",
117311=>"010111111",
117312=>"111101000",
117313=>"111011000",
117314=>"111000000",
117315=>"111111011",
117316=>"110111010",
117317=>"000111011",
117318=>"111000010",
117319=>"111111010",
117320=>"000110100",
117321=>"000111000",
117322=>"000111000",
117323=>"000010000",
117324=>"111000000",
117325=>"000011000",
117326=>"000100010",
117327=>"111000111",
117328=>"010111111",
117329=>"000111111",
117330=>"011111010",
117331=>"111011001",
117332=>"101111010",
117333=>"111011011",
117334=>"100111011",
117335=>"111101111",
117336=>"110110100",
117337=>"011011011",
117338=>"000011011",
117339=>"110111000",
117340=>"111110000",
117341=>"100111011",
117342=>"110000100",
117343=>"111101110",
117344=>"100111111",
117345=>"010010011",
117346=>"111101111",
117347=>"110100110",
117348=>"000010000",
117349=>"001010011",
117350=>"000000000",
117351=>"000111000",
117352=>"110111010",
117353=>"111111101",
117354=>"000011110",
117355=>"110101000",
117356=>"000000100",
117357=>"000111000",
117358=>"110111000",
117359=>"011111111",
117360=>"100110111",
117361=>"000000111",
117362=>"110011001",
117363=>"100001101",
117364=>"110010010",
117365=>"011110000",
117366=>"101101100",
117367=>"110111101",
117368=>"111111110",
117369=>"000111110",
117370=>"001000010",
117371=>"000000000",
117372=>"100110110",
117373=>"011110100",
117374=>"101100111",
117375=>"010000111",
117376=>"111110000",
117377=>"111100000",
117378=>"010111111",
117379=>"000011011",
117380=>"100000000",
117381=>"110110100",
117382=>"111111000",
117383=>"010111011",
117384=>"001011011",
117385=>"000001010",
117386=>"000011000",
117387=>"111111000",
117388=>"101010011",
117389=>"111101010",
117390=>"110101111",
117391=>"101001010",
117392=>"100010011",
117393=>"111111010",
117394=>"010010000",
117395=>"111111110",
117396=>"011111111",
117397=>"111101101",
117398=>"101001001",
117399=>"000110010",
117400=>"000001000",
117401=>"111111001",
117402=>"011111000",
117403=>"111000111",
117404=>"000010000",
117405=>"111001110",
117406=>"111111101",
117407=>"000000000",
117408=>"000011000",
117409=>"101111111",
117410=>"010111101",
117411=>"000100010",
117412=>"100101100",
117413=>"100110100",
117414=>"001111000",
117415=>"011100000",
117416=>"101100101",
117417=>"000110111",
117418=>"100100100",
117419=>"111000111",
117420=>"111111001",
117421=>"111011101",
117422=>"011110111",
117423=>"000000000",
117424=>"011011111",
117425=>"011011000",
117426=>"110011000",
117427=>"101110110",
117428=>"000011000",
117429=>"101111000",
117430=>"000011011",
117431=>"010010001",
117432=>"011011001",
117433=>"000011010",
117434=>"010111111",
117435=>"100110010",
117436=>"111010101",
117437=>"111001101",
117438=>"000011011",
117439=>"010001001",
117440=>"010000010",
117441=>"111111111",
117442=>"111111000",
117443=>"101111111",
117444=>"000000001",
117445=>"111111110",
117446=>"011111110",
117447=>"111111111",
117448=>"000111010",
117449=>"101111010",
117450=>"111111011",
117451=>"101101111",
117452=>"111011011",
117453=>"011011110",
117454=>"111010111",
117455=>"010111010",
117456=>"101000001",
117457=>"000010000",
117458=>"000010010",
117459=>"000011111",
117460=>"111000111",
117461=>"110110110",
117462=>"101000000",
117463=>"010111101",
117464=>"000000000",
117465=>"000111010",
117466=>"000110000",
117467=>"111000111",
117468=>"111110110",
117469=>"000000000",
117470=>"000010000",
117471=>"000011100",
117472=>"111000010",
117473=>"101100111",
117474=>"000000101",
117475=>"000001111",
117476=>"101101000",
117477=>"110110010",
117478=>"111111111",
117479=>"100110110",
117480=>"110011000",
117481=>"110111101",
117482=>"011001100",
117483=>"000000111",
117484=>"000100110",
117485=>"010111010",
117486=>"111111111",
117487=>"000110001",
117488=>"111111000",
117489=>"010110110",
117490=>"011000001",
117491=>"000110100",
117492=>"000011011",
117493=>"010000011",
117494=>"111010010",
117495=>"111111010",
117496=>"011100000",
117497=>"011010000",
117498=>"000000000",
117499=>"000111111",
117500=>"011011000",
117501=>"110110100",
117502=>"000011001",
117503=>"101000101",
117504=>"100110011",
117505=>"111011000",
117506=>"001000001",
117507=>"010011000",
117508=>"111110110",
117509=>"101101000",
117510=>"000100101",
117511=>"000011011",
117512=>"111110110",
117513=>"000111010",
117514=>"100100110",
117515=>"000000000",
117516=>"111111111",
117517=>"000000000",
117518=>"011010000",
117519=>"000000100",
117520=>"000100111",
117521=>"110100000",
117522=>"001000000",
117523=>"111110111",
117524=>"000000000",
117525=>"000100000",
117526=>"000011111",
117527=>"111111010",
117528=>"111111010",
117529=>"011000001",
117530=>"001000000",
117531=>"010100110",
117532=>"100000100",
117533=>"101000101",
117534=>"001000111",
117535=>"011111011",
117536=>"100111000",
117537=>"000010110",
117538=>"100000000",
117539=>"011000000",
117540=>"011010100",
117541=>"100101100",
117542=>"000010010",
117543=>"111000111",
117544=>"000010001",
117545=>"000000010",
117546=>"111000111",
117547=>"000111111",
117548=>"010010011",
117549=>"010010000",
117550=>"100111111",
117551=>"000000000",
117552=>"100010010",
117553=>"101111111",
117554=>"110000011",
117555=>"000010011",
117556=>"110100101",
117557=>"010100000",
117558=>"000111110",
117559=>"000110000",
117560=>"010011010",
117561=>"111101000",
117562=>"000110000",
117563=>"000100010",
117564=>"000001110",
117565=>"111111101",
117566=>"000000110",
117567=>"001101011",
117568=>"111011000",
117569=>"000000000",
117570=>"010111000",
117571=>"110111110",
117572=>"000000000",
117573=>"011001000",
117574=>"111000010",
117575=>"011100000",
117576=>"001010111",
117577=>"111001111",
117578=>"011000010",
117579=>"101000000",
117580=>"111100111",
117581=>"111111111",
117582=>"111111111",
117583=>"110111111",
117584=>"001001011",
117585=>"111111111",
117586=>"000000110",
117587=>"000011001",
117588=>"000001100",
117589=>"000011100",
117590=>"100110110",
117591=>"011000111",
117592=>"111001111",
117593=>"111111001",
117594=>"001001001",
117595=>"001000000",
117596=>"000000000",
117597=>"101111001",
117598=>"000000000",
117599=>"011111100",
117600=>"111111101",
117601=>"100000000",
117602=>"011101111",
117603=>"000000000",
117604=>"010011011",
117605=>"000001000",
117606=>"000000000",
117607=>"111111110",
117608=>"100010000",
117609=>"000100000",
117610=>"000010110",
117611=>"100000100",
117612=>"111100000",
117613=>"000100100",
117614=>"000000111",
117615=>"100100111",
117616=>"100000000",
117617=>"100100010",
117618=>"000110010",
117619=>"011110100",
117620=>"100000011",
117621=>"111000000",
117622=>"111010000",
117623=>"010000000",
117624=>"111111000",
117625=>"010111010",
117626=>"000100010",
117627=>"110011011",
117628=>"110001001",
117629=>"000011010",
117630=>"100100001",
117631=>"011101101",
117632=>"000111000",
117633=>"100111110",
117634=>"000010000",
117635=>"111111111",
117636=>"000000000",
117637=>"000010000",
117638=>"101110011",
117639=>"001000010",
117640=>"011110000",
117641=>"010101100",
117642=>"011000010",
117643=>"000111011",
117644=>"000000000",
117645=>"111100000",
117646=>"110110000",
117647=>"100000000",
117648=>"110110111",
117649=>"000010000",
117650=>"000000010",
117651=>"100000110",
117652=>"111000000",
117653=>"100111111",
117654=>"111110100",
117655=>"011111011",
117656=>"000100000",
117657=>"011111010",
117658=>"101101111",
117659=>"111110000",
117660=>"000000011",
117661=>"010111111",
117662=>"100011010",
117663=>"110111110",
117664=>"011011011",
117665=>"000110000",
117666=>"111110111",
117667=>"100111111",
117668=>"000110010",
117669=>"100110110",
117670=>"011000011",
117671=>"111100110",
117672=>"110110100",
117673=>"111111101",
117674=>"010011010",
117675=>"111111100",
117676=>"101101100",
117677=>"011101111",
117678=>"100011010",
117679=>"001111111",
117680=>"100000001",
117681=>"100111111",
117682=>"000011011",
117683=>"110111111",
117684=>"111011101",
117685=>"111010000",
117686=>"001000000",
117687=>"001100000",
117688=>"100110100",
117689=>"101010100",
117690=>"110000000",
117691=>"111000000",
117692=>"011000000",
117693=>"010101111",
117694=>"110110010",
117695=>"000000000",
117696=>"000111111",
117697=>"010111010",
117698=>"100110100",
117699=>"000000101",
117700=>"000000100",
117701=>"000110111",
117702=>"001111000",
117703=>"000000000",
117704=>"111101000",
117705=>"001000000",
117706=>"111100001",
117707=>"000100010",
117708=>"010010010",
117709=>"001100100",
117710=>"100111000",
117711=>"101111111",
117712=>"000010000",
117713=>"110111010",
117714=>"111011001",
117715=>"111111011",
117716=>"011011011",
117717=>"110111000",
117718=>"010010010",
117719=>"111111110",
117720=>"010111111",
117721=>"000000000",
117722=>"000110111",
117723=>"000000000",
117724=>"010110000",
117725=>"111001011",
117726=>"000000000",
117727=>"111001111",
117728=>"000000101",
117729=>"000011000",
117730=>"000101111",
117731=>"111011111",
117732=>"011010010",
117733=>"000000000",
117734=>"111000100",
117735=>"110111110",
117736=>"111100011",
117737=>"001001011",
117738=>"101000000",
117739=>"111110111",
117740=>"000100101",
117741=>"111101111",
117742=>"001101000",
117743=>"000010000",
117744=>"111111001",
117745=>"110011011",
117746=>"100111010",
117747=>"100110000",
117748=>"000011111",
117749=>"000000001",
117750=>"101011000",
117751=>"111010100",
117752=>"000000000",
117753=>"000000110",
117754=>"111111111",
117755=>"000100100",
117756=>"100111111",
117757=>"000001000",
117758=>"111111011",
117759=>"111000000",
117760=>"111110111",
117761=>"000000001",
117762=>"111101000",
117763=>"111111001",
117764=>"111010000",
117765=>"011011000",
117766=>"000101100",
117767=>"000111000",
117768=>"111111000",
117769=>"000000101",
117770=>"110100000",
117771=>"110111110",
117772=>"111111101",
117773=>"111111110",
117774=>"111111000",
117775=>"000011111",
117776=>"111011000",
117777=>"111101001",
117778=>"111111101",
117779=>"100101001",
117780=>"111111000",
117781=>"111111000",
117782=>"000000111",
117783=>"100001111",
117784=>"111111001",
117785=>"110000010",
117786=>"111111101",
117787=>"000000101",
117788=>"000000000",
117789=>"010111101",
117790=>"111010110",
117791=>"111000001",
117792=>"011111111",
117793=>"110010000",
117794=>"000100110",
117795=>"000000000",
117796=>"000010010",
117797=>"001001111",
117798=>"111111000",
117799=>"000000110",
117800=>"111111001",
117801=>"000111110",
117802=>"000000111",
117803=>"000000000",
117804=>"000000110",
117805=>"100101001",
117806=>"000010100",
117807=>"111001000",
117808=>"000010111",
117809=>"000010111",
117810=>"010111000",
117811=>"000010111",
117812=>"100001111",
117813=>"011101111",
117814=>"011111111",
117815=>"101010111",
117816=>"101000101",
117817=>"111100000",
117818=>"000111111",
117819=>"110101000",
117820=>"000010011",
117821=>"000111111",
117822=>"011000000",
117823=>"000000011",
117824=>"111100000",
117825=>"000010010",
117826=>"101111000",
117827=>"100101100",
117828=>"010111111",
117829=>"000011001",
117830=>"010000111",
117831=>"000000001",
117832=>"010101010",
117833=>"010011000",
117834=>"111111101",
117835=>"101111111",
117836=>"000010000",
117837=>"011000001",
117838=>"010011011",
117839=>"000111111",
117840=>"111101101",
117841=>"011011111",
117842=>"000001111",
117843=>"000110111",
117844=>"011111000",
117845=>"000010110",
117846=>"100010001",
117847=>"111111110",
117848=>"100100000",
117849=>"000000001",
117850=>"001000000",
117851=>"100000010",
117852=>"101101000",
117853=>"011110000",
117854=>"111111010",
117855=>"001001011",
117856=>"001000011",
117857=>"000111101",
117858=>"111111000",
117859=>"110110011",
117860=>"100111000",
117861=>"000101111",
117862=>"000100100",
117863=>"000000000",
117864=>"110010101",
117865=>"111111111",
117866=>"000000111",
117867=>"000000011",
117868=>"000111001",
117869=>"101000000",
117870=>"111111000",
117871=>"000000111",
117872=>"000001000",
117873=>"000000000",
117874=>"110111110",
117875=>"011111101",
117876=>"000000000",
117877=>"111101000",
117878=>"000001111",
117879=>"000001000",
117880=>"001101111",
117881=>"000000110",
117882=>"000001000",
117883=>"111110001",
117884=>"010011001",
117885=>"000011111",
117886=>"111111110",
117887=>"001000000",
117888=>"000010010",
117889=>"100011111",
117890=>"000000111",
117891=>"000111100",
117892=>"101101100",
117893=>"111101111",
117894=>"000000111",
117895=>"010110000",
117896=>"000010000",
117897=>"001101000",
117898=>"111111000",
117899=>"010111111",
117900=>"111111000",
117901=>"111001111",
117902=>"000000001",
117903=>"111111000",
117904=>"110110100",
117905=>"111101101",
117906=>"000000111",
117907=>"000110110",
117908=>"111010000",
117909=>"111000000",
117910=>"111000110",
117911=>"010110100",
117912=>"000000011",
117913=>"000000111",
117914=>"111111010",
117915=>"111111000",
117916=>"000001000",
117917=>"000110001",
117918=>"000000111",
117919=>"000111001",
117920=>"010100010",
117921=>"111000010",
117922=>"011000110",
117923=>"000000000",
117924=>"110000000",
117925=>"001011000",
117926=>"000000010",
117927=>"000001000",
117928=>"111000000",
117929=>"111101101",
117930=>"111111000",
117931=>"101111000",
117932=>"001000000",
117933=>"010111000",
117934=>"111010111",
117935=>"011010001",
117936=>"000000001",
117937=>"111001001",
117938=>"100100001",
117939=>"000000000",
117940=>"001110111",
117941=>"011101111",
117942=>"111101100",
117943=>"000001011",
117944=>"000000000",
117945=>"000000000",
117946=>"000000101",
117947=>"000010111",
117948=>"111111100",
117949=>"111010000",
117950=>"011011000",
117951=>"010111101",
117952=>"111111000",
117953=>"001000111",
117954=>"101111011",
117955=>"000110011",
117956=>"000000010",
117957=>"110001000",
117958=>"000000000",
117959=>"110110010",
117960=>"000100011",
117961=>"111100100",
117962=>"110001000",
117963=>"111000000",
117964=>"010000000",
117965=>"000110100",
117966=>"000000100",
117967=>"111110000",
117968=>"001010111",
117969=>"011011001",
117970=>"111111000",
117971=>"000011111",
117972=>"111001000",
117973=>"101110110",
117974=>"111111000",
117975=>"001110111",
117976=>"000111111",
117977=>"111111000",
117978=>"000001000",
117979=>"011111101",
117980=>"000111111",
117981=>"001100110",
117982=>"001100001",
117983=>"111110111",
117984=>"111111000",
117985=>"111101001",
117986=>"010010111",
117987=>"111111000",
117988=>"111011001",
117989=>"111000000",
117990=>"001111011",
117991=>"000010110",
117992=>"010010111",
117993=>"000000101",
117994=>"011001001",
117995=>"101001001",
117996=>"101101010",
117997=>"000000010",
117998=>"010111000",
117999=>"000110000",
118000=>"000000111",
118001=>"110010000",
118002=>"000000000",
118003=>"000111111",
118004=>"001011110",
118005=>"111110000",
118006=>"000000100",
118007=>"010111000",
118008=>"111011111",
118009=>"110000111",
118010=>"000010000",
118011=>"111110001",
118012=>"100000111",
118013=>"000000101",
118014=>"010000111",
118015=>"000000000",
118016=>"000111110",
118017=>"000100000",
118018=>"001100100",
118019=>"000110000",
118020=>"000011110",
118021=>"001010110",
118022=>"110100010",
118023=>"000000011",
118024=>"110100100",
118025=>"000000010",
118026=>"111111010",
118027=>"000011000",
118028=>"100100011",
118029=>"010111010",
118030=>"000101001",
118031=>"100000100",
118032=>"111100001",
118033=>"111110100",
118034=>"101100101",
118035=>"100000000",
118036=>"101001100",
118037=>"000011111",
118038=>"111110000",
118039=>"000011010",
118040=>"011111100",
118041=>"011010011",
118042=>"001100100",
118043=>"000100000",
118044=>"101011111",
118045=>"111011010",
118046=>"011111111",
118047=>"000000010",
118048=>"000100000",
118049=>"000000000",
118050=>"111001111",
118051=>"111111011",
118052=>"000001000",
118053=>"010000101",
118054=>"101000100",
118055=>"000111101",
118056=>"111101111",
118057=>"001000101",
118058=>"000000100",
118059=>"111100100",
118060=>"100110001",
118061=>"111111101",
118062=>"100101111",
118063=>"010111000",
118064=>"000010000",
118065=>"011011010",
118066=>"011101011",
118067=>"000111111",
118068=>"000101111",
118069=>"100010101",
118070=>"010100000",
118071=>"010011011",
118072=>"111100111",
118073=>"101111101",
118074=>"111100000",
118075=>"010011011",
118076=>"001011001",
118077=>"111111111",
118078=>"000000000",
118079=>"110111011",
118080=>"010100100",
118081=>"111011100",
118082=>"101000000",
118083=>"111000101",
118084=>"111000010",
118085=>"000000100",
118086=>"000011010",
118087=>"110001001",
118088=>"100100110",
118089=>"010011010",
118090=>"001000100",
118091=>"000011011",
118092=>"101100111",
118093=>"110000110",
118094=>"100110111",
118095=>"110010111",
118096=>"011000000",
118097=>"011010000",
118098=>"000010111",
118099=>"001001000",
118100=>"111101000",
118101=>"010000000",
118102=>"100110010",
118103=>"011111111",
118104=>"000001100",
118105=>"000100110",
118106=>"000110110",
118107=>"001011000",
118108=>"100100100",
118109=>"001001001",
118110=>"111111100",
118111=>"000111011",
118112=>"111100100",
118113=>"001000100",
118114=>"111000001",
118115=>"010111011",
118116=>"000000000",
118117=>"000100110",
118118=>"000000000",
118119=>"000000010",
118120=>"100111010",
118121=>"001001111",
118122=>"111000100",
118123=>"110001111",
118124=>"111000000",
118125=>"011111111",
118126=>"000011010",
118127=>"000000010",
118128=>"001011011",
118129=>"011000000",
118130=>"100001110",
118131=>"100100000",
118132=>"011111000",
118133=>"100101111",
118134=>"100010111",
118135=>"111000110",
118136=>"011100110",
118137=>"100000110",
118138=>"010010000",
118139=>"101111000",
118140=>"110111011",
118141=>"100111110",
118142=>"110000000",
118143=>"100011011",
118144=>"011010000",
118145=>"000000001",
118146=>"010011000",
118147=>"000011010",
118148=>"011011001",
118149=>"000011011",
118150=>"101101000",
118151=>"001101111",
118152=>"000110000",
118153=>"110111010",
118154=>"000111000",
118155=>"100111111",
118156=>"000101100",
118157=>"101000100",
118158=>"100111111",
118159=>"110101001",
118160=>"101110110",
118161=>"011000000",
118162=>"000011011",
118163=>"110010101",
118164=>"000000000",
118165=>"001101101",
118166=>"111100100",
118167=>"111100110",
118168=>"010000000",
118169=>"101101011",
118170=>"111000000",
118171=>"111011111",
118172=>"000011011",
118173=>"100111111",
118174=>"011111110",
118175=>"111101010",
118176=>"101011110",
118177=>"111110100",
118178=>"000101111",
118179=>"110111110",
118180=>"000010100",
118181=>"100110110",
118182=>"110001101",
118183=>"110100000",
118184=>"000000000",
118185=>"111111100",
118186=>"111100000",
118187=>"000101100",
118188=>"000001000",
118189=>"000001011",
118190=>"110011000",
118191=>"111001100",
118192=>"111100100",
118193=>"001011001",
118194=>"101100101",
118195=>"100100111",
118196=>"100011001",
118197=>"000000100",
118198=>"111100100",
118199=>"001100001",
118200=>"111010010",
118201=>"000011011",
118202=>"101011000",
118203=>"000111100",
118204=>"111011011",
118205=>"111111111",
118206=>"000000011",
118207=>"001000101",
118208=>"111101111",
118209=>"000000111",
118210=>"011011000",
118211=>"000000100",
118212=>"000011100",
118213=>"110110110",
118214=>"000011011",
118215=>"111101111",
118216=>"111111000",
118217=>"000000000",
118218=>"000110100",
118219=>"000011011",
118220=>"101101110",
118221=>"001111110",
118222=>"000100101",
118223=>"010001001",
118224=>"111111100",
118225=>"111011011",
118226=>"011010010",
118227=>"111111000",
118228=>"010100010",
118229=>"000100100",
118230=>"000000000",
118231=>"010011000",
118232=>"010111011",
118233=>"010111100",
118234=>"110110111",
118235=>"010100100",
118236=>"100001000",
118237=>"110100000",
118238=>"111101111",
118239=>"100000000",
118240=>"100100000",
118241=>"111111001",
118242=>"001011101",
118243=>"001011000",
118244=>"111010000",
118245=>"000010100",
118246=>"101010010",
118247=>"010111100",
118248=>"111000101",
118249=>"010101001",
118250=>"101000011",
118251=>"111101101",
118252=>"000000111",
118253=>"000000000",
118254=>"111100010",
118255=>"011100100",
118256=>"100100111",
118257=>"100011001",
118258=>"101011111",
118259=>"110101100",
118260=>"000001011",
118261=>"000101000",
118262=>"100000101",
118263=>"111111000",
118264=>"000001000",
118265=>"111000010",
118266=>"010000000",
118267=>"011011101",
118268=>"000000000",
118269=>"000011011",
118270=>"001001000",
118271=>"000011011",
118272=>"011000000",
118273=>"000010000",
118274=>"101101111",
118275=>"000100111",
118276=>"100011010",
118277=>"011000010",
118278=>"011111010",
118279=>"000011110",
118280=>"000000000",
118281=>"000000101",
118282=>"001011001",
118283=>"100111000",
118284=>"001000110",
118285=>"101111101",
118286=>"011111100",
118287=>"110001111",
118288=>"010101111",
118289=>"101111000",
118290=>"101111111",
118291=>"000010100",
118292=>"000000010",
118293=>"010010000",
118294=>"000000111",
118295=>"000111100",
118296=>"111100111",
118297=>"001001000",
118298=>"100100110",
118299=>"111000100",
118300=>"000000000",
118301=>"101000101",
118302=>"010000101",
118303=>"100111000",
118304=>"010010111",
118305=>"110110111",
118306=>"111010000",
118307=>"000000000",
118308=>"000111001",
118309=>"011000000",
118310=>"010111000",
118311=>"001010000",
118312=>"000000111",
118313=>"011110101",
118314=>"010010100",
118315=>"111101111",
118316=>"001000001",
118317=>"101000111",
118318=>"011000101",
118319=>"100000111",
118320=>"010101000",
118321=>"110001000",
118322=>"000000101",
118323=>"000000000",
118324=>"111110101",
118325=>"010001000",
118326=>"011011010",
118327=>"000000001",
118328=>"111000010",
118329=>"000000101",
118330=>"000001010",
118331=>"111000101",
118332=>"000001000",
118333=>"111010110",
118334=>"000000111",
118335=>"110000100",
118336=>"100000001",
118337=>"011000101",
118338=>"001111111",
118339=>"001001000",
118340=>"000000000",
118341=>"100000011",
118342=>"010011000",
118343=>"111111111",
118344=>"100101001",
118345=>"101000110",
118346=>"001000110",
118347=>"100101001",
118348=>"000000100",
118349=>"101100100",
118350=>"001110000",
118351=>"101000000",
118352=>"111111111",
118353=>"101111111",
118354=>"011000111",
118355=>"011000010",
118356=>"101000101",
118357=>"110111111",
118358=>"001111101",
118359=>"000011001",
118360=>"001011111",
118361=>"000011010",
118362=>"100111000",
118363=>"011111100",
118364=>"010000000",
118365=>"001101111",
118366=>"111000101",
118367=>"100100001",
118368=>"111001010",
118369=>"111000111",
118370=>"000000111",
118371=>"011001011",
118372=>"101111011",
118373=>"011011110",
118374=>"111101001",
118375=>"000000000",
118376=>"110100101",
118377=>"011011111",
118378=>"111011000",
118379=>"011111001",
118380=>"111000111",
118381=>"111011100",
118382=>"001000101",
118383=>"000111010",
118384=>"100000110",
118385=>"100010010",
118386=>"110010010",
118387=>"101000000",
118388=>"011010000",
118389=>"000100010",
118390=>"010010000",
118391=>"100101101",
118392=>"000000111",
118393=>"000111110",
118394=>"110110001",
118395=>"101111111",
118396=>"111010011",
118397=>"101000111",
118398=>"010111111",
118399=>"100000101",
118400=>"111010001",
118401=>"000000100",
118402=>"000000000",
118403=>"000010100",
118404=>"111100000",
118405=>"100000000",
118406=>"110100100",
118407=>"010111111",
118408=>"111100101",
118409=>"110000000",
118410=>"011010011",
118411=>"000111111",
118412=>"010000000",
118413=>"010101111",
118414=>"111101111",
118415=>"000001111",
118416=>"111100000",
118417=>"010110000",
118418=>"111110000",
118419=>"010010011",
118420=>"101111011",
118421=>"000010110",
118422=>"000100111",
118423=>"100100000",
118424=>"010010111",
118425=>"001000001",
118426=>"100111101",
118427=>"000000111",
118428=>"110000100",
118429=>"111101111",
118430=>"111111000",
118431=>"100101000",
118432=>"111111100",
118433=>"000000101",
118434=>"101111011",
118435=>"111111100",
118436=>"101110000",
118437=>"100111001",
118438=>"011000000",
118439=>"010001000",
118440=>"000000010",
118441=>"111101111",
118442=>"000000000",
118443=>"000010010",
118444=>"000000000",
118445=>"000001011",
118446=>"010001011",
118447=>"010000000",
118448=>"101001111",
118449=>"011110100",
118450=>"101101111",
118451=>"100110001",
118452=>"111111111",
118453=>"011000010",
118454=>"110001001",
118455=>"011011000",
118456=>"011000110",
118457=>"110111010",
118458=>"111000000",
118459=>"110000000",
118460=>"011001101",
118461=>"111011000",
118462=>"000000011",
118463=>"000000000",
118464=>"111001001",
118465=>"010101101",
118466=>"111111000",
118467=>"111011010",
118468=>"000111000",
118469=>"101111101",
118470=>"010011000",
118471=>"011000111",
118472=>"000111111",
118473=>"101100100",
118474=>"111111111",
118475=>"000110000",
118476=>"011011101",
118477=>"100010110",
118478=>"101111110",
118479=>"110101111",
118480=>"001110101",
118481=>"111011110",
118482=>"000000010",
118483=>"110111000",
118484=>"000100110",
118485=>"000001101",
118486=>"000000011",
118487=>"010100111",
118488=>"010000000",
118489=>"000010010",
118490=>"001101000",
118491=>"101001111",
118492=>"010000011",
118493=>"100101101",
118494=>"101111000",
118495=>"011101010",
118496=>"110101101",
118497=>"001001010",
118498=>"111101000",
118499=>"111111000",
118500=>"010101101",
118501=>"100010000",
118502=>"100111111",
118503=>"010110100",
118504=>"111110111",
118505=>"111000011",
118506=>"000110100",
118507=>"110110000",
118508=>"000110000",
118509=>"010010000",
118510=>"101000000",
118511=>"000001010",
118512=>"000110010",
118513=>"011111100",
118514=>"010000000",
118515=>"001000110",
118516=>"110011011",
118517=>"111000000",
118518=>"000010110",
118519=>"001000110",
118520=>"111000000",
118521=>"011101111",
118522=>"101000000",
118523=>"111111110",
118524=>"010101111",
118525=>"000010000",
118526=>"001001000",
118527=>"010000001",
118528=>"001000100",
118529=>"000111111",
118530=>"000000111",
118531=>"000000001",
118532=>"101000000",
118533=>"000000110",
118534=>"111001000",
118535=>"010000001",
118536=>"000000010",
118537=>"111000000",
118538=>"110001100",
118539=>"000101101",
118540=>"000010111",
118541=>"111101000",
118542=>"000000000",
118543=>"011101111",
118544=>"111100000",
118545=>"011010011",
118546=>"000000111",
118547=>"000010000",
118548=>"111111111",
118549=>"101101111",
118550=>"011110000",
118551=>"111111100",
118552=>"111000101",
118553=>"001001000",
118554=>"011000000",
118555=>"000010110",
118556=>"111110000",
118557=>"000000000",
118558=>"000010110",
118559=>"000000001",
118560=>"011001001",
118561=>"000111100",
118562=>"100101001",
118563=>"000000010",
118564=>"000000011",
118565=>"010100001",
118566=>"000010010",
118567=>"010101001",
118568=>"000010011",
118569=>"111111010",
118570=>"010010000",
118571=>"100000101",
118572=>"001011011",
118573=>"011110110",
118574=>"001010111",
118575=>"100001101",
118576=>"111010000",
118577=>"000010110",
118578=>"101011000",
118579=>"101000000",
118580=>"111101000",
118581=>"001101000",
118582=>"111100000",
118583=>"001101100",
118584=>"000111111",
118585=>"000000111",
118586=>"000010011",
118587=>"110110011",
118588=>"011101001",
118589=>"111111110",
118590=>"000111101",
118591=>"111000000",
118592=>"111000011",
118593=>"111111101",
118594=>"000000010",
118595=>"011001000",
118596=>"000110111",
118597=>"101111000",
118598=>"001000001",
118599=>"001000111",
118600=>"111111100",
118601=>"011000000",
118602=>"001100000",
118603=>"001111000",
118604=>"000000111",
118605=>"000000110",
118606=>"000000011",
118607=>"101000110",
118608=>"101101000",
118609=>"000101000",
118610=>"110111111",
118611=>"001000000",
118612=>"111001001",
118613=>"101100000",
118614=>"100001000",
118615=>"111000000",
118616=>"111111111",
118617=>"000110110",
118618=>"001100110",
118619=>"000011011",
118620=>"000111110",
118621=>"000110110",
118622=>"101101111",
118623=>"110100001",
118624=>"111000000",
118625=>"111101000",
118626=>"000000111",
118627=>"000011001",
118628=>"000000001",
118629=>"011111001",
118630=>"111101000",
118631=>"000001111",
118632=>"000010000",
118633=>"001111000",
118634=>"001111111",
118635=>"100001101",
118636=>"110000111",
118637=>"111111000",
118638=>"001011111",
118639=>"001010000",
118640=>"001000111",
118641=>"000111111",
118642=>"010001100",
118643=>"111101000",
118644=>"010010110",
118645=>"000001001",
118646=>"011010000",
118647=>"101001000",
118648=>"000000010",
118649=>"000110111",
118650=>"000010111",
118651=>"110010010",
118652=>"001001001",
118653=>"000000000",
118654=>"001111111",
118655=>"000001101",
118656=>"111011000",
118657=>"000110000",
118658=>"111001011",
118659=>"111100111",
118660=>"000010111",
118661=>"111101000",
118662=>"110011000",
118663=>"110100000",
118664=>"100000010",
118665=>"001000101",
118666=>"111101000",
118667=>"001001111",
118668=>"000101011",
118669=>"011011101",
118670=>"000000011",
118671=>"000001000",
118672=>"000000110",
118673=>"000000111",
118674=>"101111001",
118675=>"000101111",
118676=>"111111000",
118677=>"010010000",
118678=>"100001000",
118679=>"000010000",
118680=>"110010011",
118681=>"000111111",
118682=>"010100000",
118683=>"000000000",
118684=>"000100001",
118685=>"000000000",
118686=>"001111101",
118687=>"000000010",
118688=>"101001111",
118689=>"111111100",
118690=>"000001001",
118691=>"000100110",
118692=>"000110111",
118693=>"001110110",
118694=>"001000001",
118695=>"011001001",
118696=>"111111000",
118697=>"011001000",
118698=>"000111111",
118699=>"000010111",
118700=>"111111111",
118701=>"000101111",
118702=>"100101100",
118703=>"111000000",
118704=>"001001110",
118705=>"000101100",
118706=>"000000000",
118707=>"000001011",
118708=>"100110000",
118709=>"000000000",
118710=>"000000000",
118711=>"000000011",
118712=>"110100100",
118713=>"111011001",
118714=>"110100001",
118715=>"000000111",
118716=>"011111110",
118717=>"000000001",
118718=>"001000010",
118719=>"111111010",
118720=>"000000100",
118721=>"000000111",
118722=>"111111000",
118723=>"000000010",
118724=>"100000001",
118725=>"100100110",
118726=>"000011011",
118727=>"000000011",
118728=>"101101101",
118729=>"000111011",
118730=>"101000000",
118731=>"000001110",
118732=>"000000000",
118733=>"110100100",
118734=>"111100100",
118735=>"010111101",
118736=>"000100101",
118737=>"011111100",
118738=>"001100000",
118739=>"000000101",
118740=>"000001111",
118741=>"110111001",
118742=>"011000011",
118743=>"110000000",
118744=>"000111111",
118745=>"000000000",
118746=>"001011011",
118747=>"011000000",
118748=>"100011100",
118749=>"001111110",
118750=>"000000000",
118751=>"110000010",
118752=>"000010010",
118753=>"000011011",
118754=>"001001101",
118755=>"011111111",
118756=>"000000001",
118757=>"000000100",
118758=>"001000111",
118759=>"000001011",
118760=>"000000010",
118761=>"111111100",
118762=>"110101101",
118763=>"111001000",
118764=>"000111000",
118765=>"000000100",
118766=>"000000000",
118767=>"000110111",
118768=>"111101100",
118769=>"000011011",
118770=>"111000000",
118771=>"001011011",
118772=>"100100000",
118773=>"000101111",
118774=>"000100000",
118775=>"000000110",
118776=>"000010000",
118777=>"000010000",
118778=>"000000110",
118779=>"111111100",
118780=>"000100001",
118781=>"000000000",
118782=>"001000110",
118783=>"100000000",
118784=>"101100110",
118785=>"110111101",
118786=>"100000100",
118787=>"000001000",
118788=>"001011011",
118789=>"111001001",
118790=>"000000111",
118791=>"111111101",
118792=>"000000001",
118793=>"110000000",
118794=>"011111011",
118795=>"110100101",
118796=>"000000010",
118797=>"000001111",
118798=>"111110100",
118799=>"000000110",
118800=>"010000000",
118801=>"011010000",
118802=>"000111111",
118803=>"000111101",
118804=>"101111111",
118805=>"101100000",
118806=>"111011111",
118807=>"101101000",
118808=>"000110111",
118809=>"001000010",
118810=>"000000000",
118811=>"111000000",
118812=>"000111101",
118813=>"011101000",
118814=>"000101000",
118815=>"011011000",
118816=>"010111111",
118817=>"100000000",
118818=>"001111111",
118819=>"101001111",
118820=>"000110111",
118821=>"000001001",
118822=>"000011000",
118823=>"100000110",
118824=>"010000000",
118825=>"000010000",
118826=>"000001001",
118827=>"101000100",
118828=>"000111111",
118829=>"111011011",
118830=>"100101001",
118831=>"000011110",
118832=>"111000000",
118833=>"011001111",
118834=>"000010100",
118835=>"010010000",
118836=>"000010111",
118837=>"111011001",
118838=>"110100100",
118839=>"111100000",
118840=>"101111111",
118841=>"111010110",
118842=>"101000111",
118843=>"101100101",
118844=>"001001111",
118845=>"111000101",
118846=>"001000000",
118847=>"000111001",
118848=>"111111111",
118849=>"000111101",
118850=>"011000000",
118851=>"100010001",
118852=>"000001111",
118853=>"000100000",
118854=>"110100111",
118855=>"000000110",
118856=>"011010010",
118857=>"111101101",
118858=>"100000001",
118859=>"001000000",
118860=>"010100111",
118861=>"011011010",
118862=>"110110011",
118863=>"001101100",
118864=>"011101000",
118865=>"101111111",
118866=>"111100000",
118867=>"110111000",
118868=>"000000100",
118869=>"010000000",
118870=>"110111111",
118871=>"000010000",
118872=>"000011001",
118873=>"110001011",
118874=>"111001000",
118875=>"000000011",
118876=>"111000010",
118877=>"101111110",
118878=>"111111111",
118879=>"100000001",
118880=>"000000000",
118881=>"110111100",
118882=>"111101101",
118883=>"001111010",
118884=>"111000011",
118885=>"111101111",
118886=>"101110011",
118887=>"010010101",
118888=>"000010010",
118889=>"101111111",
118890=>"110111111",
118891=>"000000000",
118892=>"100111111",
118893=>"111111000",
118894=>"000100111",
118895=>"000111111",
118896=>"011111110",
118897=>"101001000",
118898=>"001001001",
118899=>"000000000",
118900=>"000101111",
118901=>"100111111",
118902=>"010111001",
118903=>"000111111",
118904=>"000010111",
118905=>"000011111",
118906=>"111000000",
118907=>"110111111",
118908=>"000000011",
118909=>"000011011",
118910=>"100100000",
118911=>"100100100",
118912=>"110101111",
118913=>"000000100",
118914=>"111101011",
118915=>"101111111",
118916=>"010111000",
118917=>"111111110",
118918=>"000110001",
118919=>"011000000",
118920=>"110100111",
118921=>"110100000",
118922=>"100011001",
118923=>"000100000",
118924=>"011100000",
118925=>"000000010",
118926=>"100000000",
118927=>"111000001",
118928=>"000010100",
118929=>"000101101",
118930=>"000000000",
118931=>"000000000",
118932=>"110110000",
118933=>"111101001",
118934=>"001010111",
118935=>"010000000",
118936=>"001000001",
118937=>"000111111",
118938=>"111000000",
118939=>"110000010",
118940=>"111000010",
118941=>"000000000",
118942=>"100111111",
118943=>"111101101",
118944=>"011001111",
118945=>"010000000",
118946=>"101000000",
118947=>"000010111",
118948=>"101001000",
118949=>"010000100",
118950=>"100001101",
118951=>"011001111",
118952=>"000000000",
118953=>"100010001",
118954=>"100100011",
118955=>"000000000",
118956=>"100111111",
118957=>"111101111",
118958=>"011010001",
118959=>"111000000",
118960=>"000000000",
118961=>"110100100",
118962=>"000010000",
118963=>"000000011",
118964=>"000111111",
118965=>"111111010",
118966=>"000001011",
118967=>"000000000",
118968=>"100110111",
118969=>"011001000",
118970=>"000001000",
118971=>"000000000",
118972=>"111101111",
118973=>"000000101",
118974=>"100000001",
118975=>"011101111",
118976=>"010100101",
118977=>"111000000",
118978=>"000111001",
118979=>"111101101",
118980=>"101001111",
118981=>"111001001",
118982=>"100011010",
118983=>"111000001",
118984=>"111101000",
118985=>"100000000",
118986=>"111111110",
118987=>"110010000",
118988=>"111111111",
118989=>"111100100",
118990=>"010100101",
118991=>"000011111",
118992=>"011011100",
118993=>"111111110",
118994=>"000000000",
118995=>"000000010",
118996=>"101100111",
118997=>"001000001",
118998=>"010011111",
118999=>"010110010",
119000=>"101111000",
119001=>"010011000",
119002=>"110100111",
119003=>"101001000",
119004=>"100110110",
119005=>"000010011",
119006=>"001001001",
119007=>"000111011",
119008=>"000111000",
119009=>"111111000",
119010=>"010110111",
119011=>"010000000",
119012=>"000000111",
119013=>"001111111",
119014=>"000000000",
119015=>"000011111",
119016=>"000000000",
119017=>"011111101",
119018=>"000110110",
119019=>"011100000",
119020=>"000000000",
119021=>"000000111",
119022=>"000000010",
119023=>"111000111",
119024=>"100100111",
119025=>"110100000",
119026=>"101100101",
119027=>"011011111",
119028=>"010011011",
119029=>"111111000",
119030=>"000000010",
119031=>"111000000",
119032=>"000000011",
119033=>"111111111",
119034=>"010010110",
119035=>"111111111",
119036=>"101111111",
119037=>"010000000",
119038=>"111000110",
119039=>"111110100",
119040=>"110010000",
119041=>"000010111",
119042=>"001001001",
119043=>"111001000",
119044=>"000010001",
119045=>"100001111",
119046=>"001001001",
119047=>"000011000",
119048=>"110100110",
119049=>"000000010",
119050=>"001000000",
119051=>"000000001",
119052=>"001001011",
119053=>"100110110",
119054=>"000100010",
119055=>"110110001",
119056=>"100110000",
119057=>"110000110",
119058=>"000001111",
119059=>"000100110",
119060=>"110110001",
119061=>"000001001",
119062=>"100110111",
119063=>"110000110",
119064=>"000000000",
119065=>"100111110",
119066=>"000000000",
119067=>"101001000",
119068=>"010110001",
119069=>"001001110",
119070=>"110110100",
119071=>"011011000",
119072=>"110110010",
119073=>"010110001",
119074=>"111001000",
119075=>"110011100",
119076=>"100100000",
119077=>"110111001",
119078=>"110110000",
119079=>"001000100",
119080=>"010110000",
119081=>"110110010",
119082=>"100110110",
119083=>"000000111",
119084=>"001110111",
119085=>"101100110",
119086=>"110110111",
119087=>"110001001",
119088=>"111111000",
119089=>"100111100",
119090=>"111010110",
119091=>"111011110",
119092=>"110000000",
119093=>"001001111",
119094=>"100001011",
119095=>"000001001",
119096=>"110000010",
119097=>"001110110",
119098=>"000001101",
119099=>"111001001",
119100=>"100100100",
119101=>"111111001",
119102=>"000000000",
119103=>"110110111",
119104=>"110110001",
119105=>"110110000",
119106=>"110111000",
119107=>"111100000",
119108=>"011111111",
119109=>"110110100",
119110=>"000000110",
119111=>"111100000",
119112=>"110011111",
119113=>"110110010",
119114=>"010000011",
119115=>"010000010",
119116=>"110100010",
119117=>"000011000",
119118=>"001101100",
119119=>"001000110",
119120=>"011011010",
119121=>"100111110",
119122=>"001001111",
119123=>"111001100",
119124=>"011000110",
119125=>"010110110",
119126=>"011010000",
119127=>"101101000",
119128=>"000001001",
119129=>"110100111",
119130=>"101101001",
119131=>"011100110",
119132=>"000000000",
119133=>"000011010",
119134=>"110100000",
119135=>"110110110",
119136=>"110110110",
119137=>"110110110",
119138=>"001001001",
119139=>"110111000",
119140=>"010110000",
119141=>"100000110",
119142=>"110110000",
119143=>"001000010",
119144=>"110110110",
119145=>"111001001",
119146=>"100010110",
119147=>"111110101",
119148=>"010110000",
119149=>"001000001",
119150=>"111001101",
119151=>"000000000",
119152=>"000100110",
119153=>"110000001",
119154=>"010100110",
119155=>"111111110",
119156=>"010111010",
119157=>"000000000",
119158=>"010010000",
119159=>"110111000",
119160=>"001000110",
119161=>"111001000",
119162=>"001001000",
119163=>"000000001",
119164=>"000110110",
119165=>"110100100",
119166=>"001101111",
119167=>"110000100",
119168=>"011100000",
119169=>"110001000",
119170=>"110000110",
119171=>"010111100",
119172=>"000000110",
119173=>"111000101",
119174=>"010110010",
119175=>"000110001",
119176=>"111011010",
119177=>"111111111",
119178=>"001110011",
119179=>"111000000",
119180=>"000000001",
119181=>"001011111",
119182=>"100000000",
119183=>"011000000",
119184=>"010010000",
119185=>"111111001",
119186=>"001001000",
119187=>"111000001",
119188=>"000110100",
119189=>"000000110",
119190=>"110110000",
119191=>"000010000",
119192=>"000001000",
119193=>"001111110",
119194=>"001001110",
119195=>"100000001",
119196=>"001001110",
119197=>"000110110",
119198=>"001110110",
119199=>"101001001",
119200=>"001011111",
119201=>"100110110",
119202=>"110100000",
119203=>"010000111",
119204=>"111110000",
119205=>"000011000",
119206=>"011011011",
119207=>"000010000",
119208=>"001101110",
119209=>"000000110",
119210=>"001001111",
119211=>"001010010",
119212=>"110111101",
119213=>"110110110",
119214=>"000011011",
119215=>"001001111",
119216=>"110110000",
119217=>"011011000",
119218=>"111000000",
119219=>"011000000",
119220=>"110100110",
119221=>"111111111",
119222=>"000000101",
119223=>"000010101",
119224=>"011010011",
119225=>"001110110",
119226=>"010110010",
119227=>"111110110",
119228=>"001100000",
119229=>"111001111",
119230=>"000000100",
119231=>"101001011",
119232=>"100001101",
119233=>"001001111",
119234=>"111000001",
119235=>"100100100",
119236=>"101000000",
119237=>"100000001",
119238=>"010011000",
119239=>"000110101",
119240=>"100110110",
119241=>"000111000",
119242=>"010111111",
119243=>"000000000",
119244=>"000110111",
119245=>"000110110",
119246=>"111001000",
119247=>"100110010",
119248=>"111001011",
119249=>"100110100",
119250=>"110011110",
119251=>"011010111",
119252=>"100100101",
119253=>"010001000",
119254=>"000110000",
119255=>"000110110",
119256=>"001001111",
119257=>"000000000",
119258=>"000100000",
119259=>"001001001",
119260=>"011100100",
119261=>"001110111",
119262=>"010000000",
119263=>"110000010",
119264=>"001000001",
119265=>"100000001",
119266=>"001001101",
119267=>"011011000",
119268=>"001001000",
119269=>"001001111",
119270=>"110000011",
119271=>"010111110",
119272=>"000000111",
119273=>"011111110",
119274=>"010000001",
119275=>"000001000",
119276=>"001001011",
119277=>"001001111",
119278=>"000001000",
119279=>"000001000",
119280=>"001001111",
119281=>"011001000",
119282=>"000101110",
119283=>"000010110",
119284=>"110101011",
119285=>"011001001",
119286=>"011001010",
119287=>"110000110",
119288=>"101101111",
119289=>"001000111",
119290=>"111001101",
119291=>"011001000",
119292=>"110110000",
119293=>"001001001",
119294=>"100101000",
119295=>"000000000",
119296=>"111101110",
119297=>"000010001",
119298=>"100100101",
119299=>"000101101",
119300=>"110111100",
119301=>"100000001",
119302=>"100100100",
119303=>"111111011",
119304=>"111000100",
119305=>"000000010",
119306=>"010011000",
119307=>"000011011",
119308=>"000000111",
119309=>"101000110",
119310=>"101011111",
119311=>"011111000",
119312=>"011011000",
119313=>"000111101",
119314=>"111100000",
119315=>"000010111",
119316=>"000100001",
119317=>"011011000",
119318=>"100100000",
119319=>"000111110",
119320=>"110100000",
119321=>"011111010",
119322=>"101111010",
119323=>"101100111",
119324=>"100100001",
119325=>"101100000",
119326=>"111101101",
119327=>"000100000",
119328=>"101101011",
119329=>"100100000",
119330=>"011011111",
119331=>"000100100",
119332=>"110111100",
119333=>"010000110",
119334=>"111111010",
119335=>"100100000",
119336=>"110111111",
119337=>"000000000",
119338=>"000000110",
119339=>"101110111",
119340=>"101011111",
119341=>"000000011",
119342=>"011011000",
119343=>"111001000",
119344=>"011000000",
119345=>"100111111",
119346=>"000110010",
119347=>"010011011",
119348=>"011011000",
119349=>"101101011",
119350=>"001011011",
119351=>"101100011",
119352=>"011100001",
119353=>"101100000",
119354=>"010011100",
119355=>"111100111",
119356=>"001111001",
119357=>"011100010",
119358=>"000000000",
119359=>"110111011",
119360=>"111101000",
119361=>"000000010",
119362=>"111011000",
119363=>"001001101",
119364=>"000100101",
119365=>"000100011",
119366=>"011011011",
119367=>"100000101",
119368=>"000000110",
119369=>"101100111",
119370=>"101100100",
119371=>"011011001",
119372=>"101100111",
119373=>"001001001",
119374=>"001101110",
119375=>"100111110",
119376=>"000000111",
119377=>"111110100",
119378=>"110111100",
119379=>"100000100",
119380=>"000100000",
119381=>"011011101",
119382=>"001011111",
119383=>"111111000",
119384=>"101100100",
119385=>"000100110",
119386=>"000111000",
119387=>"011011000",
119388=>"010011010",
119389=>"100101000",
119390=>"111110111",
119391=>"100110000",
119392=>"000000111",
119393=>"000011000",
119394=>"000000001",
119395=>"100101111",
119396=>"100111110",
119397=>"100101110",
119398=>"111111110",
119399=>"100000000",
119400=>"011111000",
119401=>"100111011",
119402=>"001000110",
119403=>"010010000",
119404=>"011000000",
119405=>"011011000",
119406=>"010011010",
119407=>"001000100",
119408=>"111111001",
119409=>"011111100",
119410=>"011011000",
119411=>"100000000",
119412=>"010111111",
119413=>"100100111",
119414=>"101010010",
119415=>"000000111",
119416=>"001100111",
119417=>"000000000",
119418=>"001100010",
119419=>"000000100",
119420=>"111010100",
119421=>"001000100",
119422=>"110011010",
119423=>"101100101",
119424=>"101000111",
119425=>"111001000",
119426=>"011000111",
119427=>"000100000",
119428=>"100111011",
119429=>"000000110",
119430=>"111111101",
119431=>"001011000",
119432=>"110111101",
119433=>"011111010",
119434=>"011011011",
119435=>"000000111",
119436=>"100000000",
119437=>"111001011",
119438=>"001000000",
119439=>"000001000",
119440=>"001101011",
119441=>"101111111",
119442=>"100000100",
119443=>"000100100",
119444=>"010010011",
119445=>"101011001",
119446=>"011011010",
119447=>"110110100",
119448=>"011111111",
119449=>"111011010",
119450=>"000011111",
119451=>"000000000",
119452=>"100111111",
119453=>"010010011",
119454=>"010000000",
119455=>"100100111",
119456=>"100101100",
119457=>"111101111",
119458=>"011100100",
119459=>"101000111",
119460=>"011011000",
119461=>"111010001",
119462=>"111001011",
119463=>"111000000",
119464=>"000000011",
119465=>"000000100",
119466=>"000000111",
119467=>"100101011",
119468=>"110111110",
119469=>"100100011",
119470=>"001000011",
119471=>"000010011",
119472=>"000000111",
119473=>"000000011",
119474=>"100111000",
119475=>"000001001",
119476=>"001101010",
119477=>"010011001",
119478=>"101110111",
119479=>"100111111",
119480=>"101011010",
119481=>"000011010",
119482=>"111010000",
119483=>"001011011",
119484=>"000000010",
119485=>"011000110",
119486=>"101001111",
119487=>"000000000",
119488=>"011011000",
119489=>"111100000",
119490=>"011000111",
119491=>"011100000",
119492=>"110100111",
119493=>"110100001",
119494=>"111000011",
119495=>"111011100",
119496=>"010011011",
119497=>"001100100",
119498=>"001011111",
119499=>"001111101",
119500=>"111111011",
119501=>"001011111",
119502=>"010011110",
119503=>"000011111",
119504=>"011001011",
119505=>"000001001",
119506=>"011111000",
119507=>"111111111",
119508=>"001000110",
119509=>"111111100",
119510=>"100100101",
119511=>"011011011",
119512=>"100100111",
119513=>"100110010",
119514=>"001000001",
119515=>"111111111",
119516=>"100100101",
119517=>"110001001",
119518=>"001100110",
119519=>"000000011",
119520=>"000011000",
119521=>"000100100",
119522=>"000100000",
119523=>"111111100",
119524=>"000000000",
119525=>"011000011",
119526=>"100000110",
119527=>"000000100",
119528=>"100100000",
119529=>"000110011",
119530=>"010011010",
119531=>"111111100",
119532=>"101100100",
119533=>"111100111",
119534=>"101000110",
119535=>"000000000",
119536=>"100000011",
119537=>"101110100",
119538=>"000100000",
119539=>"000000101",
119540=>"110110011",
119541=>"001111100",
119542=>"000001111",
119543=>"000000100",
119544=>"001011110",
119545=>"111001000",
119546=>"011111111",
119547=>"111011010",
119548=>"011011000",
119549=>"100100000",
119550=>"011110110",
119551=>"010011101",
119552=>"100000110",
119553=>"111000000",
119554=>"011010000",
119555=>"101101001",
119556=>"000011011",
119557=>"111101001",
119558=>"100000001",
119559=>"001111011",
119560=>"000000000",
119561=>"000000001",
119562=>"000111111",
119563=>"101101111",
119564=>"000001001",
119565=>"001000111",
119566=>"100111001",
119567=>"110111111",
119568=>"101110111",
119569=>"110010010",
119570=>"111110000",
119571=>"000101010",
119572=>"000000000",
119573=>"111110110",
119574=>"011011111",
119575=>"000100111",
119576=>"010000000",
119577=>"111110000",
119578=>"110000000",
119579=>"100111011",
119580=>"101000000",
119581=>"001001101",
119582=>"111111000",
119583=>"000000001",
119584=>"000000000",
119585=>"111101000",
119586=>"000000000",
119587=>"111001001",
119588=>"000000111",
119589=>"001001011",
119590=>"000000101",
119591=>"010001000",
119592=>"000001000",
119593=>"000000101",
119594=>"100110110",
119595=>"000000000",
119596=>"011111111",
119597=>"111110101",
119598=>"010011011",
119599=>"000000000",
119600=>"000000000",
119601=>"110110111",
119602=>"011000001",
119603=>"111011010",
119604=>"001000100",
119605=>"000001110",
119606=>"011001001",
119607=>"000000000",
119608=>"111011011",
119609=>"101000101",
119610=>"000000000",
119611=>"000000000",
119612=>"000000001",
119613=>"110111000",
119614=>"000000000",
119615=>"000001001",
119616=>"110110101",
119617=>"110010110",
119618=>"110111000",
119619=>"111111000",
119620=>"100111111",
119621=>"000001111",
119622=>"000101000",
119623=>"110000110",
119624=>"001011101",
119625=>"111111111",
119626=>"111001011",
119627=>"011111111",
119628=>"111011001",
119629=>"101100011",
119630=>"011111000",
119631=>"010011111",
119632=>"011010111",
119633=>"111010010",
119634=>"000001101",
119635=>"000000101",
119636=>"101101111",
119637=>"001111111",
119638=>"000011000",
119639=>"000111111",
119640=>"111111110",
119641=>"100100110",
119642=>"100101100",
119643=>"110111111",
119644=>"111111011",
119645=>"000000000",
119646=>"010110010",
119647=>"011010010",
119648=>"000000001",
119649=>"010111111",
119650=>"000000001",
119651=>"001111001",
119652=>"011001001",
119653=>"001011010",
119654=>"001001101",
119655=>"000000001",
119656=>"000100111",
119657=>"000000001",
119658=>"001101000",
119659=>"010101110",
119660=>"000000000",
119661=>"110111110",
119662=>"001000001",
119663=>"111011000",
119664=>"011111101",
119665=>"000001000",
119666=>"111000110",
119667=>"000000010",
119668=>"000101111",
119669=>"100000101",
119670=>"000111110",
119671=>"000000001",
119672=>"100000000",
119673=>"010010000",
119674=>"010000111",
119675=>"111101101",
119676=>"010000001",
119677=>"000000000",
119678=>"000000011",
119679=>"011111111",
119680=>"010101010",
119681=>"111111010",
119682=>"000000000",
119683=>"000111101",
119684=>"101000000",
119685=>"001001111",
119686=>"000000011",
119687=>"110010001",
119688=>"111111001",
119689=>"000000100",
119690=>"011111111",
119691=>"101101111",
119692=>"001001001",
119693=>"111111111",
119694=>"111111010",
119695=>"001000101",
119696=>"001000100",
119697=>"101111101",
119698=>"001100111",
119699=>"111000101",
119700=>"111001011",
119701=>"010000000",
119702=>"111111111",
119703=>"001001111",
119704=>"101111111",
119705=>"000000000",
119706=>"111111111",
119707=>"000000000",
119708=>"101001111",
119709=>"111111111",
119710=>"111111111",
119711=>"000001111",
119712=>"101111011",
119713=>"111111011",
119714=>"101000001",
119715=>"101111100",
119716=>"000111110",
119717=>"001101111",
119718=>"010101001",
119719=>"111011110",
119720=>"111111111",
119721=>"111001001",
119722=>"100001001",
119723=>"111101001",
119724=>"000000000",
119725=>"111001011",
119726=>"010111011",
119727=>"000111111",
119728=>"101000000",
119729=>"011110100",
119730=>"001000000",
119731=>"111001001",
119732=>"110111111",
119733=>"000000000",
119734=>"000000100",
119735=>"101000000",
119736=>"100000010",
119737=>"011010100",
119738=>"101001000",
119739=>"111010000",
119740=>"000001011",
119741=>"111110010",
119742=>"000000100",
119743=>"000000001",
119744=>"010010010",
119745=>"000110111",
119746=>"010111111",
119747=>"110001000",
119748=>"101001111",
119749=>"110110011",
119750=>"000101000",
119751=>"010111011",
119752=>"100100101",
119753=>"100110011",
119754=>"000000011",
119755=>"000001111",
119756=>"100000100",
119757=>"010000000",
119758=>"000000000",
119759=>"000000101",
119760=>"110100111",
119761=>"110111111",
119762=>"111010000",
119763=>"001001000",
119764=>"001000001",
119765=>"000000010",
119766=>"111111010",
119767=>"110110110",
119768=>"000000111",
119769=>"000001100",
119770=>"110011111",
119771=>"101101111",
119772=>"110111001",
119773=>"110001000",
119774=>"011100010",
119775=>"011000010",
119776=>"000000101",
119777=>"101001111",
119778=>"111111111",
119779=>"011111111",
119780=>"000000001",
119781=>"001001011",
119782=>"000000111",
119783=>"000110110",
119784=>"001000101",
119785=>"011010000",
119786=>"000101100",
119787=>"000000111",
119788=>"001000000",
119789=>"001101111",
119790=>"110110000",
119791=>"001000001",
119792=>"011001000",
119793=>"011111100",
119794=>"001001000",
119795=>"001011111",
119796=>"001011011",
119797=>"010111000",
119798=>"010000110",
119799=>"000000111",
119800=>"000000111",
119801=>"101111111",
119802=>"000010000",
119803=>"011010010",
119804=>"111111111",
119805=>"111101111",
119806=>"100100100",
119807=>"010011000",
119808=>"101101101",
119809=>"000011010",
119810=>"111001011",
119811=>"111011010",
119812=>"100111110",
119813=>"011001101",
119814=>"100100000",
119815=>"000100100",
119816=>"110100010",
119817=>"000000000",
119818=>"001101100",
119819=>"111011001",
119820=>"000110110",
119821=>"110011000",
119822=>"100100100",
119823=>"100100000",
119824=>"110101100",
119825=>"100000100",
119826=>"110000111",
119827=>"000001001",
119828=>"011001011",
119829=>"111001001",
119830=>"111001111",
119831=>"000100100",
119832=>"110000000",
119833=>"011001100",
119834=>"000001001",
119835=>"111001000",
119836=>"001000100",
119837=>"000000010",
119838=>"011011010",
119839=>"001111100",
119840=>"011111111",
119841=>"000001111",
119842=>"000001001",
119843=>"100110110",
119844=>"011111110",
119845=>"011001110",
119846=>"011011011",
119847=>"000110110",
119848=>"111011001",
119849=>"011011011",
119850=>"111110010",
119851=>"011001000",
119852=>"000110101",
119853=>"100010001",
119854=>"011011000",
119855=>"001000101",
119856=>"010000000",
119857=>"111001001",
119858=>"000011011",
119859=>"000111110",
119860=>"110001100",
119861=>"100100011",
119862=>"101001001",
119863=>"110110000",
119864=>"001001011",
119865=>"000000110",
119866=>"010001011",
119867=>"010100000",
119868=>"000000000",
119869=>"111110100",
119870=>"000001001",
119871=>"100110001",
119872=>"000000111",
119873=>"011111011",
119874=>"111011100",
119875=>"111101100",
119876=>"001000000",
119877=>"011111001",
119878=>"100110110",
119879=>"111110111",
119880=>"100111010",
119881=>"110000000",
119882=>"101001110",
119883=>"100110100",
119884=>"011001001",
119885=>"000000000",
119886=>"010010111",
119887=>"000111101",
119888=>"101001001",
119889=>"110001110",
119890=>"001100101",
119891=>"000101000",
119892=>"011001011",
119893=>"111101111",
119894=>"000000000",
119895=>"011111110",
119896=>"111011111",
119897=>"001101001",
119898=>"010100011",
119899=>"001001000",
119900=>"110110110",
119901=>"001000100",
119902=>"001001111",
119903=>"100011001",
119904=>"011111111",
119905=>"111011001",
119906=>"001001011",
119907=>"101100000",
119908=>"001000000",
119909=>"101111111",
119910=>"111011000",
119911=>"010110010",
119912=>"011001001",
119913=>"000000110",
119914=>"110000000",
119915=>"110110111",
119916=>"001110111",
119917=>"000100100",
119918=>"111001001",
119919=>"001001000",
119920=>"111111111",
119921=>"010010010",
119922=>"101001011",
119923=>"100111100",
119924=>"110100000",
119925=>"110010000",
119926=>"000011001",
119927=>"011001011",
119928=>"011010011",
119929=>"101000100",
119930=>"001000001",
119931=>"000000101",
119932=>"000001110",
119933=>"010000000",
119934=>"110001001",
119935=>"101110100",
119936=>"011100000",
119937=>"111000011",
119938=>"111101110",
119939=>"011111000",
119940=>"000001111",
119941=>"011011001",
119942=>"011011010",
119943=>"000100110",
119944=>"000100100",
119945=>"110100110",
119946=>"011000001",
119947=>"001110100",
119948=>"111001000",
119949=>"100000000",
119950=>"000110100",
119951=>"000000100",
119952=>"011111001",
119953=>"111011010",
119954=>"010010111",
119955=>"110001110",
119956=>"010000010",
119957=>"111001111",
119958=>"000000101",
119959=>"000000000",
119960=>"110011100",
119961=>"011011011",
119962=>"001001001",
119963=>"010001011",
119964=>"111010000",
119965=>"110101100",
119966=>"111000000",
119967=>"011100000",
119968=>"001111111",
119969=>"111110011",
119970=>"001111110",
119971=>"110000001",
119972=>"011011111",
119973=>"000100000",
119974=>"000111000",
119975=>"000101111",
119976=>"111000000",
119977=>"110010001",
119978=>"001001011",
119979=>"111011011",
119980=>"000111111",
119981=>"100100100",
119982=>"001001111",
119983=>"011110000",
119984=>"110000001",
119985=>"011111010",
119986=>"000011000",
119987=>"000011100",
119988=>"111111111",
119989=>"110101111",
119990=>"011011001",
119991=>"011011110",
119992=>"000111111",
119993=>"000000000",
119994=>"111010000",
119995=>"111111000",
119996=>"000111110",
119997=>"111001000",
119998=>"011111111",
119999=>"100000000",
120000=>"111000000",
120001=>"000000100",
120002=>"010011000",
120003=>"000000100",
120004=>"000110100",
120005=>"100001010",
120006=>"000100110",
120007=>"110000010",
120008=>"000110111",
120009=>"011010000",
120010=>"110111111",
120011=>"011001011",
120012=>"111111000",
120013=>"100100101",
120014=>"100000001",
120015=>"000000111",
120016=>"101001000",
120017=>"110111111",
120018=>"100000100",
120019=>"101111111",
120020=>"110000100",
120021=>"001001001",
120022=>"011000100",
120023=>"110000000",
120024=>"100110100",
120025=>"010010010",
120026=>"000000001",
120027=>"101101110",
120028=>"111011111",
120029=>"001011001",
120030=>"001010110",
120031=>"011011110",
120032=>"011010101",
120033=>"001000000",
120034=>"111000000",
120035=>"001111011",
120036=>"110000100",
120037=>"000100100",
120038=>"110111100",
120039=>"110110110",
120040=>"001001001",
120041=>"011001001",
120042=>"010000010",
120043=>"111111001",
120044=>"110000000",
120045=>"110000000",
120046=>"100000100",
120047=>"100110100",
120048=>"100000001",
120049=>"000101101",
120050=>"111011000",
120051=>"100000000",
120052=>"101100000",
120053=>"001011111",
120054=>"000110110",
120055=>"000001001",
120056=>"111011001",
120057=>"100011000",
120058=>"111001111",
120059=>"000010101",
120060=>"001001111",
120061=>"000100100",
120062=>"000110100",
120063=>"110110110",
120064=>"111000000",
120065=>"000101101",
120066=>"000110111",
120067=>"010100111",
120068=>"111111111",
120069=>"111111101",
120070=>"111111000",
120071=>"000000110",
120072=>"111110000",
120073=>"000000111",
120074=>"000000100",
120075=>"111111000",
120076=>"000111111",
120077=>"111111111",
120078=>"100000010",
120079=>"101110011",
120080=>"111101111",
120081=>"001000101",
120082=>"100101001",
120083=>"101000011",
120084=>"011111000",
120085=>"010010001",
120086=>"111001100",
120087=>"001000011",
120088=>"001000000",
120089=>"101111111",
120090=>"101010010",
120091=>"010101100",
120092=>"101101000",
120093=>"000010100",
120094=>"101111000",
120095=>"100100010",
120096=>"111101111",
120097=>"011111001",
120098=>"000000010",
120099=>"000010111",
120100=>"000000011",
120101=>"011111001",
120102=>"000100111",
120103=>"011111011",
120104=>"010010001",
120105=>"110100111",
120106=>"111000100",
120107=>"000100100",
120108=>"000000000",
120109=>"010100110",
120110=>"101000100",
120111=>"110001001",
120112=>"000000101",
120113=>"011101111",
120114=>"011001000",
120115=>"111010000",
120116=>"111100000",
120117=>"110111110",
120118=>"101000100",
120119=>"111010001",
120120=>"111000010",
120121=>"000010010",
120122=>"000000000",
120123=>"000000000",
120124=>"001001010",
120125=>"111111000",
120126=>"100000000",
120127=>"111111001",
120128=>"100100110",
120129=>"101101111",
120130=>"001101111",
120131=>"110110111",
120132=>"101111001",
120133=>"000100000",
120134=>"101001110",
120135=>"011000010",
120136=>"101001001",
120137=>"011111101",
120138=>"000000000",
120139=>"111101101",
120140=>"000010111",
120141=>"000001111",
120142=>"010101111",
120143=>"000000110",
120144=>"101000001",
120145=>"011000000",
120146=>"111111101",
120147=>"110100101",
120148=>"111000000",
120149=>"111011101",
120150=>"001000001",
120151=>"000000000",
120152=>"111110101",
120153=>"010001111",
120154=>"000010110",
120155=>"100100110",
120156=>"111111111",
120157=>"001001001",
120158=>"110011110",
120159=>"011011001",
120160=>"010011111",
120161=>"111011000",
120162=>"000011111",
120163=>"001000001",
120164=>"100100110",
120165=>"100101111",
120166=>"010010000",
120167=>"010010111",
120168=>"111000000",
120169=>"111000000",
120170=>"010000111",
120171=>"110111010",
120172=>"111011110",
120173=>"000000101",
120174=>"000000111",
120175=>"001001000",
120176=>"110101100",
120177=>"111000000",
120178=>"101000001",
120179=>"010111100",
120180=>"001000000",
120181=>"000000000",
120182=>"000000000",
120183=>"101110111",
120184=>"001010000",
120185=>"101101110",
120186=>"010101111",
120187=>"010101001",
120188=>"001101010",
120189=>"001000100",
120190=>"011010001",
120191=>"111111000",
120192=>"000010110",
120193=>"101100100",
120194=>"110111001",
120195=>"100111111",
120196=>"010000000",
120197=>"110101111",
120198=>"100110110",
120199=>"000000011",
120200=>"001111001",
120201=>"001001000",
120202=>"111100110",
120203=>"000001000",
120204=>"011010011",
120205=>"100000011",
120206=>"000111011",
120207=>"000000000",
120208=>"111100110",
120209=>"111101001",
120210=>"000110000",
120211=>"111101000",
120212=>"111001000",
120213=>"111000000",
120214=>"111011110",
120215=>"000011000",
120216=>"001000010",
120217=>"100000001",
120218=>"110010111",
120219=>"111111000",
120220=>"000001101",
120221=>"000000011",
120222=>"010000111",
120223=>"001000100",
120224=>"011110111",
120225=>"001110001",
120226=>"011011010",
120227=>"111000000",
120228=>"111010000",
120229=>"000001111",
120230=>"000110011",
120231=>"001011000",
120232=>"111011010",
120233=>"000111100",
120234=>"011000111",
120235=>"111000000",
120236=>"111010011",
120237=>"100000000",
120238=>"001001100",
120239=>"010111111",
120240=>"011111101",
120241=>"011100101",
120242=>"001001001",
120243=>"000100100",
120244=>"001100110",
120245=>"000011111",
120246=>"000010111",
120247=>"000111111",
120248=>"110000100",
120249=>"011100100",
120250=>"111111001",
120251=>"011000000",
120252=>"000010100",
120253=>"111111111",
120254=>"001011000",
120255=>"011000000",
120256=>"001001011",
120257=>"110000000",
120258=>"101000111",
120259=>"111100100",
120260=>"000110010",
120261=>"110100001",
120262=>"110101101",
120263=>"000010000",
120264=>"010000111",
120265=>"000000010",
120266=>"101111111",
120267=>"101101111",
120268=>"011011011",
120269=>"110001000",
120270=>"101000000",
120271=>"111111011",
120272=>"100111000",
120273=>"110111010",
120274=>"010011110",
120275=>"101101101",
120276=>"010101101",
120277=>"100100100",
120278=>"101001000",
120279=>"011001001",
120280=>"000000000",
120281=>"000111010",
120282=>"000101111",
120283=>"000000100",
120284=>"111001100",
120285=>"111010010",
120286=>"000011000",
120287=>"110011001",
120288=>"000000000",
120289=>"111000000",
120290=>"000011111",
120291=>"011001101",
120292=>"001001001",
120293=>"111001011",
120294=>"111111010",
120295=>"110000011",
120296=>"011101001",
120297=>"111011000",
120298=>"000001001",
120299=>"010000000",
120300=>"000000000",
120301=>"000010111",
120302=>"000000000",
120303=>"000100001",
120304=>"111011000",
120305=>"011001100",
120306=>"000000000",
120307=>"110101101",
120308=>"011000101",
120309=>"000000011",
120310=>"000000000",
120311=>"101000001",
120312=>"000000000",
120313=>"001000000",
120314=>"001100101",
120315=>"000101111",
120316=>"110001011",
120317=>"000000000",
120318=>"110111111",
120319=>"000000000",
120320=>"000101111",
120321=>"111111100",
120322=>"110000110",
120323=>"111001000",
120324=>"000110011",
120325=>"011001001",
120326=>"011101101",
120327=>"000000000",
120328=>"100001011",
120329=>"000000100",
120330=>"111000100",
120331=>"000000000",
120332=>"000001001",
120333=>"110110110",
120334=>"111000000",
120335=>"111011111",
120336=>"111000010",
120337=>"111001010",
120338=>"001001000",
120339=>"111111000",
120340=>"101000010",
120341=>"111110100",
120342=>"001111110",
120343=>"111011111",
120344=>"101000110",
120345=>"100111001",
120346=>"101100101",
120347=>"000111011",
120348=>"110110111",
120349=>"110110000",
120350=>"000000011",
120351=>"111101111",
120352=>"000000110",
120353=>"000100011",
120354=>"101111110",
120355=>"101111101",
120356=>"101101100",
120357=>"011111100",
120358=>"011011110",
120359=>"000000000",
120360=>"111110111",
120361=>"000110110",
120362=>"111000101",
120363=>"101111001",
120364=>"010000000",
120365=>"000000000",
120366=>"100001001",
120367=>"110011011",
120368=>"111100000",
120369=>"000001001",
120370=>"111011010",
120371=>"110110000",
120372=>"010111111",
120373=>"000010001",
120374=>"010110101",
120375=>"000101111",
120376=>"000000000",
120377=>"001001100",
120378=>"111001000",
120379=>"101110000",
120380=>"100110000",
120381=>"101111111",
120382=>"001001100",
120383=>"100010001",
120384=>"111011111",
120385=>"111111000",
120386=>"000000000",
120387=>"010110111",
120388=>"101000000",
120389=>"111101001",
120390=>"010001101",
120391=>"110110011",
120392=>"000000000",
120393=>"001111011",
120394=>"001100100",
120395=>"111001111",
120396=>"100000000",
120397=>"011010011",
120398=>"101001110",
120399=>"110010000",
120400=>"101110111",
120401=>"110111111",
120402=>"110101000",
120403=>"111011000",
120404=>"000110010",
120405=>"010000100",
120406=>"111110111",
120407=>"000100110",
120408=>"110101111",
120409=>"111001000",
120410=>"000001001",
120411=>"010000000",
120412=>"111001000",
120413=>"111000100",
120414=>"111110010",
120415=>"000111111",
120416=>"111111111",
120417=>"001000001",
120418=>"111000000",
120419=>"001111110",
120420=>"000000010",
120421=>"001110010",
120422=>"110100010",
120423=>"100110110",
120424=>"001111110",
120425=>"111101000",
120426=>"000000000",
120427=>"111110010",
120428=>"111000000",
120429=>"011000001",
120430=>"000001101",
120431=>"101111001",
120432=>"111010100",
120433=>"000000000",
120434=>"010011111",
120435=>"001001000",
120436=>"111001101",
120437=>"111001101",
120438=>"000100000",
120439=>"010010010",
120440=>"110110100",
120441=>"000111000",
120442=>"101000011",
120443=>"111001101",
120444=>"001000000",
120445=>"101111001",
120446=>"111010110",
120447=>"111000111",
120448=>"100110111",
120449=>"111100110",
120450=>"111111111",
120451=>"101000010",
120452=>"111101000",
120453=>"111000001",
120454=>"110111001",
120455=>"000000010",
120456=>"011011011",
120457=>"111000110",
120458=>"111100111",
120459=>"101110000",
120460=>"000110111",
120461=>"000000111",
120462=>"111001000",
120463=>"110001001",
120464=>"001101101",
120465=>"000101110",
120466=>"111101101",
120467=>"010110010",
120468=>"000000100",
120469=>"001000000",
120470=>"111111000",
120471=>"110001000",
120472=>"010000000",
120473=>"111011000",
120474=>"111010000",
120475=>"000000000",
120476=>"000001001",
120477=>"000000000",
120478=>"000000110",
120479=>"111100000",
120480=>"000000011",
120481=>"000111111",
120482=>"111001010",
120483=>"001000000",
120484=>"000000111",
120485=>"001000110",
120486=>"111111010",
120487=>"000000000",
120488=>"101101010",
120489=>"000101101",
120490=>"101000111",
120491=>"111011011",
120492=>"110111111",
120493=>"110000000",
120494=>"010111110",
120495=>"111001001",
120496=>"001000111",
120497=>"111101100",
120498=>"111000001",
120499=>"001001001",
120500=>"111000110",
120501=>"010111110",
120502=>"001111111",
120503=>"000011000",
120504=>"001011001",
120505=>"001000000",
120506=>"010111111",
120507=>"110101110",
120508=>"111110001",
120509=>"111001001",
120510=>"011000100",
120511=>"000101011",
120512=>"000110111",
120513=>"101000001",
120514=>"110111111",
120515=>"101111101",
120516=>"010000001",
120517=>"000000110",
120518=>"000000100",
120519=>"000110101",
120520=>"110000000",
120521=>"001111111",
120522=>"111101111",
120523=>"111000010",
120524=>"000000010",
120525=>"000000010",
120526=>"000101011",
120527=>"111001101",
120528=>"111111110",
120529=>"011001111",
120530=>"111001000",
120531=>"111111111",
120532=>"111111100",
120533=>"001011111",
120534=>"000001011",
120535=>"001001010",
120536=>"010011000",
120537=>"111000001",
120538=>"001011101",
120539=>"111000000",
120540=>"100111110",
120541=>"101101001",
120542=>"010100101",
120543=>"000110000",
120544=>"000000000",
120545=>"000000010",
120546=>"010110111",
120547=>"111000001",
120548=>"000010110",
120549=>"111001111",
120550=>"001000001",
120551=>"000111111",
120552=>"110101101",
120553=>"111111111",
120554=>"110000001",
120555=>"000101001",
120556=>"101000000",
120557=>"000010000",
120558=>"111000001",
120559=>"110000011",
120560=>"010111010",
120561=>"000000001",
120562=>"000000000",
120563=>"111100001",
120564=>"000001001",
120565=>"101000110",
120566=>"000000001",
120567=>"010010000",
120568=>"000000000",
120569=>"001101110",
120570=>"111110111",
120571=>"000000001",
120572=>"000111101",
120573=>"011100001",
120574=>"000100000",
120575=>"110000000",
120576=>"110100110",
120577=>"110110110",
120578=>"001001011",
120579=>"110100000",
120580=>"010110110",
120581=>"100110100",
120582=>"001001011",
120583=>"000001010",
120584=>"100100110",
120585=>"001001000",
120586=>"001001111",
120587=>"000000000",
120588=>"110011011",
120589=>"100001000",
120590=>"111001001",
120591=>"001010001",
120592=>"000110100",
120593=>"000001100",
120594=>"000000011",
120595=>"111000000",
120596=>"000001011",
120597=>"001011110",
120598=>"100100110",
120599=>"100000000",
120600=>"011011111",
120601=>"100000100",
120602=>"100110100",
120603=>"011011111",
120604=>"000011110",
120605=>"010010011",
120606=>"011011111",
120607=>"011000111",
120608=>"111000100",
120609=>"100100101",
120610=>"110011011",
120611=>"110110000",
120612=>"111111101",
120613=>"001001011",
120614=>"110110000",
120615=>"011011001",
120616=>"100100000",
120617=>"000100100",
120618=>"011000000",
120619=>"100110100",
120620=>"110111101",
120621=>"001011111",
120622=>"100100111",
120623=>"110011110",
120624=>"000110110",
120625=>"101100001",
120626=>"001111110",
120627=>"011011001",
120628=>"011001011",
120629=>"101010000",
120630=>"001101110",
120631=>"011101000",
120632=>"011001001",
120633=>"011001011",
120634=>"000001100",
120635=>"000011000",
120636=>"001011111",
120637=>"101101000",
120638=>"100001001",
120639=>"100100110",
120640=>"000000111",
120641=>"000111001",
120642=>"111111000",
120643=>"000110010",
120644=>"100100100",
120645=>"111011010",
120646=>"011011001",
120647=>"100101001",
120648=>"110010111",
120649=>"101001001",
120650=>"001011111",
120651=>"011011111",
120652=>"110000100",
120653=>"100000010",
120654=>"110010001",
120655=>"011011101",
120656=>"100100001",
120657=>"100110110",
120658=>"100001001",
120659=>"010000000",
120660=>"001001001",
120661=>"001011101",
120662=>"111111101",
120663=>"000001111",
120664=>"011001001",
120665=>"011001001",
120666=>"011011111",
120667=>"110101010",
120668=>"100100000",
120669=>"000110100",
120670=>"101111111",
120671=>"000100000",
120672=>"100100100",
120673=>"100100110",
120674=>"000001011",
120675=>"011011110",
120676=>"011001011",
120677=>"001001001",
120678=>"011011011",
120679=>"101101001",
120680=>"100101100",
120681=>"110011111",
120682=>"100111100",
120683=>"100111010",
120684=>"100100010",
120685=>"001100111",
120686=>"000001100",
120687=>"000011111",
120688=>"110010011",
120689=>"010000101",
120690=>"110011001",
120691=>"110110110",
120692=>"111111100",
120693=>"011011110",
120694=>"111010101",
120695=>"100101011",
120696=>"000000100",
120697=>"111110111",
120698=>"000001000",
120699=>"110101100",
120700=>"001001011",
120701=>"100000000",
120702=>"111101101",
120703=>"000011111",
120704=>"110110110",
120705=>"000000100",
120706=>"100000111",
120707=>"110010001",
120708=>"000011111",
120709=>"000000000",
120710=>"100110111",
120711=>"000000000",
120712=>"000000000",
120713=>"011011111",
120714=>"000000001",
120715=>"110000000",
120716=>"000100100",
120717=>"011000111",
120718=>"001011011",
120719=>"011001000",
120720=>"011001010",
120721=>"111011110",
120722=>"001001100",
120723=>"010011011",
120724=>"000010000",
120725=>"011111111",
120726=>"001001101",
120727=>"110110100",
120728=>"110001011",
120729=>"000100110",
120730=>"011011000",
120731=>"000100100",
120732=>"011000000",
120733=>"011011110",
120734=>"101000101",
120735=>"011001011",
120736=>"110110001",
120737=>"000101100",
120738=>"100011001",
120739=>"011010100",
120740=>"100011100",
120741=>"100000000",
120742=>"110100000",
120743=>"111100000",
120744=>"000010111",
120745=>"010100000",
120746=>"011001110",
120747=>"001101011",
120748=>"100100000",
120749=>"100100111",
120750=>"001011111",
120751=>"101100001",
120752=>"010110001",
120753=>"111110111",
120754=>"000011110",
120755=>"001001111",
120756=>"111111100",
120757=>"111011000",
120758=>"100111000",
120759=>"110001011",
120760=>"110100100",
120761=>"100010000",
120762=>"100000000",
120763=>"111000001",
120764=>"100000000",
120765=>"100100110",
120766=>"100100000",
120767=>"111111110",
120768=>"001001111",
120769=>"001000001",
120770=>"001111100",
120771=>"010000000",
120772=>"001010010",
120773=>"111111111",
120774=>"111000000",
120775=>"000100111",
120776=>"110000001",
120777=>"111110000",
120778=>"100010110",
120779=>"011011110",
120780=>"001001011",
120781=>"101000001",
120782=>"001001001",
120783=>"100100000",
120784=>"011001001",
120785=>"000100000",
120786=>"100010001",
120787=>"100110110",
120788=>"011000111",
120789=>"001000100",
120790=>"111000011",
120791=>"000111101",
120792=>"011001011",
120793=>"110010100",
120794=>"000000001",
120795=>"001001010",
120796=>"001010111",
120797=>"100110100",
120798=>"110110100",
120799=>"001001011",
120800=>"100100101",
120801=>"011011011",
120802=>"000000011",
120803=>"111110100",
120804=>"000000000",
120805=>"110110110",
120806=>"100100100",
120807=>"100011111",
120808=>"100100110",
120809=>"111010110",
120810=>"001001011",
120811=>"100010011",
120812=>"110110100",
120813=>"100100000",
120814=>"000010100",
120815=>"110110010",
120816=>"110110100",
120817=>"010010000",
120818=>"101011010",
120819=>"100100010",
120820=>"110001001",
120821=>"011001001",
120822=>"010000100",
120823=>"000100010",
120824=>"001001111",
120825=>"010011100",
120826=>"100000010",
120827=>"011110010",
120828=>"001001011",
120829=>"100110000",
120830=>"011111011",
120831=>"001001011",
120832=>"011011000",
120833=>"111111111",
120834=>"101000101",
120835=>"101100111",
120836=>"111111100",
120837=>"011101011",
120838=>"111100111",
120839=>"100000000",
120840=>"000110110",
120841=>"001000101",
120842=>"111000111",
120843=>"110101111",
120844=>"000111011",
120845=>"011111000",
120846=>"110001011",
120847=>"000000000",
120848=>"010011111",
120849=>"001000101",
120850=>"100101101",
120851=>"001111111",
120852=>"111001111",
120853=>"000110000",
120854=>"000000001",
120855=>"111000000",
120856=>"110100100",
120857=>"000111110",
120858=>"011100010",
120859=>"000001011",
120860=>"000000000",
120861=>"110110010",
120862=>"110011111",
120863=>"000110000",
120864=>"001000001",
120865=>"111111111",
120866=>"100100111",
120867=>"111110000",
120868=>"110101100",
120869=>"110100000",
120870=>"110111011",
120871=>"111010101",
120872=>"111011000",
120873=>"000000000",
120874=>"111100100",
120875=>"000001110",
120876=>"000000100",
120877=>"111111111",
120878=>"111001101",
120879=>"000111011",
120880=>"111100000",
120881=>"111111101",
120882=>"011111111",
120883=>"111101101",
120884=>"011101011",
120885=>"110111111",
120886=>"101101110",
120887=>"010111000",
120888=>"111000000",
120889=>"000110000",
120890=>"000100100",
120891=>"000000001",
120892=>"110100000",
120893=>"111111000",
120894=>"000000101",
120895=>"111110000",
120896=>"001000010",
120897=>"111111010",
120898=>"110111011",
120899=>"010101000",
120900=>"011001000",
120901=>"000000000",
120902=>"000110110",
120903=>"100000000",
120904=>"111111111",
120905=>"111001011",
120906=>"001000001",
120907=>"111000000",
120908=>"111100100",
120909=>"111101101",
120910=>"011111001",
120911=>"000000000",
120912=>"100101111",
120913=>"110111010",
120914=>"000000000",
120915=>"011001000",
120916=>"111000000",
120917=>"111110101",
120918=>"111100111",
120919=>"011111000",
120920=>"111101001",
120921=>"010000100",
120922=>"011100000",
120923=>"010000111",
120924=>"000000000",
120925=>"011001011",
120926=>"011000001",
120927=>"110001011",
120928=>"000101000",
120929=>"111111011",
120930=>"001000000",
120931=>"110111100",
120932=>"100100000",
120933=>"010011001",
120934=>"110110000",
120935=>"110110110",
120936=>"111000101",
120937=>"111110111",
120938=>"010101100",
120939=>"000110000",
120940=>"111001001",
120941=>"000000100",
120942=>"011011011",
120943=>"000000111",
120944=>"011111111",
120945=>"010000000",
120946=>"011001001",
120947=>"010110000",
120948=>"111000000",
120949=>"000001000",
120950=>"000110111",
120951=>"000001111",
120952=>"000000000",
120953=>"000000000",
120954=>"000010111",
120955=>"000101100",
120956=>"110100110",
120957=>"100100100",
120958=>"111110001",
120959=>"101101101",
120960=>"111000000",
120961=>"111000110",
120962=>"000111011",
120963=>"000000010",
120964=>"110110101",
120965=>"111100001",
120966=>"111011001",
120967=>"001011000",
120968=>"111111111",
120969=>"111001011",
120970=>"010000000",
120971=>"110110000",
120972=>"111111010",
120973=>"011000001",
120974=>"111111111",
120975=>"000000000",
120976=>"111100110",
120977=>"011111000",
120978=>"101110000",
120979=>"111110111",
120980=>"001111111",
120981=>"000000100",
120982=>"110111111",
120983=>"000011000",
120984=>"010010011",
120985=>"000110100",
120986=>"101111111",
120987=>"000000001",
120988=>"000000010",
120989=>"100001101",
120990=>"101101111",
120991=>"000000000",
120992=>"111110110",
120993=>"000000000",
120994=>"111010010",
120995=>"010111101",
120996=>"110010110",
120997=>"110110010",
120998=>"000000111",
120999=>"000111000",
121000=>"110000111",
121001=>"001111101",
121002=>"101001001",
121003=>"000000001",
121004=>"000000010",
121005=>"011010111",
121006=>"010000000",
121007=>"000001110",
121008=>"101111001",
121009=>"111111101",
121010=>"001000100",
121011=>"100100111",
121012=>"000011000",
121013=>"100000101",
121014=>"000000001",
121015=>"000000000",
121016=>"011011000",
121017=>"000111111",
121018=>"000101000",
121019=>"111101111",
121020=>"111010010",
121021=>"111001000",
121022=>"001111111",
121023=>"010111111",
121024=>"000010000",
121025=>"111111010",
121026=>"111111101",
121027=>"110001110",
121028=>"000111000",
121029=>"110110111",
121030=>"111101000",
121031=>"000000000",
121032=>"000111111",
121033=>"000000000",
121034=>"110111101",
121035=>"110001101",
121036=>"010000001",
121037=>"001010111",
121038=>"000000110",
121039=>"000001010",
121040=>"000010000",
121041=>"000101000",
121042=>"001110010",
121043=>"110101000",
121044=>"101000111",
121045=>"110111110",
121046=>"111111010",
121047=>"111000000",
121048=>"000000000",
121049=>"000001101",
121050=>"000110011",
121051=>"111100110",
121052=>"010000100",
121053=>"101010110",
121054=>"000001111",
121055=>"100110100",
121056=>"111010010",
121057=>"001000100",
121058=>"111110000",
121059=>"011101000",
121060=>"000000100",
121061=>"010111111",
121062=>"000000001",
121063=>"100100011",
121064=>"110001000",
121065=>"100010110",
121066=>"111101010",
121067=>"000000000",
121068=>"111111011",
121069=>"110111111",
121070=>"001000000",
121071=>"111001010",
121072=>"111111010",
121073=>"100010010",
121074=>"000000111",
121075=>"000100110",
121076=>"100101010",
121077=>"111000111",
121078=>"000000001",
121079=>"000000100",
121080=>"001000010",
121081=>"111111000",
121082=>"111001000",
121083=>"100110111",
121084=>"000000011",
121085=>"000000000",
121086=>"011111011",
121087=>"010101001",
121088=>"101111100",
121089=>"000000111",
121090=>"000100000",
121091=>"001001011",
121092=>"101110110",
121093=>"101011001",
121094=>"111111111",
121095=>"000000011",
121096=>"100110000",
121097=>"001000011",
121098=>"000000100",
121099=>"000000000",
121100=>"101111111",
121101=>"000001000",
121102=>"100100000",
121103=>"111011101",
121104=>"001000010",
121105=>"000000110",
121106=>"000000110",
121107=>"000000111",
121108=>"111111101",
121109=>"010110111",
121110=>"011111000",
121111=>"010000000",
121112=>"101000111",
121113=>"111101101",
121114=>"101001111",
121115=>"011000000",
121116=>"110001111",
121117=>"111110111",
121118=>"100100011",
121119=>"110001101",
121120=>"100000000",
121121=>"001001111",
121122=>"000111111",
121123=>"111111110",
121124=>"110000110",
121125=>"001111011",
121126=>"001000111",
121127=>"111000000",
121128=>"110111101",
121129=>"001111111",
121130=>"000101000",
121131=>"111001000",
121132=>"100110111",
121133=>"101000110",
121134=>"000000111",
121135=>"110111101",
121136=>"000100001",
121137=>"111100010",
121138=>"000111011",
121139=>"100011001",
121140=>"000100000",
121141=>"110000010",
121142=>"100110100",
121143=>"100111111",
121144=>"101001101",
121145=>"100000000",
121146=>"101001000",
121147=>"111111100",
121148=>"110100111",
121149=>"010111010",
121150=>"000000011",
121151=>"001100110",
121152=>"111100010",
121153=>"001100111",
121154=>"000100111",
121155=>"100000000",
121156=>"000001001",
121157=>"000101000",
121158=>"111110000",
121159=>"101000000",
121160=>"011100111",
121161=>"000000010",
121162=>"000000000",
121163=>"000001111",
121164=>"000000100",
121165=>"000100011",
121166=>"110111110",
121167=>"000000011",
121168=>"000011111",
121169=>"111010000",
121170=>"101100000",
121171=>"000010000",
121172=>"000001000",
121173=>"011011111",
121174=>"011110110",
121175=>"001000000",
121176=>"000110111",
121177=>"001011010",
121178=>"000001011",
121179=>"000000011",
121180=>"100101101",
121181=>"001100000",
121182=>"111111000",
121183=>"001000100",
121184=>"000101101",
121185=>"000000111",
121186=>"000000101",
121187=>"000110110",
121188=>"100001001",
121189=>"010101101",
121190=>"101111010",
121191=>"011111111",
121192=>"000000001",
121193=>"101000000",
121194=>"111000000",
121195=>"000000001",
121196=>"100101101",
121197=>"000000100",
121198=>"100000000",
121199=>"011011111",
121200=>"100001101",
121201=>"001101101",
121202=>"000001001",
121203=>"001000100",
121204=>"100110111",
121205=>"000000001",
121206=>"000100111",
121207=>"011111010",
121208=>"010101100",
121209=>"101111010",
121210=>"000100111",
121211=>"111010010",
121212=>"100001101",
121213=>"001001010",
121214=>"011010010",
121215=>"000000000",
121216=>"101000100",
121217=>"000000011",
121218=>"110110000",
121219=>"111010110",
121220=>"010010010",
121221=>"110000111",
121222=>"000001100",
121223=>"001100101",
121224=>"001001101",
121225=>"111110101",
121226=>"100100100",
121227=>"111100010",
121228=>"111001000",
121229=>"010011111",
121230=>"000000001",
121231=>"000000110",
121232=>"100111011",
121233=>"000000110",
121234=>"100101001",
121235=>"000000010",
121236=>"000000100",
121237=>"100000000",
121238=>"101101000",
121239=>"000110110",
121240=>"101110000",
121241=>"111111011",
121242=>"011100000",
121243=>"010000000",
121244=>"100111111",
121245=>"100000111",
121246=>"100001111",
121247=>"000001111",
121248=>"111100101",
121249=>"000000001",
121250=>"111101000",
121251=>"100101111",
121252=>"111100100",
121253=>"100100111",
121254=>"000111001",
121255=>"110001011",
121256=>"111000000",
121257=>"000001100",
121258=>"100100000",
121259=>"000100111",
121260=>"010010011",
121261=>"000000101",
121262=>"000110110",
121263=>"111111111",
121264=>"111000100",
121265=>"000101110",
121266=>"001011000",
121267=>"000101000",
121268=>"011011111",
121269=>"111011000",
121270=>"011111111",
121271=>"101101101",
121272=>"011000111",
121273=>"010000011",
121274=>"010011001",
121275=>"100101101",
121276=>"101111101",
121277=>"000101111",
121278=>"111001010",
121279=>"000000000",
121280=>"100010110",
121281=>"000000010",
121282=>"000111011",
121283=>"101110110",
121284=>"010100001",
121285=>"110011011",
121286=>"000011000",
121287=>"101100000",
121288=>"111101001",
121289=>"010111000",
121290=>"111111010",
121291=>"000100100",
121292=>"000010001",
121293=>"000000110",
121294=>"000111010",
121295=>"000111100",
121296=>"000010110",
121297=>"111011111",
121298=>"000110111",
121299=>"111011010",
121300=>"010000100",
121301=>"000111100",
121302=>"001001000",
121303=>"111001111",
121304=>"111010000",
121305=>"000110001",
121306=>"101111100",
121307=>"100000111",
121308=>"110011110",
121309=>"001011011",
121310=>"001111110",
121311=>"000111001",
121312=>"010010000",
121313=>"100101011",
121314=>"111011000",
121315=>"001100101",
121316=>"000100000",
121317=>"111111111",
121318=>"111100110",
121319=>"000011011",
121320=>"111101101",
121321=>"111110111",
121322=>"000001001",
121323=>"101111101",
121324=>"010000000",
121325=>"000000000",
121326=>"111001000",
121327=>"111101011",
121328=>"111111110",
121329=>"011110110",
121330=>"000100000",
121331=>"110110000",
121332=>"000010011",
121333=>"101000110",
121334=>"000000111",
121335=>"000010010",
121336=>"001000000",
121337=>"101000010",
121338=>"111111011",
121339=>"010011101",
121340=>"111101000",
121341=>"011011111",
121342=>"111111110",
121343=>"000000010",
121344=>"010111111",
121345=>"110000000",
121346=>"111010000",
121347=>"000000001",
121348=>"010110101",
121349=>"000110000",
121350=>"101110110",
121351=>"000000111",
121352=>"001110101",
121353=>"110100000",
121354=>"001110111",
121355=>"000100110",
121356=>"110000000",
121357=>"000001100",
121358=>"100001011",
121359=>"110000111",
121360=>"110101111",
121361=>"000000111",
121362=>"111111111",
121363=>"000111111",
121364=>"000000000",
121365=>"110111000",
121366=>"000100010",
121367=>"000000111",
121368=>"010000001",
121369=>"111010001",
121370=>"000101111",
121371=>"111110100",
121372=>"001101111",
121373=>"000010010",
121374=>"111001111",
121375=>"101101000",
121376=>"010010000",
121377=>"000000111",
121378=>"000010000",
121379=>"100000000",
121380=>"011000000",
121381=>"000000011",
121382=>"111100000",
121383=>"000011000",
121384=>"011000000",
121385=>"100111111",
121386=>"101000111",
121387=>"011000000",
121388=>"001000111",
121389=>"101010000",
121390=>"000001000",
121391=>"000011010",
121392=>"000111111",
121393=>"101110100",
121394=>"001111111",
121395=>"000100111",
121396=>"011001010",
121397=>"000001111",
121398=>"100001011",
121399=>"010011111",
121400=>"010000001",
121401=>"111101101",
121402=>"000000000",
121403=>"001001110",
121404=>"001001001",
121405=>"011011001",
121406=>"000000000",
121407=>"101100010",
121408=>"101101111",
121409=>"110010010",
121410=>"000110010",
121411=>"011111100",
121412=>"000010000",
121413=>"011111000",
121414=>"111110101",
121415=>"010010011",
121416=>"001001001",
121417=>"111101101",
121418=>"001000000",
121419=>"010101011",
121420=>"011111000",
121421=>"101101000",
121422=>"001011001",
121423=>"011111011",
121424=>"101111000",
121425=>"111111111",
121426=>"000010111",
121427=>"001100100",
121428=>"111101001",
121429=>"000000110",
121430=>"101101110",
121431=>"000000111",
121432=>"110011111",
121433=>"100000100",
121434=>"100100000",
121435=>"011001110",
121436=>"101000000",
121437=>"101101000",
121438=>"111111111",
121439=>"100001011",
121440=>"111111111",
121441=>"111111111",
121442=>"000000000",
121443=>"001101100",
121444=>"111111000",
121445=>"011011111",
121446=>"110010111",
121447=>"111111000",
121448=>"100000011",
121449=>"010000111",
121450=>"001001111",
121451=>"100111000",
121452=>"000000000",
121453=>"001100111",
121454=>"000000000",
121455=>"000000111",
121456=>"110111010",
121457=>"000000111",
121458=>"010000110",
121459=>"010010011",
121460=>"000000011",
121461=>"001000000",
121462=>"111000111",
121463=>"100000000",
121464=>"000000100",
121465=>"001001000",
121466=>"000111111",
121467=>"000000000",
121468=>"001001111",
121469=>"101011000",
121470=>"011111010",
121471=>"111101000",
121472=>"100000111",
121473=>"011111111",
121474=>"001000000",
121475=>"001001000",
121476=>"000000111",
121477=>"111110010",
121478=>"000000110",
121479=>"110001001",
121480=>"110111011",
121481=>"000000111",
121482=>"101111011",
121483=>"111010000",
121484=>"110010000",
121485=>"111011101",
121486=>"111011000",
121487=>"111000001",
121488=>"001111110",
121489=>"001111111",
121490=>"111000001",
121491=>"111111111",
121492=>"000001101",
121493=>"000000111",
121494=>"110111000",
121495=>"001001011",
121496=>"000100111",
121497=>"100010000",
121498=>"001011101",
121499=>"001100001",
121500=>"111110111",
121501=>"111111111",
121502=>"000100111",
121503=>"010110101",
121504=>"001111100",
121505=>"110011111",
121506=>"111111010",
121507=>"111011000",
121508=>"110001111",
121509=>"111010001",
121510=>"100110101",
121511=>"001000010",
121512=>"000000111",
121513=>"010000000",
121514=>"110000000",
121515=>"000111111",
121516=>"000000000",
121517=>"101101111",
121518=>"101101000",
121519=>"110110000",
121520=>"111111100",
121521=>"001101100",
121522=>"001000000",
121523=>"011100100",
121524=>"111011010",
121525=>"000000111",
121526=>"011011000",
121527=>"101101001",
121528=>"000100000",
121529=>"011101100",
121530=>"101010010",
121531=>"110111101",
121532=>"111111000",
121533=>"011010111",
121534=>"100011111",
121535=>"000000000",
121536=>"100111000",
121537=>"100111000",
121538=>"000000011",
121539=>"100011011",
121540=>"000111000",
121541=>"100000001",
121542=>"000010111",
121543=>"110000000",
121544=>"111111000",
121545=>"011010000",
121546=>"010010000",
121547=>"000001111",
121548=>"000110100",
121549=>"000001001",
121550=>"010001000",
121551=>"011011001",
121552=>"111001010",
121553=>"110100000",
121554=>"111010000",
121555=>"011010111",
121556=>"111111000",
121557=>"011001000",
121558=>"111111000",
121559=>"000000001",
121560=>"111110000",
121561=>"001001111",
121562=>"110010000",
121563=>"000000100",
121564=>"000011111",
121565=>"111000101",
121566=>"111010101",
121567=>"101111111",
121568=>"110110000",
121569=>"000001111",
121570=>"111111011",
121571=>"111011000",
121572=>"111001000",
121573=>"011000000",
121574=>"111000111",
121575=>"011011001",
121576=>"000101111",
121577=>"111000000",
121578=>"111101111",
121579=>"010110111",
121580=>"000110111",
121581=>"010101011",
121582=>"001000000",
121583=>"101101111",
121584=>"001001111",
121585=>"001010000",
121586=>"000000000",
121587=>"001000000",
121588=>"110010011",
121589=>"101011000",
121590=>"011000000",
121591=>"011111011",
121592=>"000000111",
121593=>"101001111",
121594=>"111100000",
121595=>"110001000",
121596=>"000110111",
121597=>"000011000",
121598=>"101111111",
121599=>"000000101",
121600=>"000010000",
121601=>"000000110",
121602=>"101111111",
121603=>"110000000",
121604=>"000011001",
121605=>"110110000",
121606=>"111001111",
121607=>"111010110",
121608=>"000000110",
121609=>"111000000",
121610=>"010000000",
121611=>"110110010",
121612=>"000111111",
121613=>"001001001",
121614=>"000000011",
121615=>"000110010",
121616=>"000000100",
121617=>"111111000",
121618=>"001010001",
121619=>"010000011",
121620=>"001001111",
121621=>"011111111",
121622=>"000001011",
121623=>"010001111",
121624=>"111001000",
121625=>"101111000",
121626=>"000111111",
121627=>"010000011",
121628=>"101110111",
121629=>"000101000",
121630=>"000000000",
121631=>"111101101",
121632=>"000110000",
121633=>"100000010",
121634=>"000000010",
121635=>"000110111",
121636=>"001001100",
121637=>"000000000",
121638=>"000110111",
121639=>"001001111",
121640=>"111000010",
121641=>"110010001",
121642=>"111000001",
121643=>"101000000",
121644=>"101111011",
121645=>"011001110",
121646=>"111111101",
121647=>"000001000",
121648=>"111101000",
121649=>"011011000",
121650=>"010010101",
121651=>"100110111",
121652=>"001000000",
121653=>"100110110",
121654=>"000100001",
121655=>"010001101",
121656=>"001000010",
121657=>"111000000",
121658=>"111101101",
121659=>"111000010",
121660=>"011010100",
121661=>"111001010",
121662=>"000111110",
121663=>"010110110",
121664=>"001110111",
121665=>"000100000",
121666=>"111110010",
121667=>"011011000",
121668=>"001000000",
121669=>"001000000",
121670=>"000000001",
121671=>"111111100",
121672=>"111100000",
121673=>"010010010",
121674=>"110000000",
121675=>"101101000",
121676=>"000101001",
121677=>"100001011",
121678=>"010111000",
121679=>"101001111",
121680=>"001000000",
121681=>"011011111",
121682=>"000000000",
121683=>"011000100",
121684=>"000010000",
121685=>"010011111",
121686=>"011011001",
121687=>"111110000",
121688=>"011110101",
121689=>"110110011",
121690=>"001111110",
121691=>"100111110",
121692=>"000001111",
121693=>"001001001",
121694=>"000001111",
121695=>"110100000",
121696=>"010000111",
121697=>"000000000",
121698=>"110000000",
121699=>"100001011",
121700=>"111010000",
121701=>"111000100",
121702=>"101000000",
121703=>"111001001",
121704=>"111111101",
121705=>"000100000",
121706=>"111000000",
121707=>"001001000",
121708=>"111111101",
121709=>"010000001",
121710=>"000101101",
121711=>"110000010",
121712=>"111011111",
121713=>"100000001",
121714=>"000000100",
121715=>"000110010",
121716=>"111000000",
121717=>"111000000",
121718=>"000010010",
121719=>"000100111",
121720=>"011011000",
121721=>"111111000",
121722=>"111111111",
121723=>"000111000",
121724=>"101100001",
121725=>"110100000",
121726=>"000001010",
121727=>"000001101",
121728=>"000110110",
121729=>"110111010",
121730=>"000100111",
121731=>"010000110",
121732=>"001010111",
121733=>"001001101",
121734=>"001000001",
121735=>"000010001",
121736=>"110111100",
121737=>"000101000",
121738=>"000100000",
121739=>"111100000",
121740=>"111101101",
121741=>"000111111",
121742=>"111111111",
121743=>"110000000",
121744=>"001100001",
121745=>"111110111",
121746=>"001000101",
121747=>"111100010",
121748=>"001011110",
121749=>"111010110",
121750=>"001111111",
121751=>"000111110",
121752=>"110101000",
121753=>"000000111",
121754=>"000000110",
121755=>"000000000",
121756=>"111000101",
121757=>"110111000",
121758=>"110011011",
121759=>"111010000",
121760=>"100110111",
121761=>"001000000",
121762=>"110111001",
121763=>"010111001",
121764=>"111110110",
121765=>"000111111",
121766=>"101110101",
121767=>"111111011",
121768=>"111100111",
121769=>"000010010",
121770=>"111110110",
121771=>"111110010",
121772=>"101110110",
121773=>"110111110",
121774=>"111110010",
121775=>"111011111",
121776=>"111110101",
121777=>"011011000",
121778=>"000001000",
121779=>"001001001",
121780=>"010010111",
121781=>"000111111",
121782=>"000000010",
121783=>"000110110",
121784=>"110000110",
121785=>"000100100",
121786=>"000000110",
121787=>"111001010",
121788=>"010000111",
121789=>"111111110",
121790=>"000011011",
121791=>"000000000",
121792=>"000000000",
121793=>"000100000",
121794=>"110010111",
121795=>"001111100",
121796=>"100001101",
121797=>"111001001",
121798=>"110111010",
121799=>"011000000",
121800=>"000010000",
121801=>"000000110",
121802=>"000000110",
121803=>"101000001",
121804=>"111010100",
121805=>"001001100",
121806=>"110111110",
121807=>"010101000",
121808=>"000110110",
121809=>"000110100",
121810=>"111000000",
121811=>"000110111",
121812=>"001011111",
121813=>"100100100",
121814=>"000000101",
121815=>"101001101",
121816=>"101001001",
121817=>"000000110",
121818=>"001111110",
121819=>"111001000",
121820=>"001000000",
121821=>"111110110",
121822=>"000110111",
121823=>"111001001",
121824=>"000010110",
121825=>"000000100",
121826=>"101111111",
121827=>"001111101",
121828=>"100101000",
121829=>"111111000",
121830=>"011111111",
121831=>"111011111",
121832=>"011010010",
121833=>"000000001",
121834=>"010000001",
121835=>"000000111",
121836=>"111111111",
121837=>"110110100",
121838=>"000010000",
121839=>"000100110",
121840=>"000000111",
121841=>"111000101",
121842=>"111000000",
121843=>"000001111",
121844=>"100000011",
121845=>"000000000",
121846=>"110101000",
121847=>"110000000",
121848=>"000000110",
121849=>"011111101",
121850=>"000000010",
121851=>"000000011",
121852=>"100111111",
121853=>"101000000",
121854=>"010111111",
121855=>"111100001",
121856=>"000100100",
121857=>"100000001",
121858=>"000000001",
121859=>"000001000",
121860=>"111111000",
121861=>"111111111",
121862=>"001001111",
121863=>"111010000",
121864=>"010011000",
121865=>"111101001",
121866=>"000010111",
121867=>"000000000",
121868=>"000000111",
121869=>"110111110",
121870=>"011011011",
121871=>"001000000",
121872=>"111110010",
121873=>"001000111",
121874=>"000100100",
121875=>"101001000",
121876=>"011101111",
121877=>"100100000",
121878=>"101000001",
121879=>"001001001",
121880=>"001000111",
121881=>"110111111",
121882=>"110111000",
121883=>"011000000",
121884=>"000010000",
121885=>"000001101",
121886=>"011111111",
121887=>"110000000",
121888=>"001001011",
121889=>"110110110",
121890=>"110100010",
121891=>"110010110",
121892=>"101100000",
121893=>"001011011",
121894=>"010110010",
121895=>"000000000",
121896=>"010111110",
121897=>"000000100",
121898=>"000001101",
121899=>"000000010",
121900=>"101100101",
121901=>"001010111",
121902=>"000101111",
121903=>"101001001",
121904=>"110111110",
121905=>"001100111",
121906=>"001111110",
121907=>"001111110",
121908=>"000000001",
121909=>"001100011",
121910=>"000000001",
121911=>"000000100",
121912=>"011000001",
121913=>"001000001",
121914=>"101101110",
121915=>"000001111",
121916=>"100010100",
121917=>"001111010",
121918=>"000000000",
121919=>"011111000",
121920=>"111111111",
121921=>"101101111",
121922=>"101000111",
121923=>"110111111",
121924=>"000001101",
121925=>"001110110",
121926=>"011011000",
121927=>"101101010",
121928=>"101000110",
121929=>"110010000",
121930=>"001000111",
121931=>"000001110",
121932=>"110000000",
121933=>"111100010",
121934=>"000011001",
121935=>"001000010",
121936=>"100000000",
121937=>"000011111",
121938=>"001000101",
121939=>"101100000",
121940=>"101000111",
121941=>"011110010",
121942=>"011011011",
121943=>"111111000",
121944=>"101101111",
121945=>"101100101",
121946=>"111010000",
121947=>"111001001",
121948=>"000110000",
121949=>"000000011",
121950=>"101011001",
121951=>"011111110",
121952=>"001000000",
121953=>"001111110",
121954=>"000000001",
121955=>"001000000",
121956=>"100110100",
121957=>"111110111",
121958=>"001011110",
121959=>"111101000",
121960=>"111110010",
121961=>"001001011",
121962=>"000101111",
121963=>"110110111",
121964=>"101000011",
121965=>"101111111",
121966=>"100100100",
121967=>"000000111",
121968=>"111100000",
121969=>"000111101",
121970=>"011000100",
121971=>"001001110",
121972=>"001101111",
121973=>"000000011",
121974=>"110110000",
121975=>"111111000",
121976=>"000010111",
121977=>"111010010",
121978=>"000111101",
121979=>"000001010",
121980=>"011011001",
121981=>"101000000",
121982=>"111110000",
121983=>"110110110",
121984=>"001001111",
121985=>"001010011",
121986=>"001010101",
121987=>"000101110",
121988=>"101000111",
121989=>"111101110",
121990=>"010100111",
121991=>"110110110",
121992=>"011011101",
121993=>"001011111",
121994=>"000000111",
121995=>"101001111",
121996=>"010000000",
121997=>"001110111",
121998=>"101000000",
121999=>"000000000",
122000=>"001001111",
122001=>"111110000",
122002=>"110000000",
122003=>"101000110",
122004=>"111010000",
122005=>"111101001",
122006=>"100001111",
122007=>"011011111",
122008=>"111111110",
122009=>"010110010",
122010=>"001111110",
122011=>"101100110",
122012=>"001101100",
122013=>"001000111",
122014=>"000111101",
122015=>"001001111",
122016=>"100100010",
122017=>"000010000",
122018=>"000001111",
122019=>"001101000",
122020=>"000000000",
122021=>"111100100",
122022=>"110110110",
122023=>"000000110",
122024=>"111101111",
122025=>"110110110",
122026=>"010000101",
122027=>"000000001",
122028=>"011111110",
122029=>"110010000",
122030=>"101111011",
122031=>"001000110",
122032=>"110110000",
122033=>"001001011",
122034=>"000100111",
122035=>"000101101",
122036=>"111111111",
122037=>"000000001",
122038=>"000000010",
122039=>"101111101",
122040=>"011010011",
122041=>"011101010",
122042=>"010000110",
122043=>"110110100",
122044=>"001001010",
122045=>"111110000",
122046=>"001000000",
122047=>"000101101",
122048=>"000000001",
122049=>"101001000",
122050=>"010111010",
122051=>"110110001",
122052=>"000101111",
122053=>"001101111",
122054=>"111000000",
122055=>"010010000",
122056=>"110000000",
122057=>"111110010",
122058=>"001001111",
122059=>"001000000",
122060=>"000000000",
122061=>"111000000",
122062=>"101000000",
122063=>"110110000",
122064=>"111011000",
122065=>"110100110",
122066=>"110110000",
122067=>"100000000",
122068=>"111000000",
122069=>"000000111",
122070=>"001100101",
122071=>"111111101",
122072=>"011110111",
122073=>"000000000",
122074=>"011001000",
122075=>"001001101",
122076=>"001001101",
122077=>"011001111",
122078=>"000000110",
122079=>"111101101",
122080=>"010010000",
122081=>"000001101",
122082=>"001001111",
122083=>"100101111",
122084=>"001000000",
122085=>"000001011",
122086=>"111001111",
122087=>"011100100",
122088=>"000101111",
122089=>"000000000",
122090=>"001100111",
122091=>"001001001",
122092=>"110000000",
122093=>"000111000",
122094=>"000000000",
122095=>"100110111",
122096=>"000000111",
122097=>"001101111",
122098=>"101001111",
122099=>"001011100",
122100=>"110101000",
122101=>"111001100",
122102=>"000000000",
122103=>"101011110",
122104=>"010110010",
122105=>"001001010",
122106=>"000000000",
122107=>"111001001",
122108=>"000111111",
122109=>"100101101",
122110=>"110110011",
122111=>"000010110",
122112=>"011011100",
122113=>"001001100",
122114=>"111101101",
122115=>"110010000",
122116=>"100110110",
122117=>"111000010",
122118=>"000010000",
122119=>"100010010",
122120=>"001011100",
122121=>"101100100",
122122=>"000110110",
122123=>"111101111",
122124=>"000000000",
122125=>"010111111",
122126=>"111100010",
122127=>"111011001",
122128=>"011100100",
122129=>"111000000",
122130=>"101100101",
122131=>"000000000",
122132=>"111100000",
122133=>"110000000",
122134=>"111101101",
122135=>"111111101",
122136=>"101000111",
122137=>"001010010",
122138=>"000111101",
122139=>"000001001",
122140=>"111011000",
122141=>"000000000",
122142=>"111101001",
122143=>"011111010",
122144=>"101001000",
122145=>"000111111",
122146=>"100000011",
122147=>"000010011",
122148=>"001001001",
122149=>"110010010",
122150=>"111111000",
122151=>"000010000",
122152=>"111111111",
122153=>"111111100",
122154=>"101111111",
122155=>"101000000",
122156=>"011111011",
122157=>"010010010",
122158=>"110000100",
122159=>"110110111",
122160=>"111001000",
122161=>"101100100",
122162=>"101010010",
122163=>"001010111",
122164=>"000000001",
122165=>"000100000",
122166=>"010110100",
122167=>"000000010",
122168=>"100000011",
122169=>"000011010",
122170=>"000001001",
122171=>"101101000",
122172=>"100110010",
122173=>"000111000",
122174=>"000101100",
122175=>"111111100",
122176=>"111101000",
122177=>"111111000",
122178=>"000011111",
122179=>"011101000",
122180=>"010111011",
122181=>"011000101",
122182=>"000100111",
122183=>"011011010",
122184=>"000000010",
122185=>"000000000",
122186=>"000110100",
122187=>"000010111",
122188=>"111000001",
122189=>"000110100",
122190=>"101101001",
122191=>"110111010",
122192=>"010010011",
122193=>"111101111",
122194=>"010010000",
122195=>"011000000",
122196=>"000110000",
122197=>"101000100",
122198=>"000110100",
122199=>"100100100",
122200=>"000111011",
122201=>"000111000",
122202=>"000001000",
122203=>"000101111",
122204=>"000000000",
122205=>"010101101",
122206=>"111000000",
122207=>"100000001",
122208=>"111111010",
122209=>"000000000",
122210=>"100100101",
122211=>"111110100",
122212=>"100111100",
122213=>"000110100",
122214=>"011010010",
122215=>"111000000",
122216=>"111101111",
122217=>"111111110",
122218=>"101000111",
122219=>"111010100",
122220=>"000001010",
122221=>"111111111",
122222=>"000100000",
122223=>"110110101",
122224=>"110101010",
122225=>"111101000",
122226=>"011101001",
122227=>"100010100",
122228=>"110111001",
122229=>"111100101",
122230=>"000000111",
122231=>"111100000",
122232=>"111000000",
122233=>"000111111",
122234=>"101000011",
122235=>"100100110",
122236=>"100110000",
122237=>"010010000",
122238=>"101100010",
122239=>"111100111",
122240=>"000010000",
122241=>"111100100",
122242=>"110110101",
122243=>"010111111",
122244=>"000010010",
122245=>"111111000",
122246=>"110010001",
122247=>"000100000",
122248=>"001110110",
122249=>"000100010",
122250=>"111111111",
122251=>"111100111",
122252=>"101100101",
122253=>"111000001",
122254=>"000010001",
122255=>"000000000",
122256=>"011111100",
122257=>"000000000",
122258=>"101101100",
122259=>"000000000",
122260=>"000101110",
122261=>"101100101",
122262=>"010111000",
122263=>"100100100",
122264=>"100010010",
122265=>"111111011",
122266=>"111111000",
122267=>"111000100",
122268=>"000010011",
122269=>"100101000",
122270=>"011011010",
122271=>"010111101",
122272=>"100101001",
122273=>"101100101",
122274=>"111111000",
122275=>"000000011",
122276=>"001101000",
122277=>"000111001",
122278=>"111000001",
122279=>"000010010",
122280=>"011000000",
122281=>"000101110",
122282=>"111110111",
122283=>"000111101",
122284=>"010101111",
122285=>"000000011",
122286=>"000110100",
122287=>"000000110",
122288=>"011000010",
122289=>"000001000",
122290=>"111101101",
122291=>"001001010",
122292=>"111011000",
122293=>"001010000",
122294=>"000100111",
122295=>"000001000",
122296=>"000010010",
122297=>"000000010",
122298=>"010111111",
122299=>"000010010",
122300=>"110111111",
122301=>"111101111",
122302=>"111001001",
122303=>"101101010",
122304=>"000000000",
122305=>"000000111",
122306=>"111111100",
122307=>"110001001",
122308=>"001111011",
122309=>"011001111",
122310=>"000011011",
122311=>"101100111",
122312=>"101010100",
122313=>"111101100",
122314=>"111001111",
122315=>"101000000",
122316=>"111100000",
122317=>"001001010",
122318=>"100000000",
122319=>"111111111",
122320=>"010000000",
122321=>"000011001",
122322=>"000010111",
122323=>"111111000",
122324=>"100100001",
122325=>"100000010",
122326=>"010111110",
122327=>"010111010",
122328=>"111001000",
122329=>"100010011",
122330=>"011011010",
122331=>"101100111",
122332=>"111111001",
122333=>"100011000",
122334=>"000111111",
122335=>"000000000",
122336=>"101000101",
122337=>"011000000",
122338=>"111000001",
122339=>"001001111",
122340=>"101000000",
122341=>"111000010",
122342=>"101111101",
122343=>"000010101",
122344=>"000000000",
122345=>"000010000",
122346=>"100001101",
122347=>"000000111",
122348=>"111000000",
122349=>"111000001",
122350=>"000000000",
122351=>"000110100",
122352=>"000000000",
122353=>"010100111",
122354=>"111101000",
122355=>"000011001",
122356=>"000010001",
122357=>"000000111",
122358=>"000000010",
122359=>"000000011",
122360=>"111001000",
122361=>"000010011",
122362=>"010001111",
122363=>"000111010",
122364=>"011111111",
122365=>"111100000",
122366=>"010011011",
122367=>"111111111",
122368=>"001111111",
122369=>"001000100",
122370=>"001010000",
122371=>"111011001",
122372=>"000100111",
122373=>"000001000",
122374=>"101000000",
122375=>"111011111",
122376=>"111001001",
122377=>"001010110",
122378=>"000110110",
122379=>"000000000",
122380=>"001101101",
122381=>"111000000",
122382=>"011111010",
122383=>"100110010",
122384=>"111001000",
122385=>"111000000",
122386=>"110001000",
122387=>"110110000",
122388=>"011111111",
122389=>"111111001",
122390=>"001011001",
122391=>"111000101",
122392=>"001000000",
122393=>"111001001",
122394=>"001000000",
122395=>"000110110",
122396=>"000001000",
122397=>"000111110",
122398=>"010110001",
122399=>"111001000",
122400=>"001010000",
122401=>"011000001",
122402=>"000000110",
122403=>"000000100",
122404=>"100100001",
122405=>"110100100",
122406=>"011111000",
122407=>"000000000",
122408=>"000110110",
122409=>"000000110",
122410=>"001001001",
122411=>"010111010",
122412=>"010111111",
122413=>"001111010",
122414=>"011111111",
122415=>"101000000",
122416=>"000000110",
122417=>"000101101",
122418=>"100000111",
122419=>"110110111",
122420=>"001110110",
122421=>"100110111",
122422=>"010111001",
122423=>"111001001",
122424=>"110000001",
122425=>"111001001",
122426=>"101001000",
122427=>"111110110",
122428=>"101111110",
122429=>"011011111",
122430=>"001000000",
122431=>"000101100",
122432=>"110101000",
122433=>"100100111",
122434=>"111001000",
122435=>"111001000",
122436=>"001001000",
122437=>"001000000",
122438=>"000000101",
122439=>"000000100",
122440=>"001001000",
122441=>"111000000",
122442=>"111001001",
122443=>"111001001",
122444=>"111011000",
122445=>"001100100",
122446=>"001111111",
122447=>"110110110",
122448=>"111100000",
122449=>"110111111",
122450=>"111101110",
122451=>"010000000",
122452=>"110000000",
122453=>"001110110",
122454=>"001011001",
122455=>"011000000",
122456=>"111001000",
122457=>"011100100",
122458=>"011111111",
122459=>"111111010",
122460=>"001001001",
122461=>"000000000",
122462=>"000110100",
122463=>"101000001",
122464=>"001011000",
122465=>"110001000",
122466=>"000001111",
122467=>"101101100",
122468=>"111111001",
122469=>"011000000",
122470=>"000001001",
122471=>"000110110",
122472=>"111010100",
122473=>"110010000",
122474=>"000000110",
122475=>"001001000",
122476=>"000010110",
122477=>"110110110",
122478=>"111011011",
122479=>"000000000",
122480=>"000110110",
122481=>"001000111",
122482=>"110011000",
122483=>"010110010",
122484=>"000000000",
122485=>"011001000",
122486=>"011001000",
122487=>"001110000",
122488=>"010000000",
122489=>"111110100",
122490=>"000110110",
122491=>"000000000",
122492=>"011011110",
122493=>"111100000",
122494=>"011000001",
122495=>"111100000",
122496=>"100000000",
122497=>"111001000",
122498=>"000110110",
122499=>"000000111",
122500=>"110111001",
122501=>"000110111",
122502=>"001111110",
122503=>"111101100",
122504=>"011011011",
122505=>"000110110",
122506=>"111110000",
122507=>"000101100",
122508=>"111101110",
122509=>"100110110",
122510=>"001110110",
122511=>"110101000",
122512=>"111001000",
122513=>"101101100",
122514=>"001000000",
122515=>"100111101",
122516=>"110110110",
122517=>"110000000",
122518=>"101111100",
122519=>"000001111",
122520=>"000110110",
122521=>"100001101",
122522=>"000110111",
122523=>"000000000",
122524=>"111111001",
122525=>"000110110",
122526=>"111111111",
122527=>"111001001",
122528=>"001000001",
122529=>"000000001",
122530=>"001001000",
122531=>"111000001",
122532=>"000001010",
122533=>"011010000",
122534=>"001110111",
122535=>"000110110",
122536=>"000010110",
122537=>"000101001",
122538=>"000000000",
122539=>"111010001",
122540=>"000000000",
122541=>"111101000",
122542=>"100100000",
122543=>"100001000",
122544=>"010001001",
122545=>"111001011",
122546=>"110001000",
122547=>"000001100",
122548=>"001111111",
122549=>"110000000",
122550=>"010000000",
122551=>"000110110",
122552=>"100111110",
122553=>"110111110",
122554=>"000110111",
122555=>"101000111",
122556=>"100111111",
122557=>"000110111",
122558=>"000000000",
122559=>"001000000",
122560=>"111001000",
122561=>"000000001",
122562=>"110111000",
122563=>"001011011",
122564=>"110110111",
122565=>"011101110",
122566=>"111000100",
122567=>"111001000",
122568=>"111001111",
122569=>"111001000",
122570=>"111111110",
122571=>"111001001",
122572=>"111001000",
122573=>"100100110",
122574=>"010000111",
122575=>"110001111",
122576=>"011001000",
122577=>"011101010",
122578=>"111000011",
122579=>"111111010",
122580=>"111001001",
122581=>"010001000",
122582=>"111001000",
122583=>"011000110",
122584=>"111001000",
122585=>"100000000",
122586=>"001000000",
122587=>"100100110",
122588=>"100001000",
122589=>"000110110",
122590=>"101001000",
122591=>"001110111",
122592=>"111001000",
122593=>"111001001",
122594=>"100101111",
122595=>"111001001",
122596=>"111001000",
122597=>"001011111",
122598=>"000011011",
122599=>"110110010",
122600=>"000111000",
122601=>"000010000",
122602=>"000110110",
122603=>"001001101",
122604=>"111001000",
122605=>"110001001",
122606=>"000001001",
122607=>"000110010",
122608=>"000110110",
122609=>"001010010",
122610=>"000000000",
122611=>"010010000",
122612=>"000110111",
122613=>"001001111",
122614=>"110100100",
122615=>"000110110",
122616=>"000001001",
122617=>"110111100",
122618=>"001110110",
122619=>"111111000",
122620=>"000100101",
122621=>"000110011",
122622=>"000111111",
122623=>"111001001",
122624=>"000000000",
122625=>"001011111",
122626=>"000010001",
122627=>"001000100",
122628=>"110111110",
122629=>"110101100",
122630=>"000000000",
122631=>"011111001",
122632=>"111101100",
122633=>"011000011",
122634=>"111110100",
122635=>"100001110",
122636=>"101011111",
122637=>"000000110",
122638=>"110001000",
122639=>"000011000",
122640=>"111011011",
122641=>"001000000",
122642=>"100000000",
122643=>"000000010",
122644=>"110111111",
122645=>"000100110",
122646=>"110010010",
122647=>"111000001",
122648=>"010000000",
122649=>"111111011",
122650=>"100100110",
122651=>"111110100",
122652=>"000100111",
122653=>"000110100",
122654=>"110010001",
122655=>"100101111",
122656=>"000100000",
122657=>"000000100",
122658=>"100001101",
122659=>"111101100",
122660=>"100101100",
122661=>"100001101",
122662=>"111000000",
122663=>"100010110",
122664=>"001000110",
122665=>"100101111",
122666=>"010000000",
122667=>"011011011",
122668=>"100100000",
122669=>"111001001",
122670=>"000001001",
122671=>"110111111",
122672=>"000000000",
122673=>"100100111",
122674=>"000011011",
122675=>"000001011",
122676=>"001111110",
122677=>"010100000",
122678=>"110100101",
122679=>"011010010",
122680=>"100001001",
122681=>"100110000",
122682=>"000000011",
122683=>"000011000",
122684=>"111011011",
122685=>"100100100",
122686=>"010010000",
122687=>"110111111",
122688=>"011011011",
122689=>"100110001",
122690=>"001101101",
122691=>"001010110",
122692=>"000010000",
122693=>"000010010",
122694=>"000111111",
122695=>"010111000",
122696=>"100111111",
122697=>"100100100",
122698=>"011110100",
122699=>"011011111",
122700=>"110110011",
122701=>"110011011",
122702=>"000000000",
122703=>"101111111",
122704=>"100100110",
122705=>"100000000",
122706=>"101001011",
122707=>"000010110",
122708=>"110000000",
122709=>"000110111",
122710=>"100111111",
122711=>"100000000",
122712=>"000001000",
122713=>"100110111",
122714=>"100001111",
122715=>"001001001",
122716=>"001010011",
122717=>"000001001",
122718=>"111010011",
122719=>"110100100",
122720=>"110100100",
122721=>"101110110",
122722=>"110111000",
122723=>"000001001",
122724=>"000000100",
122725=>"101001101",
122726=>"000101111",
122727=>"000011011",
122728=>"011110100",
122729=>"100000001",
122730=>"101001000",
122731=>"011111011",
122732=>"111000110",
122733=>"111000101",
122734=>"010001001",
122735=>"111000000",
122736=>"100110101",
122737=>"111111001",
122738=>"001011110",
122739=>"100110101",
122740=>"110011110",
122741=>"000101111",
122742=>"000000000",
122743=>"101001011",
122744=>"011000001",
122745=>"100000000",
122746=>"000010010",
122747=>"000011010",
122748=>"111011011",
122749=>"100100000",
122750=>"011011011",
122751=>"110110100",
122752=>"111000000",
122753=>"111000000",
122754=>"011000000",
122755=>"101100000",
122756=>"100100011",
122757=>"100100110",
122758=>"000010100",
122759=>"000000000",
122760=>"100110100",
122761=>"000100100",
122762=>"011001101",
122763=>"011011000",
122764=>"111101011",
122765=>"010001101",
122766=>"111111100",
122767=>"001000100",
122768=>"100110101",
122769=>"100011011",
122770=>"010001111",
122771=>"001001001",
122772=>"000000110",
122773=>"111000011",
122774=>"110000001",
122775=>"101101111",
122776=>"111100100",
122777=>"111011001",
122778=>"000000011",
122779=>"011000110",
122780=>"101100000",
122781=>"010010011",
122782=>"000000001",
122783=>"101001011",
122784=>"000001101",
122785=>"000111011",
122786=>"000001101",
122787=>"101110011",
122788=>"010000000",
122789=>"111111011",
122790=>"111100000",
122791=>"110111110",
122792=>"011111111",
122793=>"011000100",
122794=>"000100100",
122795=>"011000110",
122796=>"000110100",
122797=>"100100111",
122798=>"110110110",
122799=>"001010111",
122800=>"001001100",
122801=>"000011111",
122802=>"001011000",
122803=>"000001101",
122804=>"000100100",
122805=>"001001001",
122806=>"000111110",
122807=>"000111110",
122808=>"100100110",
122809=>"111001111",
122810=>"101011011",
122811=>"100011011",
122812=>"110110111",
122813=>"101100100",
122814=>"000000100",
122815=>"111010110",
122816=>"101011011",
122817=>"111011011",
122818=>"011110100",
122819=>"000110110",
122820=>"011011110",
122821=>"110110000",
122822=>"111000000",
122823=>"011011011",
122824=>"110111011",
122825=>"100100100",
122826=>"001111011",
122827=>"001000011",
122828=>"010110100",
122829=>"010110000",
122830=>"000001011",
122831=>"111011001",
122832=>"100100000",
122833=>"000001000",
122834=>"001101001",
122835=>"010010100",
122836=>"011011111",
122837=>"100100101",
122838=>"111100101",
122839=>"111000011",
122840=>"011111001",
122841=>"011110110",
122842=>"000111111",
122843=>"000000111",
122844=>"100011000",
122845=>"010100100",
122846=>"111100110",
122847=>"111001111",
122848=>"001100100",
122849=>"101011111",
122850=>"001011011",
122851=>"100101110",
122852=>"000100111",
122853=>"110100100",
122854=>"110100100",
122855=>"001001001",
122856=>"101101110",
122857=>"011011111",
122858=>"110010010",
122859=>"100111000",
122860=>"001000000",
122861=>"100111110",
122862=>"000000000",
122863=>"100100100",
122864=>"011000111",
122865=>"000001110",
122866=>"111000010",
122867=>"001011001",
122868=>"110100001",
122869=>"000101000",
122870=>"000011001",
122871=>"011010010",
122872=>"011011011",
122873=>"110100100",
122874=>"110011011",
122875=>"011010011",
122876=>"110111100",
122877=>"011011011",
122878=>"100011100",
122879=>"000001000",
122880=>"100100111",
122881=>"110011111",
122882=>"110000100",
122883=>"011011011",
122884=>"101011011",
122885=>"001100111",
122886=>"110000100",
122887=>"000111011",
122888=>"100101001",
122889=>"000000000",
122890=>"100110111",
122891=>"111101101",
122892=>"111100100",
122893=>"110100111",
122894=>"110111111",
122895=>"011111111",
122896=>"100100110",
122897=>"010011111",
122898=>"101011111",
122899=>"011011001",
122900=>"001111101",
122901=>"101000100",
122902=>"000010001",
122903=>"101111111",
122904=>"101011111",
122905=>"111100000",
122906=>"101111111",
122907=>"111111101",
122908=>"100000000",
122909=>"011111011",
122910=>"000000111",
122911=>"101100100",
122912=>"010100101",
122913=>"111111111",
122914=>"011011001",
122915=>"111000000",
122916=>"110111111",
122917=>"000000011",
122918=>"100011010",
122919=>"111111101",
122920=>"001000000",
122921=>"000111001",
122922=>"100000000",
122923=>"000000000",
122924=>"111111111",
122925=>"111111101",
122926=>"000000010",
122927=>"010110110",
122928=>"111110011",
122929=>"111110111",
122930=>"111011100",
122931=>"010111001",
122932=>"111111011",
122933=>"011011100",
122934=>"100110100",
122935=>"001011011",
122936=>"000111100",
122937=>"000001111",
122938=>"000101101",
122939=>"110010001",
122940=>"111000000",
122941=>"111011111",
122942=>"000000100",
122943=>"010011111",
122944=>"001011000",
122945=>"000000100",
122946=>"011110111",
122947=>"110100111",
122948=>"000000000",
122949=>"001111000",
122950=>"000000000",
122951=>"000000000",
122952=>"110011101",
122953=>"010001000",
122954=>"010010010",
122955=>"000000111",
122956=>"010111111",
122957=>"001111111",
122958=>"100111111",
122959=>"101000101",
122960=>"000000111",
122961=>"111111100",
122962=>"001100101",
122963=>"000110110",
122964=>"000000111",
122965=>"011111001",
122966=>"000110111",
122967=>"111000000",
122968=>"100000000",
122969=>"011011001",
122970=>"000000111",
122971=>"110010110",
122972=>"000111111",
122973=>"000110100",
122974=>"000111010",
122975=>"111000001",
122976=>"000000001",
122977=>"111000000",
122978=>"111000000",
122979=>"001110100",
122980=>"000001000",
122981=>"000000000",
122982=>"101111101",
122983=>"001000000",
122984=>"010010101",
122985=>"000111011",
122986=>"010010010",
122987=>"101100101",
122988=>"000010111",
122989=>"010011011",
122990=>"100100101",
122991=>"101010111",
122992=>"011101101",
122993=>"010000000",
122994=>"100111101",
122995=>"010010000",
122996=>"010010010",
122997=>"110101101",
122998=>"001001000",
122999=>"111001000",
123000=>"000000110",
123001=>"000101001",
123002=>"010000000",
123003=>"111110100",
123004=>"011011011",
123005=>"000001011",
123006=>"001001101",
123007=>"100100101",
123008=>"110100110",
123009=>"000000000",
123010=>"010011111",
123011=>"111111011",
123012=>"101110111",
123013=>"000101000",
123014=>"000000100",
123015=>"111100100",
123016=>"100100000",
123017=>"111111101",
123018=>"000011111",
123019=>"001001011",
123020=>"110000000",
123021=>"000100101",
123022=>"001000000",
123023=>"001000000",
123024=>"010011011",
123025=>"000111111",
123026=>"000111100",
123027=>"110001000",
123028=>"001001111",
123029=>"111001000",
123030=>"000010110",
123031=>"111110100",
123032=>"000101000",
123033=>"011001000",
123034=>"100000000",
123035=>"000100100",
123036=>"110100100",
123037=>"111100000",
123038=>"000100110",
123039=>"100100100",
123040=>"000001111",
123041=>"111111111",
123042=>"000000001",
123043=>"110000111",
123044=>"111111010",
123045=>"100110100",
123046=>"101001000",
123047=>"100000101",
123048=>"000011010",
123049=>"001111001",
123050=>"110101101",
123051=>"101101111",
123052=>"001011111",
123053=>"000111010",
123054=>"010000100",
123055=>"101100101",
123056=>"111100000",
123057=>"100110100",
123058=>"111010000",
123059=>"011000000",
123060=>"101111111",
123061=>"011010011",
123062=>"000001001",
123063=>"101000000",
123064=>"110100100",
123065=>"110011111",
123066=>"010111011",
123067=>"110110100",
123068=>"111101000",
123069=>"101000000",
123070=>"100100100",
123071=>"111010110",
123072=>"000000011",
123073=>"000011000",
123074=>"000100101",
123075=>"001100110",
123076=>"011010001",
123077=>"111111101",
123078=>"000011011",
123079=>"111000110",
123080=>"111101101",
123081=>"000000000",
123082=>"110110100",
123083=>"000100000",
123084=>"100000100",
123085=>"111110100",
123086=>"100011011",
123087=>"110111010",
123088=>"111111111",
123089=>"000111111",
123090=>"111110000",
123091=>"011000111",
123092=>"011101101",
123093=>"000111111",
123094=>"000010101",
123095=>"000000111",
123096=>"000000000",
123097=>"111000000",
123098=>"011100000",
123099=>"000000011",
123100=>"000111110",
123101=>"000101000",
123102=>"000000000",
123103=>"010111111",
123104=>"111100100",
123105=>"011100110",
123106=>"111000100",
123107=>"011011111",
123108=>"100000000",
123109=>"010010011",
123110=>"111100000",
123111=>"001000010",
123112=>"111100100",
123113=>"000000000",
123114=>"100111111",
123115=>"100010111",
123116=>"111000000",
123117=>"000000111",
123118=>"001000011",
123119=>"000000000",
123120=>"100100101",
123121=>"000011100",
123122=>"001000101",
123123=>"110111110",
123124=>"011010011",
123125=>"101111011",
123126=>"000000111",
123127=>"111000000",
123128=>"111000000",
123129=>"010100111",
123130=>"110100111",
123131=>"000101010",
123132=>"111011110",
123133=>"000000000",
123134=>"000111110",
123135=>"011000000",
123136=>"001000000",
123137=>"000000101",
123138=>"001110000",
123139=>"111110000",
123140=>"000001011",
123141=>"000000000",
123142=>"111101011",
123143=>"101001000",
123144=>"111001011",
123145=>"101001001",
123146=>"011011110",
123147=>"000001101",
123148=>"111001111",
123149=>"111111011",
123150=>"001000011",
123151=>"111111110",
123152=>"001001000",
123153=>"000000000",
123154=>"000000000",
123155=>"010001011",
123156=>"001000000",
123157=>"001100100",
123158=>"000100111",
123159=>"100111111",
123160=>"100000011",
123161=>"111110000",
123162=>"001000000",
123163=>"000000000",
123164=>"000101101",
123165=>"101111111",
123166=>"010000011",
123167=>"111111000",
123168=>"101111010",
123169=>"000000011",
123170=>"000011111",
123171=>"110111111",
123172=>"100100111",
123173=>"011000000",
123174=>"000111010",
123175=>"010101001",
123176=>"010010000",
123177=>"010000001",
123178=>"010000001",
123179=>"100000101",
123180=>"010000110",
123181=>"000111111",
123182=>"000111111",
123183=>"000000011",
123184=>"010010011",
123185=>"001011100",
123186=>"000010101",
123187=>"110010000",
123188=>"000000000",
123189=>"110110100",
123190=>"001001011",
123191=>"010101111",
123192=>"010000010",
123193=>"000000000",
123194=>"000000101",
123195=>"000111111",
123196=>"110000100",
123197=>"111101000",
123198=>"100000000",
123199=>"011001001",
123200=>"011000000",
123201=>"000000000",
123202=>"111111111",
123203=>"110001000",
123204=>"000010010",
123205=>"010000000",
123206=>"111111111",
123207=>"110000000",
123208=>"000001100",
123209=>"010010000",
123210=>"000001000",
123211=>"010001001",
123212=>"010011010",
123213=>"111111101",
123214=>"110100000",
123215=>"000000011",
123216=>"000001111",
123217=>"110111000",
123218=>"000001000",
123219=>"000100111",
123220=>"010110111",
123221=>"010001010",
123222=>"011011111",
123223=>"111110010",
123224=>"111110111",
123225=>"001101001",
123226=>"110000011",
123227=>"001000000",
123228=>"111010000",
123229=>"001001001",
123230=>"111111010",
123231=>"110100000",
123232=>"010011000",
123233=>"110010000",
123234=>"000000000",
123235=>"111111101",
123236=>"100000101",
123237=>"100100101",
123238=>"110111001",
123239=>"111001010",
123240=>"110111110",
123241=>"000000000",
123242=>"110101101",
123243=>"000101000",
123244=>"000000010",
123245=>"000010111",
123246=>"110011000",
123247=>"010000010",
123248=>"111111110",
123249=>"000000000",
123250=>"100100100",
123251=>"111111010",
123252=>"000011111",
123253=>"000000000",
123254=>"110110010",
123255=>"111000000",
123256=>"000110010",
123257=>"000000111",
123258=>"000111111",
123259=>"000000111",
123260=>"110110100",
123261=>"100001011",
123262=>"000111111",
123263=>"100111100",
123264=>"001100100",
123265=>"111000000",
123266=>"010000100",
123267=>"111100101",
123268=>"000000000",
123269=>"111111111",
123270=>"000000000",
123271=>"111011010",
123272=>"101001011",
123273=>"000010111",
123274=>"000000001",
123275=>"010000000",
123276=>"111111000",
123277=>"000100000",
123278=>"000000111",
123279=>"001000000",
123280=>"011111111",
123281=>"010110000",
123282=>"010111011",
123283=>"101001011",
123284=>"111111111",
123285=>"011011111",
123286=>"011011000",
123287=>"000000100",
123288=>"110000000",
123289=>"010010010",
123290=>"011111000",
123291=>"001101111",
123292=>"010111111",
123293=>"010000000",
123294=>"100010111",
123295=>"000100101",
123296=>"100100001",
123297=>"000000011",
123298=>"111111001",
123299=>"000000101",
123300=>"000000001",
123301=>"011100100",
123302=>"110110101",
123303=>"010010111",
123304=>"110110111",
123305=>"010101111",
123306=>"000000001",
123307=>"010000000",
123308=>"111000000",
123309=>"111111000",
123310=>"000011001",
123311=>"111111110",
123312=>"101000000",
123313=>"001001111",
123314=>"101110000",
123315=>"000000100",
123316=>"101100111",
123317=>"111111111",
123318=>"111110000",
123319=>"111111100",
123320=>"011001001",
123321=>"110110111",
123322=>"101111100",
123323=>"011111111",
123324=>"111000000",
123325=>"111111011",
123326=>"100100110",
123327=>"000000000",
123328=>"010111000",
123329=>"010010000",
123330=>"110101111",
123331=>"001101100",
123332=>"000010111",
123333=>"000001110",
123334=>"111100000",
123335=>"110100000",
123336=>"111111010",
123337=>"111111011",
123338=>"001000010",
123339=>"111110111",
123340=>"010010010",
123341=>"011011001",
123342=>"000111010",
123343=>"011101110",
123344=>"011111000",
123345=>"000001011",
123346=>"110010010",
123347=>"010101011",
123348=>"010000000",
123349=>"000000111",
123350=>"111110111",
123351=>"000001111",
123352=>"001011010",
123353=>"110101110",
123354=>"000001000",
123355=>"011010011",
123356=>"011011000",
123357=>"010000111",
123358=>"011110010",
123359=>"111000010",
123360=>"000000000",
123361=>"000001101",
123362=>"111110010",
123363=>"000001101",
123364=>"010111000",
123365=>"000000111",
123366=>"100111111",
123367=>"001101101",
123368=>"110100000",
123369=>"110010000",
123370=>"100100111",
123371=>"111111100",
123372=>"001000100",
123373=>"111111110",
123374=>"000000000",
123375=>"001000010",
123376=>"100011010",
123377=>"101110010",
123378=>"000000000",
123379=>"001001111",
123380=>"100100110",
123381=>"000000111",
123382=>"110001000",
123383=>"001111011",
123384=>"010110111",
123385=>"001011111",
123386=>"000100000",
123387=>"111011000",
123388=>"001111111",
123389=>"000000000",
123390=>"100100111",
123391=>"100000101",
123392=>"111101111",
123393=>"000000111",
123394=>"000000110",
123395=>"111111000",
123396=>"101000001",
123397=>"110000000",
123398=>"010111000",
123399=>"000111111",
123400=>"010000000",
123401=>"010010110",
123402=>"001011011",
123403=>"000001110",
123404=>"000000000",
123405=>"011001001",
123406=>"000010011",
123407=>"100000111",
123408=>"111111000",
123409=>"111110010",
123410=>"100100111",
123411=>"101000100",
123412=>"010011111",
123413=>"000110110",
123414=>"100101101",
123415=>"101000000",
123416=>"001000000",
123417=>"111101101",
123418=>"101000000",
123419=>"010000000",
123420=>"100100101",
123421=>"011111101",
123422=>"111111010",
123423=>"110111001",
123424=>"001000001",
123425=>"001001001",
123426=>"000000100",
123427=>"000110111",
123428=>"001000000",
123429=>"100000010",
123430=>"000010110",
123431=>"100000000",
123432=>"011111101",
123433=>"100001001",
123434=>"000111011",
123435=>"110000000",
123436=>"111000000",
123437=>"111111101",
123438=>"000010000",
123439=>"110111111",
123440=>"011110000",
123441=>"101000100",
123442=>"101000111",
123443=>"000100111",
123444=>"000000111",
123445=>"101000101",
123446=>"000111111",
123447=>"111111111",
123448=>"001101000",
123449=>"111111111",
123450=>"000000000",
123451=>"000000000",
123452=>"100001000",
123453=>"111111111",
123454=>"000000000",
123455=>"110110100",
123456=>"000000000",
123457=>"110000010",
123458=>"011011111",
123459=>"011011011",
123460=>"011000001",
123461=>"111001101",
123462=>"100110111",
123463=>"100111111",
123464=>"111101111",
123465=>"010111000",
123466=>"101011111",
123467=>"000000001",
123468=>"101000010",
123469=>"100100000",
123470=>"011000001",
123471=>"000101000",
123472=>"010110110",
123473=>"111111101",
123474=>"000000110",
123475=>"011001100",
123476=>"000000000",
123477=>"110100000",
123478=>"111011001",
123479=>"000111110",
123480=>"001000000",
123481=>"000100100",
123482=>"001001001",
123483=>"011001000",
123484=>"000110000",
123485=>"111001001",
123486=>"010010111",
123487=>"110110111",
123488=>"101100100",
123489=>"000000000",
123490=>"111000000",
123491=>"100100000",
123492=>"100110100",
123493=>"111000110",
123494=>"111101111",
123495=>"110111010",
123496=>"000011111",
123497=>"101111111",
123498=>"011001100",
123499=>"010100111",
123500=>"101111110",
123501=>"000111000",
123502=>"000110110",
123503=>"011001000",
123504=>"100101001",
123505=>"000001000",
123506=>"000100100",
123507=>"111111010",
123508=>"000100100",
123509=>"001000101",
123510=>"111111111",
123511=>"000000000",
123512=>"000000001",
123513=>"000010011",
123514=>"000000101",
123515=>"010100000",
123516=>"000110100",
123517=>"111101010",
123518=>"000010100",
123519=>"000000001",
123520=>"000000010",
123521=>"111101100",
123522=>"111111101",
123523=>"111111101",
123524=>"000101111",
123525=>"110111001",
123526=>"001000000",
123527=>"000000000",
123528=>"001011001",
123529=>"000010000",
123530=>"111111000",
123531=>"011111110",
123532=>"001010000",
123533=>"010111111",
123534=>"110111111",
123535=>"000001000",
123536=>"111001001",
123537=>"101010111",
123538=>"101000001",
123539=>"000111111",
123540=>"000100001",
123541=>"000111010",
123542=>"110111111",
123543=>"100000000",
123544=>"011101110",
123545=>"001001000",
123546=>"000111111",
123547=>"010111000",
123548=>"111101100",
123549=>"001110111",
123550=>"110111001",
123551=>"101100111",
123552=>"001111101",
123553=>"111000000",
123554=>"010111111",
123555=>"110001000",
123556=>"101011111",
123557=>"100000000",
123558=>"001000001",
123559=>"111010000",
123560=>"011011000",
123561=>"000111110",
123562=>"111101100",
123563=>"001000000",
123564=>"111101101",
123565=>"010010010",
123566=>"010010011",
123567=>"010110110",
123568=>"101111111",
123569=>"101001100",
123570=>"011001001",
123571=>"001100100",
123572=>"011010100",
123573=>"111111000",
123574=>"101000000",
123575=>"000101101",
123576=>"111110000",
123577=>"010000000",
123578=>"110111101",
123579=>"010101111",
123580=>"100111110",
123581=>"111000100",
123582=>"101001101",
123583=>"011110110",
123584=>"000110010",
123585=>"111000000",
123586=>"111111110",
123587=>"000000110",
123588=>"000000011",
123589=>"100110001",
123590=>"110110011",
123591=>"101101101",
123592=>"101111101",
123593=>"110001101",
123594=>"000111111",
123595=>"110111111",
123596=>"110111110",
123597=>"101011011",
123598=>"001000000",
123599=>"001111010",
123600=>"001000011",
123601=>"001001000",
123602=>"000101001",
123603=>"010100111",
123604=>"101101111",
123605=>"000110100",
123606=>"111000000",
123607=>"010000101",
123608=>"000000100",
123609=>"000000001",
123610=>"100011001",
123611=>"000110100",
123612=>"001000001",
123613=>"101101000",
123614=>"010000000",
123615=>"010111101",
123616=>"000010011",
123617=>"011111111",
123618=>"111001101",
123619=>"000000101",
123620=>"101000010",
123621=>"111001011",
123622=>"101000111",
123623=>"101000000",
123624=>"010001100",
123625=>"101000101",
123626=>"000110100",
123627=>"001000000",
123628=>"000011111",
123629=>"000000001",
123630=>"001000100",
123631=>"000000000",
123632=>"000000100",
123633=>"011011000",
123634=>"000000111",
123635=>"100000001",
123636=>"010110010",
123637=>"000111111",
123638=>"000000010",
123639=>"000000100",
123640=>"111000000",
123641=>"111111110",
123642=>"000000001",
123643=>"000000100",
123644=>"111111111",
123645=>"111111111",
123646=>"001000101",
123647=>"111111111",
123648=>"111011111",
123649=>"010111010",
123650=>"100000101",
123651=>"111001101",
123652=>"101000000",
123653=>"111101110",
123654=>"101011101",
123655=>"011111101",
123656=>"000101101",
123657=>"111100110",
123658=>"000010100",
123659=>"110001000",
123660=>"111001000",
123661=>"110111000",
123662=>"000000000",
123663=>"110110110",
123664=>"111111100",
123665=>"111111001",
123666=>"111111000",
123667=>"011001001",
123668=>"001000000",
123669=>"111101101",
123670=>"001011111",
123671=>"111110110",
123672=>"101000000",
123673=>"111001111",
123674=>"011110110",
123675=>"000111111",
123676=>"101000000",
123677=>"001111000",
123678=>"011000101",
123679=>"110110100",
123680=>"111001001",
123681=>"001100111",
123682=>"110110100",
123683=>"110110001",
123684=>"011011011",
123685=>"000000000",
123686=>"111101101",
123687=>"011011000",
123688=>"111101111",
123689=>"000000000",
123690=>"100101000",
123691=>"000010000",
123692=>"011111101",
123693=>"110110000",
123694=>"111111111",
123695=>"011101000",
123696=>"111100000",
123697=>"111001001",
123698=>"110000100",
123699=>"001000000",
123700=>"101010010",
123701=>"000101111",
123702=>"010011010",
123703=>"010000000",
123704=>"111001101",
123705=>"000000000",
123706=>"000111100",
123707=>"000011110",
123708=>"110110111",
123709=>"101110110",
123710=>"000000100",
123711=>"000000101",
123712=>"011001000",
123713=>"000010110",
123714=>"110001101",
123715=>"100101001",
123716=>"000110111",
123717=>"000000100",
123718=>"000110000",
123719=>"000110110",
123720=>"111011111",
123721=>"000101101",
123722=>"010000001",
123723=>"111011010",
123724=>"000001101",
123725=>"000101100",
123726=>"000100100",
123727=>"000010100",
123728=>"010000111",
123729=>"111111010",
123730=>"000000000",
123731=>"000011011",
123732=>"110100111",
123733=>"110100011",
123734=>"111110110",
123735=>"110100000",
123736=>"110000100",
123737=>"011001000",
123738=>"001001001",
123739=>"001000000",
123740=>"000010111",
123741=>"011011010",
123742=>"111011111",
123743=>"001001111",
123744=>"011000000",
123745=>"010100110",
123746=>"010001101",
123747=>"100110000",
123748=>"100000000",
123749=>"111101000",
123750=>"101011110",
123751=>"000000000",
123752=>"111101111",
123753=>"000100010",
123754=>"111100101",
123755=>"001010110",
123756=>"110001000",
123757=>"000001000",
123758=>"000000001",
123759=>"011111111",
123760=>"001001000",
123761=>"111100000",
123762=>"000110111",
123763=>"100000000",
123764=>"010111000",
123765=>"100000000",
123766=>"111001000",
123767=>"101101000",
123768=>"111110110",
123769=>"011001110",
123770=>"111100001",
123771=>"000010101",
123772=>"001100100",
123773=>"100110110",
123774=>"101011110",
123775=>"010000010",
123776=>"111101000",
123777=>"110000000",
123778=>"000001100",
123779=>"001110100",
123780=>"000100111",
123781=>"111001000",
123782=>"100000001",
123783=>"111001001",
123784=>"100100100",
123785=>"000000011",
123786=>"011010000",
123787=>"110101100",
123788=>"000001111",
123789=>"000000100",
123790=>"111111101",
123791=>"001101000",
123792=>"001000000",
123793=>"000000100",
123794=>"111010010",
123795=>"011011000",
123796=>"111111000",
123797=>"000000000",
123798=>"010111000",
123799=>"110100100",
123800=>"011100011",
123801=>"000110110",
123802=>"111101101",
123803=>"000000001",
123804=>"101101101",
123805=>"111101111",
123806=>"010101011",
123807=>"101111111",
123808=>"001011011",
123809=>"101111010",
123810=>"111111010",
123811=>"111001000",
123812=>"111001001",
123813=>"000100100",
123814=>"000111000",
123815=>"111100111",
123816=>"111111111",
123817=>"110110000",
123818=>"000111110",
123819=>"011001111",
123820=>"111111101",
123821=>"111101001",
123822=>"110010011",
123823=>"110000000",
123824=>"110101000",
123825=>"111001111",
123826=>"101001010",
123827=>"100000000",
123828=>"001010000",
123829=>"111111111",
123830=>"100111110",
123831=>"111010111",
123832=>"110001110",
123833=>"100111001",
123834=>"111011000",
123835=>"111001110",
123836=>"100000010",
123837=>"010111111",
123838=>"100101101",
123839=>"000010000",
123840=>"011000000",
123841=>"010000100",
123842=>"000000001",
123843=>"111100100",
123844=>"111100000",
123845=>"001110100",
123846=>"000000011",
123847=>"111101101",
123848=>"110111111",
123849=>"000111100",
123850=>"101111000",
123851=>"000010011",
123852=>"001010001",
123853=>"110000000",
123854=>"000110000",
123855=>"001000000",
123856=>"110110000",
123857=>"110011011",
123858=>"010101100",
123859=>"000011111",
123860=>"011001001",
123861=>"110110110",
123862=>"010111010",
123863=>"111010000",
123864=>"000000000",
123865=>"100001000",
123866=>"000110110",
123867=>"000101101",
123868=>"011111101",
123869=>"000000101",
123870=>"111101000",
123871=>"111111101",
123872=>"000110110",
123873=>"010000101",
123874=>"110000000",
123875=>"111111011",
123876=>"111000000",
123877=>"000110111",
123878=>"111001000",
123879=>"111110110",
123880=>"111001100",
123881=>"010011011",
123882=>"100010010",
123883=>"101100101",
123884=>"001000100",
123885=>"110110010",
123886=>"111000101",
123887=>"011001000",
123888=>"110000000",
123889=>"011001011",
123890=>"000111010",
123891=>"000110100",
123892=>"111011101",
123893=>"000110010",
123894=>"001000000",
123895=>"011110000",
123896=>"111001000",
123897=>"101000010",
123898=>"000101011",
123899=>"000011010",
123900=>"111111111",
123901=>"000000000",
123902=>"000000001",
123903=>"000000000",
123904=>"001000100",
123905=>"000000000",
123906=>"000010010",
123907=>"000000001",
123908=>"000111011",
123909=>"100011111",
123910=>"010000000",
123911=>"000111111",
123912=>"010001101",
123913=>"000000010",
123914=>"001011111",
123915=>"010000000",
123916=>"110000000",
123917=>"011111100",
123918=>"100100111",
123919=>"111111111",
123920=>"100111111",
123921=>"000000000",
123922=>"000000000",
123923=>"100000000",
123924=>"111001011",
123925=>"000000111",
123926=>"100000001",
123927=>"101111111",
123928=>"101000000",
123929=>"010000000",
123930=>"001000000",
123931=>"000111110",
123932=>"111101100",
123933=>"111001111",
123934=>"101111111",
123935=>"011111101",
123936=>"100000011",
123937=>"000000101",
123938=>"101111011",
123939=>"001111111",
123940=>"011101101",
123941=>"001001011",
123942=>"000110111",
123943=>"110111000",
123944=>"100110010",
123945=>"000110110",
123946=>"100010111",
123947=>"000000000",
123948=>"010100100",
123949=>"111111111",
123950=>"010000000",
123951=>"000111001",
123952=>"111111110",
123953=>"001101111",
123954=>"001000000",
123955=>"111111000",
123956=>"000011111",
123957=>"001101111",
123958=>"100011011",
123959=>"010010000",
123960=>"000000000",
123961=>"010010011",
123962=>"111001000",
123963=>"101011100",
123964=>"010111001",
123965=>"111111110",
123966=>"111001000",
123967=>"001011111",
123968=>"100000000",
123969=>"011101111",
123970=>"111100000",
123971=>"000111111",
123972=>"011000000",
123973=>"011000101",
123974=>"000011001",
123975=>"000101000",
123976=>"110110111",
123977=>"000000001",
123978=>"111000000",
123979=>"000000010",
123980=>"111010000",
123981=>"001001001",
123982=>"100000010",
123983=>"111111001",
123984=>"101000000",
123985=>"111100000",
123986=>"111000000",
123987=>"001001000",
123988=>"111000000",
123989=>"100110110",
123990=>"110011001",
123991=>"101111110",
123992=>"110010010",
123993=>"000001111",
123994=>"001100110",
123995=>"110110100",
123996=>"000000000",
123997=>"110000000",
123998=>"000111111",
123999=>"100110101",
124000=>"111111111",
124001=>"110111101",
124002=>"111000000",
124003=>"111000011",
124004=>"011100101",
124005=>"011010000",
124006=>"011000000",
124007=>"101110100",
124008=>"000110100",
124009=>"111111100",
124010=>"110111100",
124011=>"011111111",
124012=>"101001000",
124013=>"001111011",
124014=>"000000000",
124015=>"100000100",
124016=>"001001011",
124017=>"011000010",
124018=>"001111110",
124019=>"101000111",
124020=>"000000000",
124021=>"000000000",
124022=>"000110110",
124023=>"000001111",
124024=>"010110010",
124025=>"011101000",
124026=>"011001001",
124027=>"001111100",
124028=>"010000001",
124029=>"110100000",
124030=>"010111000",
124031=>"000000000",
124032=>"000000000",
124033=>"000000000",
124034=>"001000100",
124035=>"111101111",
124036=>"111000000",
124037=>"011000111",
124038=>"100100110",
124039=>"000110010",
124040=>"100100010",
124041=>"000111111",
124042=>"100111000",
124043=>"111001000",
124044=>"000000000",
124045=>"000000100",
124046=>"100000110",
124047=>"010000000",
124048=>"111011001",
124049=>"010010110",
124050=>"000000111",
124051=>"011111010",
124052=>"100111110",
124053=>"101000100",
124054=>"000011111",
124055=>"100001001",
124056=>"011100110",
124057=>"000001011",
124058=>"000110110",
124059=>"100001000",
124060=>"000000000",
124061=>"010000000",
124062=>"000000001",
124063=>"101000111",
124064=>"100101110",
124065=>"001111000",
124066=>"001111111",
124067=>"101101111",
124068=>"111111110",
124069=>"101101101",
124070=>"001101111",
124071=>"000111111",
124072=>"111000111",
124073=>"100001101",
124074=>"111101100",
124075=>"000000000",
124076=>"111111100",
124077=>"110000000",
124078=>"010111001",
124079=>"111000010",
124080=>"011100100",
124081=>"111010100",
124082=>"000000000",
124083=>"000000100",
124084=>"111111111",
124085=>"101111100",
124086=>"011010000",
124087=>"011000000",
124088=>"011111100",
124089=>"000011010",
124090=>"000000000",
124091=>"000111100",
124092=>"111001100",
124093=>"100000010",
124094=>"001100110",
124095=>"000000000",
124096=>"111000000",
124097=>"000100010",
124098=>"111110000",
124099=>"110101100",
124100=>"000000000",
124101=>"111110001",
124102=>"010000000",
124103=>"000010000",
124104=>"111101000",
124105=>"000111010",
124106=>"101110010",
124107=>"000011011",
124108=>"000111111",
124109=>"111000101",
124110=>"000010010",
124111=>"111011000",
124112=>"000000110",
124113=>"000010110",
124114=>"000010110",
124115=>"011101111",
124116=>"111001100",
124117=>"010010001",
124118=>"000011000",
124119=>"000000101",
124120=>"000011111",
124121=>"011000000",
124122=>"001101110",
124123=>"111001000",
124124=>"001000000",
124125=>"100000101",
124126=>"101000101",
124127=>"000000000",
124128=>"111111000",
124129=>"111001000",
124130=>"110100110",
124131=>"011111111",
124132=>"111000000",
124133=>"100110010",
124134=>"011000011",
124135=>"111110000",
124136=>"110101000",
124137=>"000000011",
124138=>"100110110",
124139=>"001001000",
124140=>"000111111",
124141=>"110000000",
124142=>"101000000",
124143=>"000000000",
124144=>"110000100",
124145=>"011011010",
124146=>"111001001",
124147=>"100001101",
124148=>"000100000",
124149=>"001000101",
124150=>"101000000",
124151=>"000000000",
124152=>"000010010",
124153=>"100100101",
124154=>"111100111",
124155=>"011111101",
124156=>"100110010",
124157=>"111111000",
124158=>"110100101",
124159=>"011000000",
124160=>"000001001",
124161=>"101100011",
124162=>"000000101",
124163=>"111101111",
124164=>"100101011",
124165=>"110000000",
124166=>"100001000",
124167=>"101100000",
124168=>"000000000",
124169=>"000000100",
124170=>"000110000",
124171=>"010100011",
124172=>"101000100",
124173=>"000000000",
124174=>"101100000",
124175=>"011010000",
124176=>"000011001",
124177=>"110101010",
124178=>"100000000",
124179=>"101111101",
124180=>"000011000",
124181=>"000000001",
124182=>"110001101",
124183=>"010001000",
124184=>"001111001",
124185=>"000100100",
124186=>"000010010",
124187=>"101101110",
124188=>"000100000",
124189=>"000100100",
124190=>"111011101",
124191=>"000000000",
124192=>"100011011",
124193=>"000010000",
124194=>"011000010",
124195=>"111010000",
124196=>"111111011",
124197=>"101100000",
124198=>"000111111",
124199=>"111111111",
124200=>"010110110",
124201=>"000010110",
124202=>"011000001",
124203=>"111101000",
124204=>"001011011",
124205=>"011101000",
124206=>"001101100",
124207=>"000000000",
124208=>"000001001",
124209=>"000100110",
124210=>"000000010",
124211=>"000000111",
124212=>"000110111",
124213=>"110101100",
124214=>"000010110",
124215=>"000000000",
124216=>"011101000",
124217=>"101001000",
124218=>"101100110",
124219=>"101100111",
124220=>"001001000",
124221=>"010111101",
124222=>"001101000",
124223=>"111000000",
124224=>"101111011",
124225=>"010100010",
124226=>"111111111",
124227=>"110111111",
124228=>"011010010",
124229=>"000100101",
124230=>"110111010",
124231=>"010000001",
124232=>"000000000",
124233=>"000011011",
124234=>"000010001",
124235=>"110010111",
124236=>"000000000",
124237=>"100111000",
124238=>"000101101",
124239=>"000101000",
124240=>"010011010",
124241=>"110111111",
124242=>"110111010",
124243=>"001001001",
124244=>"111101101",
124245=>"100001110",
124246=>"111111100",
124247=>"001001100",
124248=>"110110000",
124249=>"101100100",
124250=>"001001000",
124251=>"111110100",
124252=>"010010010",
124253=>"011001001",
124254=>"101100111",
124255=>"001011111",
124256=>"011011010",
124257=>"010111110",
124258=>"101101100",
124259=>"110110000",
124260=>"110111110",
124261=>"010000000",
124262=>"110110011",
124263=>"000000000",
124264=>"010010001",
124265=>"000100100",
124266=>"111011110",
124267=>"000100000",
124268=>"000010111",
124269=>"010010010",
124270=>"000000111",
124271=>"011000000",
124272=>"100100101",
124273=>"111000000",
124274=>"100110111",
124275=>"101100111",
124276=>"111001000",
124277=>"100000100",
124278=>"111110101",
124279=>"011101111",
124280=>"000000000",
124281=>"111111100",
124282=>"011000001",
124283=>"101000100",
124284=>"100110111",
124285=>"000000000",
124286=>"000001111",
124287=>"010010010",
124288=>"101111101",
124289=>"100101101",
124290=>"101101111",
124291=>"111111100",
124292=>"000001001",
124293=>"111101111",
124294=>"001100101",
124295=>"110000000",
124296=>"011001111",
124297=>"010010000",
124298=>"011111011",
124299=>"100101111",
124300=>"100000011",
124301=>"000110000",
124302=>"111000000",
124303=>"000000000",
124304=>"001011001",
124305=>"110010000",
124306=>"000001111",
124307=>"010000001",
124308=>"101001000",
124309=>"100000100",
124310=>"010110111",
124311=>"011100110",
124312=>"010110000",
124313=>"101100100",
124314=>"100100101",
124315=>"100101000",
124316=>"111111111",
124317=>"111100001",
124318=>"111000000",
124319=>"100111000",
124320=>"100100111",
124321=>"100101111",
124322=>"101100000",
124323=>"111001000",
124324=>"101111100",
124325=>"010011111",
124326=>"101001011",
124327=>"000011010",
124328=>"111111111",
124329=>"111111010",
124330=>"000101101",
124331=>"000101111",
124332=>"111101111",
124333=>"111010110",
124334=>"001111111",
124335=>"010011010",
124336=>"101000001",
124337=>"011011011",
124338=>"111101011",
124339=>"101000001",
124340=>"110110111",
124341=>"011111000",
124342=>"001011000",
124343=>"011100000",
124344=>"000100000",
124345=>"110010000",
124346=>"111000000",
124347=>"100000001",
124348=>"000000000",
124349=>"001111111",
124350=>"111001001",
124351=>"111000000",
124352=>"001001101",
124353=>"111100001",
124354=>"100000000",
124355=>"100110100",
124356=>"111111011",
124357=>"100111011",
124358=>"000101111",
124359=>"110100100",
124360=>"000001110",
124361=>"100100101",
124362=>"111111010",
124363=>"111000101",
124364=>"011011111",
124365=>"001011111",
124366=>"000000000",
124367=>"011011001",
124368=>"000101111",
124369=>"111110010",
124370=>"010010000",
124371=>"000000010",
124372=>"100101111",
124373=>"110110110",
124374=>"011011000",
124375=>"101011011",
124376=>"101101101",
124377=>"010011000",
124378=>"101001101",
124379=>"000111000",
124380=>"001101011",
124381=>"001001000",
124382=>"110111010",
124383=>"000000100",
124384=>"000000011",
124385=>"010010010",
124386=>"101001101",
124387=>"111111100",
124388=>"000000000",
124389=>"000101111",
124390=>"011111110",
124391=>"000111111",
124392=>"000110110",
124393=>"000000000",
124394=>"010011011",
124395=>"111110010",
124396=>"110110111",
124397=>"011011000",
124398=>"000000000",
124399=>"000100100",
124400=>"110101000",
124401=>"001110110",
124402=>"011000111",
124403=>"001001001",
124404=>"011110100",
124405=>"111111111",
124406=>"000000101",
124407=>"010000100",
124408=>"101000000",
124409=>"000001110",
124410=>"111101000",
124411=>"111111011",
124412=>"101111111",
124413=>"111000000",
124414=>"011110100",
124415=>"000001000",
124416=>"110110100",
124417=>"000000010",
124418=>"101000000",
124419=>"110000010",
124420=>"000000001",
124421=>"111101000",
124422=>"000000110",
124423=>"110111111",
124424=>"000000101",
124425=>"000000111",
124426=>"011001000",
124427=>"010000010",
124428=>"101000000",
124429=>"001101111",
124430=>"100100100",
124431=>"101001010",
124432=>"111001000",
124433=>"111000000",
124434=>"110101001",
124435=>"000101011",
124436=>"100000000",
124437=>"000111111",
124438=>"000100111",
124439=>"101000100",
124440=>"100001000",
124441=>"001110000",
124442=>"000000111",
124443=>"000001101",
124444=>"000110000",
124445=>"011101001",
124446=>"000001001",
124447=>"000111010",
124448=>"000100101",
124449=>"000001111",
124450=>"000111111",
124451=>"100111110",
124452=>"000001011",
124453=>"000011100",
124454=>"000010011",
124455=>"000000000",
124456=>"100111111",
124457=>"111111000",
124458=>"111000111",
124459=>"010111011",
124460=>"111111010",
124461=>"111010010",
124462=>"110110000",
124463=>"100101000",
124464=>"101110000",
124465=>"000001111",
124466=>"000000000",
124467=>"101001111",
124468=>"101101111",
124469=>"111111001",
124470=>"011001000",
124471=>"000000000",
124472=>"111110100",
124473=>"000101000",
124474=>"111111000",
124475=>"100101100",
124476=>"011010001",
124477=>"011111001",
124478=>"111000001",
124479=>"100100010",
124480=>"000000011",
124481=>"000101100",
124482=>"111000101",
124483=>"100100000",
124484=>"111000011",
124485=>"100001000",
124486=>"000110111",
124487=>"110111011",
124488=>"001111111",
124489=>"011001011",
124490=>"111101000",
124491=>"000100001",
124492=>"000000010",
124493=>"100100111",
124494=>"000000110",
124495=>"111100000",
124496=>"111110000",
124497=>"110010000",
124498=>"001111010",
124499=>"111100001",
124500=>"010000101",
124501=>"000010010",
124502=>"000101101",
124503=>"111010000",
124504=>"001101110",
124505=>"011011000",
124506=>"111011010",
124507=>"000000000",
124508=>"010000000",
124509=>"000001001",
124510=>"010000011",
124511=>"011001001",
124512=>"111000101",
124513=>"001011111",
124514=>"111000000",
124515=>"111111001",
124516=>"011000000",
124517=>"011100001",
124518=>"111001111",
124519=>"010111000",
124520=>"011010111",
124521=>"010000000",
124522=>"000000010",
124523=>"101000011",
124524=>"000111110",
124525=>"111101111",
124526=>"100101100",
124527=>"000000001",
124528=>"100010110",
124529=>"000000000",
124530=>"110101001",
124531=>"010111001",
124532=>"010011111",
124533=>"101000000",
124534=>"001000101",
124535=>"101001011",
124536=>"111010000",
124537=>"010111111",
124538=>"000000000",
124539=>"111000111",
124540=>"110110110",
124541=>"011001001",
124542=>"101111111",
124543=>"111110101",
124544=>"101101101",
124545=>"111111100",
124546=>"000000101",
124547=>"000000000",
124548=>"011011010",
124549=>"111001000",
124550=>"100100001",
124551=>"000000000",
124552=>"011001001",
124553=>"001101111",
124554=>"111010010",
124555=>"111001000",
124556=>"000000111",
124557=>"111111111",
124558=>"010001001",
124559=>"001001000",
124560=>"111001111",
124561=>"000110111",
124562=>"000100110",
124563=>"111011101",
124564=>"100000001",
124565=>"101001000",
124566=>"101000000",
124567=>"000100001",
124568=>"010001100",
124569=>"100100010",
124570=>"101110000",
124571=>"111010010",
124572=>"110101111",
124573=>"111000001",
124574=>"111111101",
124575=>"001001001",
124576=>"000000110",
124577=>"000101111",
124578=>"011001111",
124579=>"000010000",
124580=>"110110010",
124581=>"101001100",
124582=>"001000010",
124583=>"101001111",
124584=>"010111100",
124585=>"101111111",
124586=>"111100000",
124587=>"111100000",
124588=>"110111111",
124589=>"111101000",
124590=>"011011110",
124591=>"101011111",
124592=>"000011010",
124593=>"110100111",
124594=>"011001111",
124595=>"000010010",
124596=>"011001010",
124597=>"111011111",
124598=>"011111101",
124599=>"000001111",
124600=>"110110100",
124601=>"000000010",
124602=>"111111010",
124603=>"011111111",
124604=>"011111110",
124605=>"111101111",
124606=>"001001001",
124607=>"100010010",
124608=>"111111101",
124609=>"000000011",
124610=>"001001010",
124611=>"100000101",
124612=>"101100111",
124613=>"010001001",
124614=>"011010000",
124615=>"110111100",
124616=>"111100101",
124617=>"111111010",
124618=>"111111100",
124619=>"000000111",
124620=>"000000000",
124621=>"011011001",
124622=>"101111001",
124623=>"000000000",
124624=>"101000001",
124625=>"011100110",
124626=>"000000000",
124627=>"100000000",
124628=>"100000000",
124629=>"001100101",
124630=>"111110000",
124631=>"101011000",
124632=>"000010111",
124633=>"000000010",
124634=>"111001101",
124635=>"111000111",
124636=>"000001100",
124637=>"111111000",
124638=>"000000000",
124639=>"000100110",
124640=>"111010100",
124641=>"111000000",
124642=>"100011111",
124643=>"100000110",
124644=>"001000001",
124645=>"111010010",
124646=>"111101111",
124647=>"110100101",
124648=>"010111111",
124649=>"000101001",
124650=>"100100001",
124651=>"110011011",
124652=>"000000101",
124653=>"000101111",
124654=>"000001000",
124655=>"110001111",
124656=>"101111111",
124657=>"100100100",
124658=>"000000000",
124659=>"100000110",
124660=>"001001101",
124661=>"110000000",
124662=>"111000000",
124663=>"011001001",
124664=>"100100101",
124665=>"111010111",
124666=>"011011000",
124667=>"001100110",
124668=>"000000000",
124669=>"000010111",
124670=>"011000000",
124671=>"000000101",
124672=>"001000001",
124673=>"110111110",
124674=>"111000111",
124675=>"110111111",
124676=>"000100000",
124677=>"011000110",
124678=>"101111100",
124679=>"101001111",
124680=>"000000000",
124681=>"111000001",
124682=>"100110011",
124683=>"111111000",
124684=>"101101101",
124685=>"100111100",
124686=>"000001110",
124687=>"111001111",
124688=>"110000101",
124689=>"111010111",
124690=>"101000000",
124691=>"110111111",
124692=>"111000110",
124693=>"100111011",
124694=>"111101100",
124695=>"111110111",
124696=>"000000000",
124697=>"111111111",
124698=>"111111111",
124699=>"000011000",
124700=>"110100110",
124701=>"000000000",
124702=>"111111111",
124703=>"000000000",
124704=>"000101101",
124705=>"101000000",
124706=>"000000000",
124707=>"111110100",
124708=>"000000000",
124709=>"000001001",
124710=>"000111111",
124711=>"101000000",
124712=>"111110010",
124713=>"000000000",
124714=>"111111000",
124715=>"000010110",
124716=>"100111110",
124717=>"111110001",
124718=>"111101000",
124719=>"000001010",
124720=>"111000000",
124721=>"000000000",
124722=>"110000111",
124723=>"111111111",
124724=>"000000000",
124725=>"111111000",
124726=>"010000011",
124727=>"000000000",
124728=>"010111111",
124729=>"000001101",
124730=>"110000010",
124731=>"000000100",
124732=>"111111111",
124733=>"111000000",
124734=>"000011000",
124735=>"001011111",
124736=>"111111001",
124737=>"000110010",
124738=>"111111111",
124739=>"100110010",
124740=>"111000000",
124741=>"100001111",
124742=>"000111111",
124743=>"111110010",
124744=>"100011011",
124745=>"111111111",
124746=>"010000011",
124747=>"000001000",
124748=>"111000000",
124749=>"000000000",
124750=>"000000000",
124751=>"100101101",
124752=>"000010000",
124753=>"111010100",
124754=>"111100101",
124755=>"001100110",
124756=>"111010000",
124757=>"111111101",
124758=>"000010100",
124759=>"101101101",
124760=>"010001000",
124761=>"000000011",
124762=>"000001011",
124763=>"111111111",
124764=>"111011111",
124765=>"000000010",
124766=>"111111111",
124767=>"010010111",
124768=>"111111111",
124769=>"101101111",
124770=>"010000010",
124771=>"000100110",
124772=>"000000000",
124773=>"111000011",
124774=>"011111111",
124775=>"111001011",
124776=>"010001011",
124777=>"111111111",
124778=>"111111111",
124779=>"000000111",
124780=>"101001111",
124781=>"010010011",
124782=>"100000000",
124783=>"010000110",
124784=>"000000000",
124785=>"110111111",
124786=>"100000110",
124787=>"001001111",
124788=>"111000010",
124789=>"000101110",
124790=>"111111111",
124791=>"001111001",
124792=>"111111111",
124793=>"011001110",
124794=>"110000010",
124795=>"000000000",
124796=>"000000000",
124797=>"000000000",
124798=>"000000000",
124799=>"000000000",
124800=>"111111010",
124801=>"111000000",
124802=>"111111111",
124803=>"111010000",
124804=>"111000000",
124805=>"000010010",
124806=>"001100100",
124807=>"100100100",
124808=>"000000000",
124809=>"000000000",
124810=>"111111100",
124811=>"001001111",
124812=>"001111111",
124813=>"000001001",
124814=>"011111101",
124815=>"001001001",
124816=>"000001001",
124817=>"000000110",
124818=>"000101111",
124819=>"000000101",
124820=>"000000001",
124821=>"111000111",
124822=>"111100111",
124823=>"000000000",
124824=>"011110110",
124825=>"110111011",
124826=>"111110000",
124827=>"000010010",
124828=>"100111100",
124829=>"111110010",
124830=>"110111111",
124831=>"000000111",
124832=>"111001000",
124833=>"011000001",
124834=>"111001000",
124835=>"111011111",
124836=>"111111010",
124837=>"000001000",
124838=>"100111111",
124839=>"010111111",
124840=>"111000000",
124841=>"000000111",
124842=>"110000000",
124843=>"010000010",
124844=>"000011011",
124845=>"010010000",
124846=>"000000000",
124847=>"111111111",
124848=>"000000111",
124849=>"000000100",
124850=>"000000000",
124851=>"010000010",
124852=>"010110110",
124853=>"110000001",
124854=>"111111110",
124855=>"000111100",
124856=>"111111111",
124857=>"001001000",
124858=>"101111111",
124859=>"111000001",
124860=>"000111110",
124861=>"111110111",
124862=>"000110110",
124863=>"110000000",
124864=>"111100101",
124865=>"010110111",
124866=>"111000111",
124867=>"000000000",
124868=>"000001000",
124869=>"001011001",
124870=>"001100111",
124871=>"111110010",
124872=>"111011001",
124873=>"000001000",
124874=>"011001001",
124875=>"011111111",
124876=>"000111011",
124877=>"110001000",
124878=>"000000010",
124879=>"011001111",
124880=>"000000000",
124881=>"000000100",
124882=>"111111100",
124883=>"010100001",
124884=>"000111100",
124885=>"000100100",
124886=>"111101110",
124887=>"111101111",
124888=>"101101101",
124889=>"110011101",
124890=>"011000000",
124891=>"111010000",
124892=>"111011011",
124893=>"110010011",
124894=>"010101100",
124895=>"111111101",
124896=>"000010111",
124897=>"111000111",
124898=>"111001000",
124899=>"011011010",
124900=>"000011111",
124901=>"010111111",
124902=>"000101110",
124903=>"000000000",
124904=>"111110111",
124905=>"111101110",
124906=>"011011110",
124907=>"111111111",
124908=>"000001111",
124909=>"111001000",
124910=>"100000000",
124911=>"000000111",
124912=>"101111111",
124913=>"111111100",
124914=>"101001000",
124915=>"001011110",
124916=>"000100000",
124917=>"000101110",
124918=>"101001100",
124919=>"111111010",
124920=>"111111101",
124921=>"000000100",
124922=>"111010100",
124923=>"000000000",
124924=>"110010000",
124925=>"100111000",
124926=>"000000000",
124927=>"000111110",
124928=>"011001101",
124929=>"000100110",
124930=>"101101111",
124931=>"000000010",
124932=>"100000011",
124933=>"000000110",
124934=>"011111000",
124935=>"011000100",
124936=>"010001100",
124937=>"101100000",
124938=>"100101001",
124939=>"110010000",
124940=>"010111110",
124941=>"010011000",
124942=>"101111011",
124943=>"111000001",
124944=>"100000101",
124945=>"000111111",
124946=>"000000000",
124947=>"000000000",
124948=>"101100000",
124949=>"101000111",
124950=>"001011100",
124951=>"101010001",
124952=>"001101001",
124953=>"000101111",
124954=>"111100111",
124955=>"111101100",
124956=>"000101000",
124957=>"000000000",
124958=>"011010010",
124959=>"001011000",
124960=>"010111101",
124961=>"010010000",
124962=>"010100000",
124963=>"000101111",
124964=>"110110100",
124965=>"001100110",
124966=>"000000111",
124967=>"000111010",
124968=>"000111111",
124969=>"011111000",
124970=>"000010001",
124971=>"000000101",
124972=>"111110001",
124973=>"000101011",
124974=>"011000111",
124975=>"011010111",
124976=>"010000000",
124977=>"000011001",
124978=>"111111010",
124979=>"000000110",
124980=>"000000000",
124981=>"100000100",
124982=>"010100101",
124983=>"000101111",
124984=>"111000010",
124985=>"000000000",
124986=>"000111000",
124987=>"000000000",
124988=>"110110000",
124989=>"111111101",
124990=>"000000001",
124991=>"001001110",
124992=>"000101000",
124993=>"101110110",
124994=>"000111111",
124995=>"000001000",
124996=>"001010011",
124997=>"100000010",
124998=>"011110100",
124999=>"110101101",
125000=>"001111001",
125001=>"011100000",
125002=>"000010001",
125003=>"111101111",
125004=>"100000000",
125005=>"011011101",
125006=>"000100100",
125007=>"000010111",
125008=>"101111001",
125009=>"111101001",
125010=>"111000010",
125011=>"011001010",
125012=>"100101101",
125013=>"000100011",
125014=>"011011011",
125015=>"001001111",
125016=>"100101000",
125017=>"001011011",
125018=>"110000001",
125019=>"000011001",
125020=>"000000010",
125021=>"001001110",
125022=>"011011010",
125023=>"000000001",
125024=>"000100000",
125025=>"010000000",
125026=>"111100101",
125027=>"100100111",
125028=>"101101001",
125029=>"010100100",
125030=>"000000010",
125031=>"111111000",
125032=>"000101110",
125033=>"101111101",
125034=>"111110110",
125035=>"010110100",
125036=>"001000111",
125037=>"011010010",
125038=>"011010000",
125039=>"000000000",
125040=>"110110000",
125041=>"000011010",
125042=>"000000111",
125043=>"001001000",
125044=>"101111111",
125045=>"000100010",
125046=>"111111110",
125047=>"110010000",
125048=>"101000011",
125049=>"101101111",
125050=>"000011111",
125051=>"000011000",
125052=>"000110110",
125053=>"110100001",
125054=>"010010101",
125055=>"101101101",
125056=>"010000000",
125057=>"110000001",
125058=>"111010000",
125059=>"001010111",
125060=>"000000111",
125061=>"111111000",
125062=>"100000101",
125063=>"001001001",
125064=>"011001000",
125065=>"110110000",
125066=>"101000101",
125067=>"011010000",
125068=>"000000000",
125069=>"101000111",
125070=>"000010010",
125071=>"000000101",
125072=>"110110111",
125073=>"001111101",
125074=>"001000000",
125075=>"000000001",
125076=>"000101101",
125077=>"001000110",
125078=>"111110001",
125079=>"110111100",
125080=>"010000010",
125081=>"000010010",
125082=>"111100000",
125083=>"001100111",
125084=>"011010111",
125085=>"010000000",
125086=>"110010011",
125087=>"101000111",
125088=>"011111000",
125089=>"111001100",
125090=>"111110000",
125091=>"101111111",
125092=>"010000101",
125093=>"000100100",
125094=>"110110000",
125095=>"000000111",
125096=>"000000011",
125097=>"000101101",
125098=>"000100011",
125099=>"000000001",
125100=>"010011000",
125101=>"000101101",
125102=>"001000010",
125103=>"000010111",
125104=>"000000010",
125105=>"000110110",
125106=>"001000000",
125107=>"100110100",
125108=>"001011010",
125109=>"111101111",
125110=>"111000000",
125111=>"010011000",
125112=>"001001000",
125113=>"000101100",
125114=>"010010000",
125115=>"101111111",
125116=>"000010110",
125117=>"110100000",
125118=>"001000011",
125119=>"000010010",
125120=>"000101111",
125121=>"001101011",
125122=>"101111111",
125123=>"011111111",
125124=>"000011010",
125125=>"010001000",
125126=>"000000000",
125127=>"010111100",
125128=>"111111010",
125129=>"101000101",
125130=>"101011010",
125131=>"111111010",
125132=>"000000000",
125133=>"000011110",
125134=>"111111101",
125135=>"000110011",
125136=>"101111111",
125137=>"100110100",
125138=>"000010111",
125139=>"101010000",
125140=>"010000000",
125141=>"110111011",
125142=>"000000111",
125143=>"110000100",
125144=>"001000000",
125145=>"001000111",
125146=>"100111100",
125147=>"111101111",
125148=>"100100000",
125149=>"000001010",
125150=>"011101010",
125151=>"010000000",
125152=>"101101101",
125153=>"010101110",
125154=>"010010010",
125155=>"010100111",
125156=>"001101111",
125157=>"000100111",
125158=>"111000010",
125159=>"010100010",
125160=>"000010000",
125161=>"111000110",
125162=>"001000100",
125163=>"101101101",
125164=>"101101111",
125165=>"010010000",
125166=>"101000000",
125167=>"000001101",
125168=>"101000111",
125169=>"110101100",
125170=>"000010111",
125171=>"100110110",
125172=>"010111010",
125173=>"111111111",
125174=>"000010000",
125175=>"000010011",
125176=>"000010010",
125177=>"010010001",
125178=>"000001000",
125179=>"100001011",
125180=>"111011000",
125181=>"000000111",
125182=>"011011011",
125183=>"000000111",
125184=>"111111011",
125185=>"000000000",
125186=>"000000101",
125187=>"010010000",
125188=>"111100100",
125189=>"101000110",
125190=>"111101101",
125191=>"000110011",
125192=>"011001000",
125193=>"000000001",
125194=>"001000000",
125195=>"101101000",
125196=>"000010000",
125197=>"001000000",
125198=>"011111011",
125199=>"101111010",
125200=>"000111000",
125201=>"111000000",
125202=>"100000000",
125203=>"000001011",
125204=>"100000000",
125205=>"000000100",
125206=>"111000000",
125207=>"111111110",
125208=>"000111110",
125209=>"111001101",
125210=>"100000000",
125211=>"011000000",
125212=>"000111000",
125213=>"010000000",
125214=>"111111010",
125215=>"111110000",
125216=>"010101000",
125217=>"110101010",
125218=>"111101000",
125219=>"000010000",
125220=>"100000000",
125221=>"111010000",
125222=>"000010110",
125223=>"001011100",
125224=>"000001000",
125225=>"111001001",
125226=>"001011001",
125227=>"111111111",
125228=>"001111001",
125229=>"101001111",
125230=>"111111001",
125231=>"111001111",
125232=>"110000000",
125233=>"010100100",
125234=>"100110100",
125235=>"100111010",
125236=>"001001111",
125237=>"001011110",
125238=>"110000001",
125239=>"000010000",
125240=>"110101000",
125241=>"001001000",
125242=>"100100101",
125243=>"001001010",
125244=>"100010100",
125245=>"010101101",
125246=>"000000000",
125247=>"011000000",
125248=>"001110111",
125249=>"011010000",
125250=>"000111111",
125251=>"001001001",
125252=>"000000111",
125253=>"010000100",
125254=>"001000001",
125255=>"110010111",
125256=>"010100100",
125257=>"010010010",
125258=>"001101001",
125259=>"000001111",
125260=>"001111010",
125261=>"100100110",
125262=>"001011011",
125263=>"100111111",
125264=>"110010000",
125265=>"111000010",
125266=>"000010000",
125267=>"011001110",
125268=>"000000111",
125269=>"100011100",
125270=>"011011000",
125271=>"000101100",
125272=>"001000000",
125273=>"001101000",
125274=>"111011000",
125275=>"011101100",
125276=>"110111000",
125277=>"001101000",
125278=>"000000101",
125279=>"100100000",
125280=>"000010110",
125281=>"110000000",
125282=>"000010111",
125283=>"100001011",
125284=>"100111100",
125285=>"111110110",
125286=>"001000110",
125287=>"000000000",
125288=>"100111111",
125289=>"111111111",
125290=>"000000111",
125291=>"111101111",
125292=>"111100000",
125293=>"111111011",
125294=>"001000000",
125295=>"111111000",
125296=>"100011001",
125297=>"111111000",
125298=>"001000110",
125299=>"110111111",
125300=>"000111111",
125301=>"000000100",
125302=>"000110111",
125303=>"001000100",
125304=>"101010010",
125305=>"000111111",
125306=>"110000000",
125307=>"101000001",
125308=>"000100110",
125309=>"100100010",
125310=>"010111111",
125311=>"111000110",
125312=>"010111011",
125313=>"111101000",
125314=>"111000000",
125315=>"111110011",
125316=>"000111111",
125317=>"000001011",
125318=>"110011000",
125319=>"000110000",
125320=>"101100101",
125321=>"010110100",
125322=>"110100100",
125323=>"101100111",
125324=>"001000001",
125325=>"111101111",
125326=>"111110000",
125327=>"110001001",
125328=>"101011000",
125329=>"010111000",
125330=>"001001011",
125331=>"000010010",
125332=>"000011111",
125333=>"000111010",
125334=>"110111011",
125335=>"111110100",
125336=>"110111000",
125337=>"000000010",
125338=>"110111111",
125339=>"000000000",
125340=>"110000000",
125341=>"000111111",
125342=>"111110000",
125343=>"000110111",
125344=>"000010000",
125345=>"111111010",
125346=>"001000101",
125347=>"101111111",
125348=>"001011001",
125349=>"011011011",
125350=>"100001011",
125351=>"001110110",
125352=>"111100101",
125353=>"001100111",
125354=>"111100000",
125355=>"110000000",
125356=>"111111111",
125357=>"011111110",
125358=>"010110011",
125359=>"010110111",
125360=>"010000000",
125361=>"011001111",
125362=>"011000000",
125363=>"001001000",
125364=>"000110110",
125365=>"000100111",
125366=>"100001101",
125367=>"010110100",
125368=>"001010001",
125369=>"000110111",
125370=>"110110101",
125371=>"101001101",
125372=>"010111010",
125373=>"000100111",
125374=>"111100100",
125375=>"101001101",
125376=>"001000101",
125377=>"000000000",
125378=>"010000110",
125379=>"000000100",
125380=>"010010111",
125381=>"111111011",
125382=>"111111000",
125383=>"000001101",
125384=>"101111101",
125385=>"000001111",
125386=>"110111111",
125387=>"010000101",
125388=>"101000010",
125389=>"001011011",
125390=>"011001010",
125391=>"110011111",
125392=>"000000000",
125393=>"110011111",
125394=>"000010001",
125395=>"111111110",
125396=>"000100111",
125397=>"010100110",
125398=>"000000000",
125399=>"000000111",
125400=>"101111001",
125401=>"000000000",
125402=>"000110100",
125403=>"001110000",
125404=>"011001000",
125405=>"100100011",
125406=>"000000000",
125407=>"001000000",
125408=>"000000000",
125409=>"110000000",
125410=>"010010000",
125411=>"011111100",
125412=>"000001111",
125413=>"011000001",
125414=>"111000000",
125415=>"011011101",
125416=>"000000010",
125417=>"100101111",
125418=>"000000011",
125419=>"111111111",
125420=>"000001000",
125421=>"110101111",
125422=>"000000000",
125423=>"100100000",
125424=>"000000010",
125425=>"011111100",
125426=>"111100000",
125427=>"001011011",
125428=>"110110111",
125429=>"011101000",
125430=>"001000011",
125431=>"010011010",
125432=>"111000000",
125433=>"111000000",
125434=>"111100100",
125435=>"000111111",
125436=>"111111111",
125437=>"111100101",
125438=>"001001001",
125439=>"000110111",
125440=>"100000010",
125441=>"110000010",
125442=>"001010000",
125443=>"000000000",
125444=>"100000111",
125445=>"001111000",
125446=>"011110000",
125447=>"101101000",
125448=>"110110101",
125449=>"000010010",
125450=>"110111011",
125451=>"111000000",
125452=>"000000001",
125453=>"000000000",
125454=>"011111001",
125455=>"111110110",
125456=>"101111110",
125457=>"010111110",
125458=>"000100000",
125459=>"000010111",
125460=>"001101011",
125461=>"000001111",
125462=>"010011011",
125463=>"000111111",
125464=>"011101010",
125465=>"000000110",
125466=>"000101111",
125467=>"000000001",
125468=>"011110111",
125469=>"000111001",
125470=>"011000000",
125471=>"110111100",
125472=>"000000101",
125473=>"000000010",
125474=>"010010110",
125475=>"000000001",
125476=>"010110110",
125477=>"000001000",
125478=>"001001111",
125479=>"001111101",
125480=>"000111111",
125481=>"111110000",
125482=>"000010010",
125483=>"010000000",
125484=>"111111001",
125485=>"101111111",
125486=>"000101101",
125487=>"000000110",
125488=>"100111110",
125489=>"100000011",
125490=>"111000010",
125491=>"010110111",
125492=>"000001111",
125493=>"000111111",
125494=>"000111010",
125495=>"000000111",
125496=>"110111001",
125497=>"000101111",
125498=>"101111101",
125499=>"010010110",
125500=>"110101111",
125501=>"111111010",
125502=>"100110000",
125503=>"110100011",
125504=>"111111111",
125505=>"110000001",
125506=>"001111100",
125507=>"100000111",
125508=>"111000000",
125509=>"111111101",
125510=>"011010000",
125511=>"000000000",
125512=>"001011011",
125513=>"000000001",
125514=>"111001000",
125515=>"100111111",
125516=>"111110000",
125517=>"011011111",
125518=>"111000100",
125519=>"111001001",
125520=>"010110010",
125521=>"010000000",
125522=>"010111001",
125523=>"000000101",
125524=>"001110110",
125525=>"111000000",
125526=>"000100000",
125527=>"110000000",
125528=>"111001000",
125529=>"100110000",
125530=>"111111000",
125531=>"111110111",
125532=>"000000000",
125533=>"100000001",
125534=>"000000110",
125535=>"011001110",
125536=>"010000101",
125537=>"010000000",
125538=>"111001000",
125539=>"111011101",
125540=>"010101101",
125541=>"011111100",
125542=>"000001111",
125543=>"010101111",
125544=>"001010010",
125545=>"011101101",
125546=>"110111011",
125547=>"000101000",
125548=>"001001000",
125549=>"110011101",
125550=>"111111000",
125551=>"110000001",
125552=>"101000110",
125553=>"001111001",
125554=>"001111011",
125555=>"110000000",
125556=>"101101111",
125557=>"101101101",
125558=>"111110010",
125559=>"111111111",
125560=>"000000101",
125561=>"010000000",
125562=>"111111000",
125563=>"000000111",
125564=>"100101101",
125565=>"000100101",
125566=>"011000100",
125567=>"110000000",
125568=>"110100110",
125569=>"010010001",
125570=>"010100001",
125571=>"000000101",
125572=>"101001101",
125573=>"111111011",
125574=>"001100100",
125575=>"100011001",
125576=>"101001001",
125577=>"010101110",
125578=>"010000000",
125579=>"111000101",
125580=>"001000111",
125581=>"010000000",
125582=>"111000101",
125583=>"111100100",
125584=>"100100011",
125585=>"000111111",
125586=>"000000010",
125587=>"101001001",
125588=>"001000010",
125589=>"110111000",
125590=>"111110010",
125591=>"111111000",
125592=>"110110000",
125593=>"010000010",
125594=>"001000111",
125595=>"100000100",
125596=>"111110001",
125597=>"110000000",
125598=>"111000111",
125599=>"011001000",
125600=>"100111001",
125601=>"111111000",
125602=>"110000000",
125603=>"011011010",
125604=>"000111010",
125605=>"001011110",
125606=>"001111111",
125607=>"111111000",
125608=>"010111111",
125609=>"000000001",
125610=>"000111110",
125611=>"001110000",
125612=>"011111110",
125613=>"110111000",
125614=>"010100000",
125615=>"111000000",
125616=>"011000001",
125617=>"110110010",
125618=>"000001000",
125619=>"111000000",
125620=>"011001001",
125621=>"000111010",
125622=>"000100100",
125623=>"000010000",
125624=>"011011000",
125625=>"100000010",
125626=>"000000000",
125627=>"100001000",
125628=>"101101111",
125629=>"111000111",
125630=>"011111101",
125631=>"000000101",
125632=>"000101111",
125633=>"111111010",
125634=>"000011101",
125635=>"001011000",
125636=>"111001111",
125637=>"111001000",
125638=>"111111000",
125639=>"011000010",
125640=>"000011111",
125641=>"001000001",
125642=>"000001011",
125643=>"000111111",
125644=>"000000000",
125645=>"011010011",
125646=>"101010000",
125647=>"001100000",
125648=>"110010000",
125649=>"101000110",
125650=>"001000000",
125651=>"110100010",
125652=>"001001101",
125653=>"001011110",
125654=>"111101000",
125655=>"010001000",
125656=>"000101111",
125657=>"101001111",
125658=>"011010111",
125659=>"101111110",
125660=>"110110000",
125661=>"001000000",
125662=>"101101101",
125663=>"110101001",
125664=>"011100100",
125665=>"011111101",
125666=>"010000101",
125667=>"000110111",
125668=>"000000000",
125669=>"010000011",
125670=>"001101111",
125671=>"100010000",
125672=>"001111000",
125673=>"101101010",
125674=>"111101110",
125675=>"110111111",
125676=>"101111101",
125677=>"101000111",
125678=>"000000000",
125679=>"111001101",
125680=>"001000010",
125681=>"011000000",
125682=>"011111101",
125683=>"100000111",
125684=>"011000100",
125685=>"101101000",
125686=>"111000000",
125687=>"000100100",
125688=>"001100110",
125689=>"001111111",
125690=>"110110000",
125691=>"000111101",
125692=>"000111111",
125693=>"010000000",
125694=>"111101100",
125695=>"010001001",
125696=>"011011001",
125697=>"111000000",
125698=>"101000101",
125699=>"110000110",
125700=>"100111111",
125701=>"010000000",
125702=>"000000101",
125703=>"111111000",
125704=>"110000001",
125705=>"000000101",
125706=>"101000010",
125707=>"110110110",
125708=>"000000000",
125709=>"000110110",
125710=>"100110010",
125711=>"111001000",
125712=>"111110100",
125713=>"111001000",
125714=>"110111110",
125715=>"110000000",
125716=>"100000001",
125717=>"000000001",
125718=>"000001111",
125719=>"111000000",
125720=>"000001001",
125721=>"000110000",
125722=>"000110010",
125723=>"000010101",
125724=>"000101110",
125725=>"000101010",
125726=>"010011011",
125727=>"010010011",
125728=>"000110111",
125729=>"100110110",
125730=>"000000000",
125731=>"101000111",
125732=>"101100100",
125733=>"010110100",
125734=>"010111000",
125735=>"100110110",
125736=>"111111000",
125737=>"001001000",
125738=>"011000111",
125739=>"000011010",
125740=>"001100000",
125741=>"100110101",
125742=>"111000001",
125743=>"111010111",
125744=>"000000000",
125745=>"001111011",
125746=>"110111111",
125747=>"111001000",
125748=>"000000100",
125749=>"000000000",
125750=>"000000001",
125751=>"111001101",
125752=>"001000001",
125753=>"000000000",
125754=>"101001101",
125755=>"000000000",
125756=>"110110110",
125757=>"100111111",
125758=>"000000000",
125759=>"010110110",
125760=>"000001001",
125761=>"111111101",
125762=>"101000001",
125763=>"100111011",
125764=>"101001111",
125765=>"010110110",
125766=>"010101110",
125767=>"000110010",
125768=>"010111110",
125769=>"000110010",
125770=>"111110111",
125771=>"111111111",
125772=>"110000111",
125773=>"101001001",
125774=>"100101100",
125775=>"111101000",
125776=>"101110111",
125777=>"111111111",
125778=>"111011111",
125779=>"011011001",
125780=>"001000000",
125781=>"110010110",
125782=>"011011011",
125783=>"001111001",
125784=>"100110110",
125785=>"001111011",
125786=>"001011111",
125787=>"110110111",
125788=>"101001001",
125789=>"000000011",
125790=>"001001001",
125791=>"110111101",
125792=>"000000000",
125793=>"000110010",
125794=>"101000101",
125795=>"000100110",
125796=>"111111110",
125797=>"101000000",
125798=>"110110000",
125799=>"001001101",
125800=>"000101111",
125801=>"111111000",
125802=>"111001111",
125803=>"110111111",
125804=>"001111011",
125805=>"001001001",
125806=>"000000000",
125807=>"000000111",
125808=>"000100100",
125809=>"011011111",
125810=>"001001100",
125811=>"000101111",
125812=>"001000111",
125813=>"000000000",
125814=>"001000111",
125815=>"000111001",
125816=>"000000000",
125817=>"000001011",
125818=>"111111111",
125819=>"000000000",
125820=>"100101110",
125821=>"010100000",
125822=>"010110110",
125823=>"110110110",
125824=>"010010100",
125825=>"110110000",
125826=>"111000101",
125827=>"000000101",
125828=>"111110000",
125829=>"000000101",
125830=>"000010011",
125831=>"000100010",
125832=>"100001001",
125833=>"000011010",
125834=>"000100100",
125835=>"110010000",
125836=>"001000001",
125837=>"000001000",
125838=>"000000101",
125839=>"000000000",
125840=>"000000100",
125841=>"000111000",
125842=>"111110000",
125843=>"000100110",
125844=>"100111110",
125845=>"111000001",
125846=>"111001001",
125847=>"000000010",
125848=>"010111110",
125849=>"111011001",
125850=>"010111110",
125851=>"000000000",
125852=>"011101101",
125853=>"001111011",
125854=>"000001100",
125855=>"111001101",
125856=>"110110010",
125857=>"010000000",
125858=>"000001111",
125859=>"111001000",
125860=>"001000010",
125861=>"011001010",
125862=>"001111010",
125863=>"100100100",
125864=>"011111000",
125865=>"111111010",
125866=>"010000110",
125867=>"111000000",
125868=>"111111101",
125869=>"000000101",
125870=>"100101011",
125871=>"011000001",
125872=>"001000000",
125873=>"011010100",
125874=>"000101110",
125875=>"010000111",
125876=>"110101110",
125877=>"101001001",
125878=>"000110110",
125879=>"000111111",
125880=>"010011011",
125881=>"001111111",
125882=>"110111111",
125883=>"000000110",
125884=>"000100000",
125885=>"110110000",
125886=>"010001000",
125887=>"000001101",
125888=>"111000000",
125889=>"000000111",
125890=>"111111110",
125891=>"001100100",
125892=>"001000000",
125893=>"110111101",
125894=>"111101111",
125895=>"010000001",
125896=>"000000010",
125897=>"010000000",
125898=>"000001101",
125899=>"101000000",
125900=>"010010000",
125901=>"001111110",
125902=>"001101101",
125903=>"000111111",
125904=>"100010000",
125905=>"000110100",
125906=>"110111111",
125907=>"001001000",
125908=>"110110000",
125909=>"001000000",
125910=>"110001000",
125911=>"000000111",
125912=>"001001001",
125913=>"010010000",
125914=>"000011100",
125915=>"101001001",
125916=>"010100010",
125917=>"001011011",
125918=>"110111110",
125919=>"111110101",
125920=>"111000000",
125921=>"101011101",
125922=>"000111110",
125923=>"001101000",
125924=>"101000000",
125925=>"101001001",
125926=>"101001110",
125927=>"000010000",
125928=>"000000100",
125929=>"000000101",
125930=>"001000010",
125931=>"001001111",
125932=>"000010000",
125933=>"001000000",
125934=>"000101000",
125935=>"010110110",
125936=>"111000001",
125937=>"101110010",
125938=>"010000111",
125939=>"100100110",
125940=>"110110011",
125941=>"000000011",
125942=>"010110000",
125943=>"000111111",
125944=>"000111110",
125945=>"111101000",
125946=>"111111111",
125947=>"000111111",
125948=>"000100111",
125949=>"001000010",
125950=>"001111110",
125951=>"111100111",
125952=>"001000100",
125953=>"101110000",
125954=>"100000101",
125955=>"011111000",
125956=>"011001000",
125957=>"000101100",
125958=>"000000000",
125959=>"001000111",
125960=>"111110111",
125961=>"000000111",
125962=>"111011110",
125963=>"000101100",
125964=>"111010010",
125965=>"111010010",
125966=>"011011000",
125967=>"111101111",
125968=>"110010010",
125969=>"000101000",
125970=>"000101110",
125971=>"100000011",
125972=>"100000000",
125973=>"000111111",
125974=>"111100100",
125975=>"010111110",
125976=>"100000000",
125977=>"110000110",
125978=>"001000101",
125979=>"111010110",
125980=>"000000111",
125981=>"101111000",
125982=>"000001010",
125983=>"111000000",
125984=>"000000000",
125985=>"111111010",
125986=>"001101010",
125987=>"000000000",
125988=>"010001001",
125989=>"100101001",
125990=>"011110100",
125991=>"000011101",
125992=>"100110100",
125993=>"000010111",
125994=>"101000001",
125995=>"000000010",
125996=>"000101001",
125997=>"000100000",
125998=>"010100010",
125999=>"010001000",
126000=>"111111000",
126001=>"001001001",
126002=>"000111111",
126003=>"101110110",
126004=>"100100100",
126005=>"010110110",
126006=>"010110001",
126007=>"101000000",
126008=>"101000110",
126009=>"101101111",
126010=>"101101000",
126011=>"111011111",
126012=>"100100011",
126013=>"011000011",
126014=>"000000000",
126015=>"000100100",
126016=>"111111111",
126017=>"000101000",
126018=>"111111010",
126019=>"100100000",
126020=>"101111000",
126021=>"000000000",
126022=>"111101000",
126023=>"010100000",
126024=>"011111111",
126025=>"111111111",
126026=>"000101100",
126027=>"000000001",
126028=>"000000001",
126029=>"010101111",
126030=>"000001100",
126031=>"101100110",
126032=>"001111000",
126033=>"010111110",
126034=>"111111000",
126035=>"110000000",
126036=>"010000100",
126037=>"000010111",
126038=>"111001100",
126039=>"000000111",
126040=>"111111111",
126041=>"111100001",
126042=>"100000000",
126043=>"111100100",
126044=>"000000000",
126045=>"001011010",
126046=>"011000111",
126047=>"001001000",
126048=>"010010000",
126049=>"010010010",
126050=>"000000111",
126051=>"001000000",
126052=>"110010000",
126053=>"111100111",
126054=>"101110110",
126055=>"111000101",
126056=>"111111000",
126057=>"000111111",
126058=>"101000011",
126059=>"111111111",
126060=>"000011110",
126061=>"111111011",
126062=>"010000111",
126063=>"000100000",
126064=>"001000000",
126065=>"101101010",
126066=>"010011100",
126067=>"111101000",
126068=>"000111111",
126069=>"101101111",
126070=>"101001000",
126071=>"111011001",
126072=>"111000000",
126073=>"001010000",
126074=>"001000001",
126075=>"000111111",
126076=>"111000000",
126077=>"010100000",
126078=>"000001111",
126079=>"010010001",
126080=>"111111110",
126081=>"001001111",
126082=>"000100000",
126083=>"011010010",
126084=>"000010010",
126085=>"111001000",
126086=>"000110000",
126087=>"111001011",
126088=>"000001100",
126089=>"001111001",
126090=>"100000000",
126091=>"011000100",
126092=>"110010001",
126093=>"111111101",
126094=>"011111100",
126095=>"110100000",
126096=>"110100100",
126097=>"001001000",
126098=>"010001111",
126099=>"111000000",
126100=>"001010000",
126101=>"101000111",
126102=>"101101101",
126103=>"011000000",
126104=>"010000111",
126105=>"000000111",
126106=>"000001111",
126107=>"110111010",
126108=>"001001111",
126109=>"000111000",
126110=>"000001111",
126111=>"101101101",
126112=>"111110011",
126113=>"100101000",
126114=>"111010000",
126115=>"001000111",
126116=>"000111110",
126117=>"111001001",
126118=>"100000001",
126119=>"000111110",
126120=>"010111111",
126121=>"111000000",
126122=>"111101111",
126123=>"001000000",
126124=>"111010000",
126125=>"111010000",
126126=>"001000000",
126127=>"011010000",
126128=>"001100110",
126129=>"011011110",
126130=>"100100000",
126131=>"100000100",
126132=>"001001011",
126133=>"000000110",
126134=>"000110000",
126135=>"110000111",
126136=>"011010010",
126137=>"111000110",
126138=>"010000000",
126139=>"000100000",
126140=>"000000000",
126141=>"111111000",
126142=>"111011000",
126143=>"001101111",
126144=>"000000111",
126145=>"001010111",
126146=>"111111000",
126147=>"011100000",
126148=>"011010010",
126149=>"000010000",
126150=>"111101011",
126151=>"000000100",
126152=>"001000111",
126153=>"000000000",
126154=>"111100100",
126155=>"000101101",
126156=>"111111101",
126157=>"111000000",
126158=>"000000000",
126159=>"010100000",
126160=>"111010111",
126161=>"110110100",
126162=>"111111010",
126163=>"111101111",
126164=>"100000111",
126165=>"100111000",
126166=>"000000000",
126167=>"001111010",
126168=>"000000101",
126169=>"110010000",
126170=>"111111111",
126171=>"000100010",
126172=>"101001011",
126173=>"111111110",
126174=>"000010001",
126175=>"001101101",
126176=>"111010010",
126177=>"100010110",
126178=>"111011001",
126179=>"111111001",
126180=>"000000101",
126181=>"000010010",
126182=>"010010110",
126183=>"001011111",
126184=>"000000010",
126185=>"000000000",
126186=>"001101111",
126187=>"111100000",
126188=>"000010000",
126189=>"100001001",
126190=>"000000000",
126191=>"100000000",
126192=>"001000000",
126193=>"001010000",
126194=>"000001011",
126195=>"110100000",
126196=>"101000011",
126197=>"111111001",
126198=>"000000010",
126199=>"000000110",
126200=>"001000000",
126201=>"101111110",
126202=>"111110000",
126203=>"001010000",
126204=>"111111111",
126205=>"001000001",
126206=>"110001001",
126207=>"111101000",
126208=>"100011011",
126209=>"000100110",
126210=>"001000001",
126211=>"000000110",
126212=>"100110100",
126213=>"001001001",
126214=>"111110111",
126215=>"000110110",
126216=>"110000000",
126217=>"011001011",
126218=>"000100101",
126219=>"000000001",
126220=>"000000101",
126221=>"110110000",
126222=>"000010100",
126223=>"111111001",
126224=>"000100100",
126225=>"001100110",
126226=>"011001000",
126227=>"111100110",
126228=>"001001101",
126229=>"001001111",
126230=>"001011011",
126231=>"100110110",
126232=>"011001001",
126233=>"111111011",
126234=>"111111110",
126235=>"000111101",
126236=>"000111011",
126237=>"110110100",
126238=>"001011100",
126239=>"000010110",
126240=>"001001001",
126241=>"000001001",
126242=>"000000100",
126243=>"000000100",
126244=>"001001001",
126245=>"100100010",
126246=>"101100110",
126247=>"110110000",
126248=>"011010010",
126249=>"000000000",
126250=>"000110100",
126251=>"110000010",
126252=>"100101110",
126253=>"011011101",
126254=>"100001011",
126255=>"111011100",
126256=>"110011011",
126257=>"110111011",
126258=>"011111001",
126259=>"011001000",
126260=>"100110110",
126261=>"100100100",
126262=>"000000110",
126263=>"100110100",
126264=>"010011001",
126265=>"000000110",
126266=>"011001000",
126267=>"100100101",
126268=>"000100000",
126269=>"000111010",
126270=>"001001000",
126271=>"100010100",
126272=>"111001101",
126273=>"100100110",
126274=>"001111111",
126275=>"100110011",
126276=>"010001010",
126277=>"100000000",
126278=>"111111001",
126279=>"011011010",
126280=>"110011010",
126281=>"010011001",
126282=>"001100111",
126283=>"111100111",
126284=>"111001100",
126285=>"000011011",
126286=>"000001001",
126287=>"111010010",
126288=>"000000010",
126289=>"110111111",
126290=>"011011011",
126291=>"110011001",
126292=>"001001011",
126293=>"000111001",
126294=>"000001100",
126295=>"011000000",
126296=>"011111111",
126297=>"101011011",
126298=>"000000001",
126299=>"111111101",
126300=>"000010010",
126301=>"110011011",
126302=>"100110100",
126303=>"111100000",
126304=>"110000011",
126305=>"100000110",
126306=>"011001101",
126307=>"001111111",
126308=>"110010000",
126309=>"110110000",
126310=>"000000010",
126311=>"000110100",
126312=>"000001111",
126313=>"011011111",
126314=>"110000000",
126315=>"101001111",
126316=>"011001111",
126317=>"101100100",
126318=>"000000000",
126319=>"000011111",
126320=>"100011001",
126321=>"010110110",
126322=>"010000101",
126323=>"001000100",
126324=>"111111010",
126325=>"011001100",
126326=>"011000111",
126327=>"110000011",
126328=>"011111001",
126329=>"001111110",
126330=>"111111011",
126331=>"110011011",
126332=>"000100110",
126333=>"100000000",
126334=>"111110010",
126335=>"001000001",
126336=>"100000111",
126337=>"011001000",
126338=>"001001000",
126339=>"100000000",
126340=>"001110100",
126341=>"101001101",
126342=>"100101111",
126343=>"000000001",
126344=>"000000000",
126345=>"100110010",
126346=>"111011001",
126347=>"110001001",
126348=>"000100110",
126349=>"001001011",
126350=>"011111000",
126351=>"000000000",
126352=>"111011001",
126353=>"000100100",
126354=>"110110011",
126355=>"000110010",
126356=>"010100010",
126357=>"001001100",
126358=>"000100100",
126359=>"110100100",
126360=>"110010000",
126361=>"011011001",
126362=>"001011110",
126363=>"011011000",
126364=>"100110111",
126365=>"111001111",
126366=>"110110010",
126367=>"000100100",
126368=>"011011001",
126369=>"001101111",
126370=>"100011011",
126371=>"000011010",
126372=>"011011111",
126373=>"000000000",
126374=>"101001100",
126375=>"100100100",
126376=>"101001110",
126377=>"011001011",
126378=>"011001001",
126379=>"001000100",
126380=>"000001000",
126381=>"110010011",
126382=>"000100100",
126383=>"000011111",
126384=>"000000010",
126385=>"111110000",
126386=>"110011011",
126387=>"000001000",
126388=>"110111101",
126389=>"010101000",
126390=>"000101011",
126391=>"110010010",
126392=>"110101111",
126393=>"100100000",
126394=>"110010111",
126395=>"011011011",
126396=>"001110010",
126397=>"011101001",
126398=>"010000011",
126399=>"000100111",
126400=>"011001001",
126401=>"000000010",
126402=>"001101110",
126403=>"110011011",
126404=>"100010000",
126405=>"010011011",
126406=>"110111111",
126407=>"011101111",
126408=>"110010011",
126409=>"000100110",
126410=>"011001000",
126411=>"000100001",
126412=>"100110010",
126413=>"010000100",
126414=>"000100000",
126415=>"111101000",
126416=>"000100000",
126417=>"100010100",
126418=>"001100011",
126419=>"111111000",
126420=>"100101001",
126421=>"001000001",
126422=>"000010001",
126423=>"100101111",
126424=>"100110110",
126425=>"110100100",
126426=>"000001001",
126427=>"011001101",
126428=>"000010000",
126429=>"001101011",
126430=>"000101111",
126431=>"100011000",
126432=>"000100000",
126433=>"001001000",
126434=>"100110110",
126435=>"111001001",
126436=>"001000011",
126437=>"111011011",
126438=>"100110110",
126439=>"110111011",
126440=>"111111100",
126441=>"100110101",
126442=>"101110010",
126443=>"011001001",
126444=>"100100100",
126445=>"100110110",
126446=>"000000001",
126447=>"100010010",
126448=>"100110110",
126449=>"111011011",
126450=>"000111000",
126451=>"100010000",
126452=>"101101001",
126453=>"011000001",
126454=>"101000000",
126455=>"010110010",
126456=>"000100110",
126457=>"000110110",
126458=>"111001111",
126459=>"110111001",
126460=>"001111011",
126461=>"000001010",
126462=>"111001001",
126463=>"100110010",
126464=>"100000110",
126465=>"000000001",
126466=>"011000001",
126467=>"111111111",
126468=>"101101001",
126469=>"100001000",
126470=>"000111111",
126471=>"111001110",
126472=>"000000000",
126473=>"000000000",
126474=>"100100100",
126475=>"000000111",
126476=>"000000111",
126477=>"111010111",
126478=>"100000100",
126479=>"100000000",
126480=>"001001001",
126481=>"000000000",
126482=>"000000000",
126483=>"000000000",
126484=>"001000011",
126485=>"111001111",
126486=>"101001001",
126487=>"000000100",
126488=>"001000000",
126489=>"111111010",
126490=>"100001000",
126491=>"000001000",
126492=>"110101001",
126493=>"111101100",
126494=>"000001000",
126495=>"110010010",
126496=>"001001000",
126497=>"111101111",
126498=>"110011111",
126499=>"000001010",
126500=>"111111111",
126501=>"000000011",
126502=>"001100001",
126503=>"000001111",
126504=>"111101000",
126505=>"110100000",
126506=>"000000010",
126507=>"011010001",
126508=>"101000100",
126509=>"000000111",
126510=>"101101100",
126511=>"111011001",
126512=>"000000000",
126513=>"001000000",
126514=>"000111110",
126515=>"111110110",
126516=>"000100100",
126517=>"110101111",
126518=>"000000100",
126519=>"000111111",
126520=>"000000011",
126521=>"100100111",
126522=>"101100111",
126523=>"000100010",
126524=>"001001111",
126525=>"110010010",
126526=>"000001101",
126527=>"000100110",
126528=>"111100001",
126529=>"000000101",
126530=>"111101101",
126531=>"000000000",
126532=>"111011111",
126533=>"111100001",
126534=>"000110100",
126535=>"011100010",
126536=>"001001111",
126537=>"000000000",
126538=>"001000110",
126539=>"111111010",
126540=>"000000000",
126541=>"001001001",
126542=>"100101100",
126543=>"111111010",
126544=>"010110000",
126545=>"110000000",
126546=>"010001101",
126547=>"001000010",
126548=>"110100000",
126549=>"001010011",
126550=>"111111110",
126551=>"000010110",
126552=>"000000000",
126553=>"001000000",
126554=>"001001001",
126555=>"101100100",
126556=>"000000000",
126557=>"000000000",
126558=>"111111111",
126559=>"000000000",
126560=>"000010000",
126561=>"110010011",
126562=>"000001000",
126563=>"001000000",
126564=>"000000011",
126565=>"101111100",
126566=>"000011111",
126567=>"111110100",
126568=>"001101111",
126569=>"100001111",
126570=>"000000000",
126571=>"100001111",
126572=>"110110101",
126573=>"111100000",
126574=>"001000001",
126575=>"101000000",
126576=>"001001100",
126577=>"000000001",
126578=>"000000000",
126579=>"111000000",
126580=>"000000010",
126581=>"100000100",
126582=>"011001000",
126583=>"001111111",
126584=>"001000000",
126585=>"111000000",
126586=>"111111111",
126587=>"000010011",
126588=>"011001001",
126589=>"000001010",
126590=>"000001101",
126591=>"001001000",
126592=>"101000000",
126593=>"000000000",
126594=>"000000000",
126595=>"111110010",
126596=>"111001000",
126597=>"111011000",
126598=>"000000000",
126599=>"100100101",
126600=>"000001100",
126601=>"101000001",
126602=>"101111111",
126603=>"000000000",
126604=>"111111000",
126605=>"000000000",
126606=>"001101101",
126607=>"001001001",
126608=>"100100100",
126609=>"000000000",
126610=>"000000111",
126611=>"001001111",
126612=>"111000000",
126613=>"000000000",
126614=>"111001111",
126615=>"001100101",
126616=>"111001000",
126617=>"001101011",
126618=>"000000000",
126619=>"111111011",
126620=>"100111111",
126621=>"101101111",
126622=>"010110111",
126623=>"000000001",
126624=>"111111111",
126625=>"111101001",
126626=>"000000010",
126627=>"001111011",
126628=>"000000011",
126629=>"011011111",
126630=>"011000000",
126631=>"110000010",
126632=>"000000101",
126633=>"001001001",
126634=>"101101000",
126635=>"000001000",
126636=>"111001000",
126637=>"001111001",
126638=>"100100100",
126639=>"111111111",
126640=>"111111111",
126641=>"100110111",
126642=>"001010101",
126643=>"000000100",
126644=>"100000010",
126645=>"100111110",
126646=>"111110001",
126647=>"100111111",
126648=>"100101111",
126649=>"000000010",
126650=>"101111011",
126651=>"000000010",
126652=>"111111111",
126653=>"111110110",
126654=>"100110011",
126655=>"000001000",
126656=>"000000100",
126657=>"000101111",
126658=>"000000111",
126659=>"111111110",
126660=>"000000011",
126661=>"100000011",
126662=>"000000001",
126663=>"000000000",
126664=>"010010001",
126665=>"101101101",
126666=>"000001110",
126667=>"000111110",
126668=>"000101101",
126669=>"110100000",
126670=>"111111111",
126671=>"001110010",
126672=>"110000110",
126673=>"011111011",
126674=>"111101111",
126675=>"101000010",
126676=>"000000001",
126677=>"011111110",
126678=>"000001111",
126679=>"000010010",
126680=>"000000111",
126681=>"110100110",
126682=>"111111111",
126683=>"111110000",
126684=>"000001000",
126685=>"111111111",
126686=>"110110000",
126687=>"011110111",
126688=>"100000000",
126689=>"111111101",
126690=>"111111111",
126691=>"011010011",
126692=>"000100111",
126693=>"011111111",
126694=>"000000000",
126695=>"001011001",
126696=>"111000011",
126697=>"000000000",
126698=>"001001001",
126699=>"000101000",
126700=>"111101111",
126701=>"111110011",
126702=>"010000000",
126703=>"000000111",
126704=>"000000010",
126705=>"001001101",
126706=>"000000111",
126707=>"000000000",
126708=>"000110101",
126709=>"111011111",
126710=>"000000010",
126711=>"111000011",
126712=>"000000101",
126713=>"000010110",
126714=>"111110010",
126715=>"000000111",
126716=>"101101101",
126717=>"100111001",
126718=>"101000000",
126719=>"111101010",
126720=>"001010110",
126721=>"000111111",
126722=>"001100111",
126723=>"000111111",
126724=>"011001000",
126725=>"000000000",
126726=>"101111111",
126727=>"111010000",
126728=>"110001111",
126729=>"100000111",
126730=>"100111110",
126731=>"110000000",
126732=>"111110000",
126733=>"110010000",
126734=>"110110011",
126735=>"110000000",
126736=>"011001000",
126737=>"111000000",
126738=>"001101111",
126739=>"000001101",
126740=>"110111111",
126741=>"000000111",
126742=>"000100111",
126743=>"111010111",
126744=>"111111111",
126745=>"110011000",
126746=>"110110111",
126747=>"110000011",
126748=>"111111000",
126749=>"100111111",
126750=>"000101101",
126751=>"011111111",
126752=>"000000010",
126753=>"000000001",
126754=>"000001000",
126755=>"101111000",
126756=>"011000001",
126757=>"000000010",
126758=>"000001111",
126759=>"111000000",
126760=>"101111111",
126761=>"110010110",
126762=>"000010000",
126763=>"000101111",
126764=>"111000111",
126765=>"101110111",
126766=>"111001001",
126767=>"011010001",
126768=>"000010000",
126769=>"011011001",
126770=>"000111101",
126771=>"111111101",
126772=>"101110110",
126773=>"101110011",
126774=>"000001111",
126775=>"110101011",
126776=>"011100011",
126777=>"010000000",
126778=>"000111011",
126779=>"010011011",
126780=>"110000000",
126781=>"111110000",
126782=>"000001011",
126783=>"100100000",
126784=>"100100101",
126785=>"010110000",
126786=>"000101010",
126787=>"000000000",
126788=>"010000000",
126789=>"111110000",
126790=>"000000000",
126791=>"101101101",
126792=>"101111001",
126793=>"011111111",
126794=>"000000000",
126795=>"111111010",
126796=>"111100100",
126797=>"100001000",
126798=>"110100000",
126799=>"101111111",
126800=>"001000111",
126801=>"111110000",
126802=>"101000000",
126803=>"001001001",
126804=>"000011000",
126805=>"000111111",
126806=>"110110010",
126807=>"111001000",
126808=>"110001001",
126809=>"001011101",
126810=>"111111111",
126811=>"100000000",
126812=>"000100111",
126813=>"001000011",
126814=>"111111110",
126815=>"000000110",
126816=>"100111111",
126817=>"001011111",
126818=>"100000000",
126819=>"001100100",
126820=>"001001000",
126821=>"111101100",
126822=>"110111111",
126823=>"010001011",
126824=>"000111111",
126825=>"001001000",
126826=>"111000100",
126827=>"101100000",
126828=>"110100111",
126829=>"001000010",
126830=>"000100111",
126831=>"001111111",
126832=>"001000001",
126833=>"000110000",
126834=>"000100010",
126835=>"101011000",
126836=>"010000000",
126837=>"000000000",
126838=>"110110000",
126839=>"100010010",
126840=>"000110011",
126841=>"110100000",
126842=>"001000000",
126843=>"011010000",
126844=>"100000000",
126845=>"100000010",
126846=>"000000111",
126847=>"111111110",
126848=>"000000000",
126849=>"101101000",
126850=>"100000100",
126851=>"000111111",
126852=>"110000100",
126853=>"111010110",
126854=>"100000110",
126855=>"011000000",
126856=>"110110100",
126857=>"010001011",
126858=>"111011011",
126859=>"010000001",
126860=>"001001110",
126861=>"100000100",
126862=>"000000000",
126863=>"000010010",
126864=>"111101000",
126865=>"111000000",
126866=>"001001011",
126867=>"000110011",
126868=>"110000000",
126869=>"101001001",
126870=>"101101010",
126871=>"011010100",
126872=>"000000000",
126873=>"000001001",
126874=>"000100111",
126875=>"101000000",
126876=>"101011111",
126877=>"010000000",
126878=>"000011000",
126879=>"111110100",
126880=>"001011011",
126881=>"000000111",
126882=>"011010111",
126883=>"001001000",
126884=>"000001111",
126885=>"110000100",
126886=>"001111010",
126887=>"000101111",
126888=>"100100001",
126889=>"110110100",
126890=>"101101111",
126891=>"010000100",
126892=>"110111110",
126893=>"111000000",
126894=>"000010111",
126895=>"101100000",
126896=>"000000000",
126897=>"000000000",
126898=>"111000010",
126899=>"110000101",
126900=>"001011111",
126901=>"101111111",
126902=>"000000001",
126903=>"110011010",
126904=>"011100111",
126905=>"010111000",
126906=>"010000111",
126907=>"111011111",
126908=>"001000010",
126909=>"111000100",
126910=>"000000000",
126911=>"000011111",
126912=>"101101111",
126913=>"000000010",
126914=>"100000000",
126915=>"001011000",
126916=>"011011111",
126917=>"000100010",
126918=>"011011000",
126919=>"000101110",
126920=>"010000000",
126921=>"100100000",
126922=>"001110111",
126923=>"110000000",
126924=>"011111000",
126925=>"001010110",
126926=>"000000000",
126927=>"000100111",
126928=>"000110000",
126929=>"000110010",
126930=>"010011001",
126931=>"111000110",
126932=>"111000000",
126933=>"000111011",
126934=>"110110111",
126935=>"001101110",
126936=>"111011000",
126937=>"000100100",
126938=>"110101111",
126939=>"101111011",
126940=>"001100110",
126941=>"011010111",
126942=>"000100000",
126943=>"001000000",
126944=>"011101010",
126945=>"101001011",
126946=>"111110100",
126947=>"011111111",
126948=>"111001000",
126949=>"111000000",
126950=>"111100000",
126951=>"100000010",
126952=>"101000000",
126953=>"001000101",
126954=>"101111111",
126955=>"000101110",
126956=>"111110010",
126957=>"011111001",
126958=>"111000000",
126959=>"111100000",
126960=>"101111011",
126961=>"011011111",
126962=>"111000110",
126963=>"110100000",
126964=>"101000011",
126965=>"101010011",
126966=>"111000000",
126967=>"100000000",
126968=>"000000000",
126969=>"110110111",
126970=>"101000000",
126971=>"101001000",
126972=>"000000010",
126973=>"010000000",
126974=>"001000011",
126975=>"010000000",
126976=>"111011111",
126977=>"111110000",
126978=>"101000000",
126979=>"000110110",
126980=>"100110110",
126981=>"000100111",
126982=>"110111000",
126983=>"111011111",
126984=>"100110011",
126985=>"000000100",
126986=>"101000000",
126987=>"000000000",
126988=>"100001001",
126989=>"111110000",
126990=>"011000011",
126991=>"001000000",
126992=>"110111100",
126993=>"001000000",
126994=>"100001000",
126995=>"001111110",
126996=>"111101101",
126997=>"110110110",
126998=>"010000000",
126999=>"001011111",
127000=>"101001000",
127001=>"000000000",
127002=>"000000011",
127003=>"001111111",
127004=>"000000101",
127005=>"011001000",
127006=>"111111111",
127007=>"011000000",
127008=>"000000000",
127009=>"110101000",
127010=>"000000101",
127011=>"000000000",
127012=>"100111101",
127013=>"110111111",
127014=>"110010000",
127015=>"111111111",
127016=>"111001111",
127017=>"111111111",
127018=>"101111111",
127019=>"001000000",
127020=>"110100100",
127021=>"000110010",
127022=>"110110101",
127023=>"000101000",
127024=>"111111110",
127025=>"110100000",
127026=>"000010010",
127027=>"000110111",
127028=>"000000000",
127029=>"001001001",
127030=>"000000001",
127031=>"110111110",
127032=>"000111111",
127033=>"110110010",
127034=>"000101111",
127035=>"000000000",
127036=>"100001000",
127037=>"111111011",
127038=>"001000100",
127039=>"110111001",
127040=>"110011001",
127041=>"001001101",
127042=>"111111100",
127043=>"110110001",
127044=>"001111100",
127045=>"001101000",
127046=>"000111010",
127047=>"000111110",
127048=>"110111011",
127049=>"010000001",
127050=>"111001000",
127051=>"111111110",
127052=>"111111111",
127053=>"100011011",
127054=>"010011101",
127055=>"001001101",
127056=>"001100111",
127057=>"111111111",
127058=>"111111111",
127059=>"111101101",
127060=>"001001010",
127061=>"001111110",
127062=>"001011111",
127063=>"001000001",
127064=>"100100100",
127065=>"000100110",
127066=>"000101001",
127067=>"011011111",
127068=>"111111110",
127069=>"001001001",
127070=>"000110010",
127071=>"110110100",
127072=>"000000001",
127073=>"010110111",
127074=>"000000000",
127075=>"000011001",
127076=>"110111111",
127077=>"010100100",
127078=>"101001001",
127079=>"111111000",
127080=>"110010010",
127081=>"001000000",
127082=>"111111111",
127083=>"110001101",
127084=>"111000001",
127085=>"001001000",
127086=>"010111110",
127087=>"100101111",
127088=>"011111011",
127089=>"010101111",
127090=>"000100010",
127091=>"101001001",
127092=>"111110110",
127093=>"001000001",
127094=>"110111101",
127095=>"100001111",
127096=>"000000000",
127097=>"111001000",
127098=>"001011010",
127099=>"110111100",
127100=>"110100100",
127101=>"110100100",
127102=>"000101000",
127103=>"101110000",
127104=>"000001001",
127105=>"111111111",
127106=>"111010010",
127107=>"111111111",
127108=>"000111110",
127109=>"000111110",
127110=>"010000101",
127111=>"001001001",
127112=>"110110111",
127113=>"111000010",
127114=>"101101100",
127115=>"001101000",
127116=>"000000000",
127117=>"111101000",
127118=>"000110010",
127119=>"000001001",
127120=>"000001010",
127121=>"000100111",
127122=>"011010011",
127123=>"110101001",
127124=>"111010010",
127125=>"000000001",
127126=>"000000000",
127127=>"110011110",
127128=>"000000000",
127129=>"100001101",
127130=>"010111110",
127131=>"000000000",
127132=>"001111111",
127133=>"000001000",
127134=>"111111111",
127135=>"101001001",
127136=>"100000100",
127137=>"010001010",
127138=>"111111100",
127139=>"010011000",
127140=>"111111111",
127141=>"001001011",
127142=>"100110100",
127143=>"111011100",
127144=>"001100110",
127145=>"111111101",
127146=>"001001001",
127147=>"001000000",
127148=>"000111111",
127149=>"111110110",
127150=>"100101111",
127151=>"100101111",
127152=>"111111100",
127153=>"011011001",
127154=>"111011011",
127155=>"110100100",
127156=>"111101100",
127157=>"000000000",
127158=>"000000000",
127159=>"000000000",
127160=>"001000000",
127161=>"101100100",
127162=>"010010000",
127163=>"110000011",
127164=>"000001000",
127165=>"001010011",
127166=>"001111000",
127167=>"111011001",
127168=>"000110010",
127169=>"000000000",
127170=>"010110111",
127171=>"111011001",
127172=>"001000111",
127173=>"001100110",
127174=>"111110001",
127175=>"100110111",
127176=>"110010111",
127177=>"110110111",
127178=>"000000000",
127179=>"000010000",
127180=>"111010000",
127181=>"011001001",
127182=>"000000000",
127183=>"111000000",
127184=>"110111111",
127185=>"110101011",
127186=>"000000111",
127187=>"011101111",
127188=>"000000111",
127189=>"100001000",
127190=>"101110111",
127191=>"111101111",
127192=>"000000000",
127193=>"000000010",
127194=>"010000010",
127195=>"001001101",
127196=>"001100110",
127197=>"001001000",
127198=>"110100110",
127199=>"110111100",
127200=>"111110001",
127201=>"000100000",
127202=>"000000001",
127203=>"101001000",
127204=>"000000000",
127205=>"000001101",
127206=>"000100110",
127207=>"111011101",
127208=>"111001101",
127209=>"000001001",
127210=>"001000000",
127211=>"001000001",
127212=>"000000000",
127213=>"000111001",
127214=>"111000000",
127215=>"111000001",
127216=>"000000000",
127217=>"000011110",
127218=>"111111110",
127219=>"011011011",
127220=>"101100100",
127221=>"001000010",
127222=>"011000001",
127223=>"000111010",
127224=>"100111111",
127225=>"011111101",
127226=>"101111010",
127227=>"001001000",
127228=>"110110110",
127229=>"001000000",
127230=>"111100111",
127231=>"111000001",
127232=>"011001011",
127233=>"110111111",
127234=>"000001111",
127235=>"000000000",
127236=>"001000011",
127237=>"000111101",
127238=>"111000000",
127239=>"111111101",
127240=>"010010000",
127241=>"000000000",
127242=>"001000110",
127243=>"000011000",
127244=>"000100111",
127245=>"000000001",
127246=>"100011001",
127247=>"001000000",
127248=>"111111111",
127249=>"000000110",
127250=>"000001000",
127251=>"101111110",
127252=>"011000000",
127253=>"000000111",
127254=>"101011111",
127255=>"100111111",
127256=>"000010000",
127257=>"000001000",
127258=>"000101111",
127259=>"000000101",
127260=>"001000000",
127261=>"100101111",
127262=>"000000000",
127263=>"000101000",
127264=>"010101101",
127265=>"011111111",
127266=>"100101100",
127267=>"000000111",
127268=>"011001011",
127269=>"101111000",
127270=>"000101111",
127271=>"001000010",
127272=>"100111111",
127273=>"000111111",
127274=>"111000000",
127275=>"110110110",
127276=>"111011000",
127277=>"110010000",
127278=>"010110111",
127279=>"000000000",
127280=>"100111000",
127281=>"001000000",
127282=>"010000100",
127283=>"000111000",
127284=>"000111111",
127285=>"111111111",
127286=>"001111100",
127287=>"110010000",
127288=>"010000000",
127289=>"000100110",
127290=>"100100100",
127291=>"000000000",
127292=>"111110010",
127293=>"110110110",
127294=>"000000011",
127295=>"111110000",
127296=>"110011111",
127297=>"111111001",
127298=>"010010010",
127299=>"011000000",
127300=>"100110110",
127301=>"000000010",
127302=>"001001000",
127303=>"110100001",
127304=>"100010001",
127305=>"111000000",
127306=>"000000010",
127307=>"000010111",
127308=>"000001000",
127309=>"111000000",
127310=>"111000000",
127311=>"001000010",
127312=>"111101010",
127313=>"111010010",
127314=>"100111111",
127315=>"001001000",
127316=>"001111000",
127317=>"001010110",
127318=>"010100111",
127319=>"101101101",
127320=>"000011011",
127321=>"100110111",
127322=>"111110101",
127323=>"100100110",
127324=>"110000000",
127325=>"001011011",
127326=>"111110000",
127327=>"100001010",
127328=>"010000000",
127329=>"000000000",
127330=>"001101111",
127331=>"010010110",
127332=>"101000000",
127333=>"001001010",
127334=>"110111000",
127335=>"101111011",
127336=>"110110010",
127337=>"010000000",
127338=>"110111110",
127339=>"111010111",
127340=>"111111111",
127341=>"111101011",
127342=>"101000000",
127343=>"000010001",
127344=>"111000001",
127345=>"000000111",
127346=>"001110011",
127347=>"001001001",
127348=>"000000000",
127349=>"000101001",
127350=>"101001110",
127351=>"000000010",
127352=>"000001111",
127353=>"010000010",
127354=>"110011101",
127355=>"111000000",
127356=>"011111110",
127357=>"100000100",
127358=>"000000111",
127359=>"000000010",
127360=>"001001000",
127361=>"101001001",
127362=>"010010000",
127363=>"111000010",
127364=>"100110010",
127365=>"111000000",
127366=>"111111001",
127367=>"111000100",
127368=>"110110001",
127369=>"000111111",
127370=>"000001101",
127371=>"011000101",
127372=>"000000110",
127373=>"111110000",
127374=>"111010000",
127375=>"000000000",
127376=>"101111011",
127377=>"110010011",
127378=>"000110111",
127379=>"010001000",
127380=>"010111110",
127381=>"000000111",
127382=>"111000000",
127383=>"011011001",
127384=>"010011000",
127385=>"010110000",
127386=>"000010111",
127387=>"111000000",
127388=>"011010111",
127389=>"010010000",
127390=>"000001000",
127391=>"101101111",
127392=>"011001001",
127393=>"000111111",
127394=>"110000000",
127395=>"100101101",
127396=>"011001000",
127397=>"101000000",
127398=>"110000001",
127399=>"111000000",
127400=>"000000101",
127401=>"110110000",
127402=>"001101111",
127403=>"000000000",
127404=>"110000000",
127405=>"100111100",
127406=>"110110011",
127407=>"110001000",
127408=>"010001000",
127409=>"110000000",
127410=>"101001101",
127411=>"001000110",
127412=>"111011000",
127413=>"000000110",
127414=>"000000000",
127415=>"000011100",
127416=>"010101010",
127417=>"111011000",
127418=>"111010000",
127419=>"110000100",
127420=>"110001001",
127421=>"101111111",
127422=>"110000000",
127423=>"000000000",
127424=>"000101111",
127425=>"100111111",
127426=>"011111000",
127427=>"001011111",
127428=>"100000000",
127429=>"100101100",
127430=>"111111010",
127431=>"001111111",
127432=>"001000100",
127433=>"110111101",
127434=>"000101111",
127435=>"111011000",
127436=>"010010000",
127437=>"111100110",
127438=>"000001111",
127439=>"101000000",
127440=>"000101111",
127441=>"110110110",
127442=>"000000110",
127443=>"011000000",
127444=>"001011011",
127445=>"110110110",
127446=>"000010111",
127447=>"010110111",
127448=>"000001110",
127449=>"110111000",
127450=>"100100110",
127451=>"000000111",
127452=>"000100011",
127453=>"010000000",
127454=>"000000010",
127455=>"000000000",
127456=>"000101111",
127457=>"000100000",
127458=>"000001001",
127459=>"011011001",
127460=>"000111111",
127461=>"010111010",
127462=>"000000101",
127463=>"010000100",
127464=>"111011101",
127465=>"010111111",
127466=>"000100011",
127467=>"000100111",
127468=>"000000101",
127469=>"000111111",
127470=>"101000010",
127471=>"101100100",
127472=>"000000000",
127473=>"011011011",
127474=>"000001001",
127475=>"011011000",
127476=>"111010000",
127477=>"000111111",
127478=>"000110111",
127479=>"100000000",
127480=>"111111010",
127481=>"000101000",
127482=>"100110111",
127483=>"011111101",
127484=>"000000111",
127485=>"111010000",
127486=>"011011100",
127487=>"110101000",
127488=>"011000100",
127489=>"011000001",
127490=>"001001111",
127491=>"000010010",
127492=>"111111000",
127493=>"110110000",
127494=>"010000001",
127495=>"111111110",
127496=>"100110000",
127497=>"101001100",
127498=>"100000001",
127499=>"111000000",
127500=>"000001110",
127501=>"110110000",
127502=>"011001101",
127503=>"000000000",
127504=>"110110000",
127505=>"000001101",
127506=>"000111111",
127507=>"110110000",
127508=>"000001100",
127509=>"111111111",
127510=>"011111111",
127511=>"011111111",
127512=>"100110110",
127513=>"111111111",
127514=>"101000111",
127515=>"000101111",
127516=>"100100001",
127517=>"110101000",
127518=>"100001001",
127519=>"000111111",
127520=>"001001001",
127521=>"111110001",
127522=>"000000000",
127523=>"100110110",
127524=>"000001000",
127525=>"110100000",
127526=>"001000110",
127527=>"000110000",
127528=>"011111010",
127529=>"101110111",
127530=>"000001111",
127531=>"000000000",
127532=>"010011000",
127533=>"000010011",
127534=>"111000000",
127535=>"000110111",
127536=>"000111110",
127537=>"111111010",
127538=>"001001000",
127539=>"001111111",
127540=>"011001111",
127541=>"111101000",
127542=>"110100001",
127543=>"001001001",
127544=>"001000010",
127545=>"001001111",
127546=>"011111110",
127547=>"011111011",
127548=>"000110100",
127549=>"010111010",
127550=>"000000011",
127551=>"000010000",
127552=>"111111101",
127553=>"111111111",
127554=>"110000001",
127555=>"110111001",
127556=>"010000010",
127557=>"100100000",
127558=>"110111111",
127559=>"111111001",
127560=>"001110000",
127561=>"110001110",
127562=>"111001111",
127563=>"101001101",
127564=>"101000000",
127565=>"111111100",
127566=>"100110100",
127567=>"111011001",
127568=>"110110000",
127569=>"101001110",
127570=>"001000000",
127571=>"010010000",
127572=>"000000110",
127573=>"101110011",
127574=>"011011010",
127575=>"111001111",
127576=>"100100111",
127577=>"001011111",
127578=>"110100100",
127579=>"011101000",
127580=>"000001111",
127581=>"000000000",
127582=>"111110000",
127583=>"110110101",
127584=>"000010000",
127585=>"000010111",
127586=>"000000011",
127587=>"011000011",
127588=>"000000000",
127589=>"011111000",
127590=>"000101000",
127591=>"000101000",
127592=>"110111110",
127593=>"111000000",
127594=>"110110000",
127595=>"111011001",
127596=>"100110111",
127597=>"001001101",
127598=>"000001100",
127599=>"001111110",
127600=>"101001100",
127601=>"111001001",
127602=>"001111100",
127603=>"000001111",
127604=>"010000000",
127605=>"000001001",
127606=>"110000001",
127607=>"000110000",
127608=>"000010110",
127609=>"010000000",
127610=>"001000000",
127611=>"110110001",
127612=>"100000110",
127613=>"110111000",
127614=>"010100111",
127615=>"101110101",
127616=>"111001000",
127617=>"110000001",
127618=>"101000000",
127619=>"000011010",
127620=>"110110101",
127621=>"001001111",
127622=>"011011000",
127623=>"001001011",
127624=>"101001011",
127625=>"010110000",
127626=>"001001111",
127627=>"111110111",
127628=>"000000000",
127629=>"001001001",
127630=>"000000111",
127631=>"001001001",
127632=>"111111000",
127633=>"000100100",
127634=>"001000000",
127635=>"010111111",
127636=>"001111100",
127637=>"111001101",
127638=>"101101111",
127639=>"011010000",
127640=>"001111111",
127641=>"001110110",
127642=>"111101101",
127643=>"010000000",
127644=>"001001001",
127645=>"000000000",
127646=>"001111110",
127647=>"001000111",
127648=>"101011111",
127649=>"110110111",
127650=>"000000000",
127651=>"000011101",
127652=>"000111001",
127653=>"001000100",
127654=>"000000000",
127655=>"111000000",
127656=>"001001001",
127657=>"100000001",
127658=>"111111111",
127659=>"001000001",
127660=>"001111101",
127661=>"001000110",
127662=>"110100011",
127663=>"000000001",
127664=>"010111101",
127665=>"101011000",
127666=>"010010010",
127667=>"000000000",
127668=>"000110000",
127669=>"010010010",
127670=>"010111010",
127671=>"110000101",
127672=>"010011011",
127673=>"000100101",
127674=>"011001001",
127675=>"110010110",
127676=>"000001000",
127677=>"010010000",
127678=>"010110000",
127679=>"000000100",
127680=>"100000001",
127681=>"000001111",
127682=>"110101001",
127683=>"111010000",
127684=>"000001011",
127685=>"101000101",
127686=>"110000000",
127687=>"110000000",
127688=>"110110110",
127689=>"111011001",
127690=>"110110110",
127691=>"000111110",
127692=>"000111110",
127693=>"011000001",
127694=>"001000010",
127695=>"110111110",
127696=>"110010000",
127697=>"110101110",
127698=>"101111111",
127699=>"101101101",
127700=>"000000001",
127701=>"000000010",
127702=>"101000101",
127703=>"010001111",
127704=>"001101110",
127705=>"000000000",
127706=>"011110100",
127707=>"101101111",
127708=>"101101110",
127709=>"011110111",
127710=>"000001001",
127711=>"101001111",
127712=>"111111010",
127713=>"001000111",
127714=>"110111000",
127715=>"011111000",
127716=>"000000001",
127717=>"110010000",
127718=>"111000000",
127719=>"000001111",
127720=>"001000000",
127721=>"000000000",
127722=>"001001000",
127723=>"111111111",
127724=>"000000000",
127725=>"011100001",
127726=>"000000010",
127727=>"111010010",
127728=>"111101110",
127729=>"011001011",
127730=>"000100101",
127731=>"110110110",
127732=>"110000100",
127733=>"001000000",
127734=>"101000101",
127735=>"000011000",
127736=>"000111010",
127737=>"110110000",
127738=>"101001011",
127739=>"001011010",
127740=>"100101111",
127741=>"111111110",
127742=>"100100000",
127743=>"001000111",
127744=>"000000000",
127745=>"100000001",
127746=>"001000101",
127747=>"101001011",
127748=>"000111000",
127749=>"100101001",
127750=>"000111111",
127751=>"110111111",
127752=>"010011110",
127753=>"111001111",
127754=>"011011010",
127755=>"111111111",
127756=>"100000000",
127757=>"111111101",
127758=>"100110100",
127759=>"011011111",
127760=>"011101110",
127761=>"011001000",
127762=>"000000000",
127763=>"000011010",
127764=>"101111000",
127765=>"001000001",
127766=>"001000000",
127767=>"111111001",
127768=>"000000100",
127769=>"111000011",
127770=>"010000101",
127771=>"000111101",
127772=>"001000101",
127773=>"000000010",
127774=>"000000000",
127775=>"111111111",
127776=>"111100010",
127777=>"111111111",
127778=>"000000111",
127779=>"000001000",
127780=>"001111011",
127781=>"011000001",
127782=>"001101001",
127783=>"000010110",
127784=>"000001011",
127785=>"100101111",
127786=>"000000000",
127787=>"101101101",
127788=>"110001011",
127789=>"001010000",
127790=>"001000000",
127791=>"110110100",
127792=>"000111100",
127793=>"001000011",
127794=>"000111111",
127795=>"011001101",
127796=>"000111000",
127797=>"101001000",
127798=>"110110100",
127799=>"000000100",
127800=>"111111111",
127801=>"000000000",
127802=>"000000001",
127803=>"000000110",
127804=>"001000111",
127805=>"111110011",
127806=>"000001101",
127807=>"100100100",
127808=>"101001111",
127809=>"000000000",
127810=>"111111010",
127811=>"010000001",
127812=>"000000011",
127813=>"000000000",
127814=>"000011100",
127815=>"101111111",
127816=>"000010000",
127817=>"000110111",
127818=>"100000001",
127819=>"011111010",
127820=>"111111110",
127821=>"001101100",
127822=>"001111110",
127823=>"000000010",
127824=>"000000001",
127825=>"011110111",
127826=>"101101000",
127827=>"110011011",
127828=>"100100101",
127829=>"001001000",
127830=>"000010010",
127831=>"101001101",
127832=>"111001000",
127833=>"010111011",
127834=>"010000000",
127835=>"111110000",
127836=>"000000100",
127837=>"000000010",
127838=>"110010000",
127839=>"000000000",
127840=>"000010000",
127841=>"001000101",
127842=>"000000011",
127843=>"011000010",
127844=>"111111111",
127845=>"010011110",
127846=>"011111111",
127847=>"001000111",
127848=>"011111101",
127849=>"111111111",
127850=>"111000000",
127851=>"000000001",
127852=>"001100110",
127853=>"111111101",
127854=>"111000001",
127855=>"010111111",
127856=>"110011110",
127857=>"111111011",
127858=>"011011111",
127859=>"000000000",
127860=>"111010000",
127861=>"000000111",
127862=>"011110000",
127863=>"000000111",
127864=>"101000000",
127865=>"011111100",
127866=>"111111111",
127867=>"001110110",
127868=>"011001011",
127869=>"001001000",
127870=>"010101111",
127871=>"000000010",
127872=>"000000001",
127873=>"101100111",
127874=>"000000000",
127875=>"000000010",
127876=>"011001001",
127877=>"111101011",
127878=>"100000100",
127879=>"111111111",
127880=>"000010010",
127881=>"010111000",
127882=>"011111000",
127883=>"001000101",
127884=>"111100000",
127885=>"000000000",
127886=>"111000000",
127887=>"000000111",
127888=>"111011011",
127889=>"000000000",
127890=>"111111000",
127891=>"000000011",
127892=>"111111101",
127893=>"101001001",
127894=>"111111100",
127895=>"110100001",
127896=>"000000001",
127897=>"000011001",
127898=>"101000101",
127899=>"100111101",
127900=>"100110100",
127901=>"010000010",
127902=>"101111111",
127903=>"100000111",
127904=>"000000000",
127905=>"111101000",
127906=>"101111111",
127907=>"000010000",
127908=>"001111101",
127909=>"010111111",
127910=>"000000010",
127911=>"101101111",
127912=>"101001001",
127913=>"111101001",
127914=>"111100101",
127915=>"101000000",
127916=>"110010000",
127917=>"000011001",
127918=>"011111111",
127919=>"010100111",
127920=>"001000101",
127921=>"100100111",
127922=>"101111001",
127923=>"001011111",
127924=>"110010110",
127925=>"010000000",
127926=>"000000000",
127927=>"111000011",
127928=>"000000011",
127929=>"111111111",
127930=>"000100111",
127931=>"010011111",
127932=>"100000000",
127933=>"101011000",
127934=>"001010010",
127935=>"000101100",
127936=>"000000000",
127937=>"001000000",
127938=>"111111010",
127939=>"000100000",
127940=>"000111001",
127941=>"111111111",
127942=>"110011111",
127943=>"111111111",
127944=>"000000010",
127945=>"101101000",
127946=>"000011000",
127947=>"100010000",
127948=>"000111100",
127949=>"100100110",
127950=>"111101111",
127951=>"010000100",
127952=>"111011100",
127953=>"000010100",
127954=>"111111111",
127955=>"111111010",
127956=>"111001101",
127957=>"001001000",
127958=>"101100000",
127959=>"110111101",
127960=>"000001001",
127961=>"000101010",
127962=>"001011011",
127963=>"101101001",
127964=>"100000110",
127965=>"110011101",
127966=>"110101010",
127967=>"000101110",
127968=>"000000000",
127969=>"111110000",
127970=>"110010000",
127971=>"000011011",
127972=>"000000000",
127973=>"000010111",
127974=>"101111100",
127975=>"100010011",
127976=>"110001100",
127977=>"111110100",
127978=>"100100000",
127979=>"000000001",
127980=>"001000111",
127981=>"101101001",
127982=>"111011011",
127983=>"000000001",
127984=>"011001001",
127985=>"111111111",
127986=>"000000101",
127987=>"011111010",
127988=>"000000111",
127989=>"010010010",
127990=>"000000111",
127991=>"000000000",
127992=>"100000101",
127993=>"111111000",
127994=>"111101000",
127995=>"111111111",
127996=>"011111011",
127997=>"000010000",
127998=>"000000000",
127999=>"000000000",
128000=>"010100110",
128001=>"010111111",
128002=>"101000100",
128003=>"010000000",
128004=>"111011011",
128005=>"011000000",
128006=>"111111011",
128007=>"000111011",
128008=>"000000100",
128009=>"000101001",
128010=>"111101101",
128011=>"111100000",
128012=>"100111111",
128013=>"111111000",
128014=>"111101100",
128015=>"000010000",
128016=>"010000000",
128017=>"101000100",
128018=>"000101000",
128019=>"110100000",
128020=>"000011111",
128021=>"000100110",
128022=>"000101101",
128023=>"101101101",
128024=>"111000100",
128025=>"110010000",
128026=>"010100000",
128027=>"111000000",
128028=>"111101001",
128029=>"000100111",
128030=>"110000000",
128031=>"000110111",
128032=>"011101000",
128033=>"111111011",
128034=>"000100111",
128035=>"000110000",
128036=>"011000001",
128037=>"011001010",
128038=>"000000001",
128039=>"111011000",
128040=>"111111001",
128041=>"100111010",
128042=>"000001000",
128043=>"110000000",
128044=>"111110100",
128045=>"101010101",
128046=>"000000000",
128047=>"101111101",
128048=>"000001111",
128049=>"111100000",
128050=>"000111111",
128051=>"011000111",
128052=>"111001000",
128053=>"111111101",
128054=>"110000000",
128055=>"000110111",
128056=>"100010001",
128057=>"000000000",
128058=>"011100101",
128059=>"000100001",
128060=>"110000000",
128061=>"000111111",
128062=>"100000000",
128063=>"111111111",
128064=>"100101100",
128065=>"110000011",
128066=>"010010010",
128067=>"011100000",
128068=>"000000000",
128069=>"000011100",
128070=>"111000000",
128071=>"001000101",
128072=>"000101111",
128073=>"011000000",
128074=>"001000111",
128075=>"000000000",
128076=>"111000000",
128077=>"000001100",
128078=>"110111100",
128079=>"111110101",
128080=>"101101000",
128081=>"111100000",
128082=>"010101100",
128083=>"010011001",
128084=>"101101100",
128085=>"001110111",
128086=>"001001000",
128087=>"111000000",
128088=>"111111000",
128089=>"111101100",
128090=>"111111101",
128091=>"001011011",
128092=>"000000010",
128093=>"000001001",
128094=>"000111111",
128095=>"000000000",
128096=>"011111110",
128097=>"001111110",
128098=>"111100000",
128099=>"100101111",
128100=>"100001010",
128101=>"010000000",
128102=>"111000000",
128103=>"000000011",
128104=>"111100110",
128105=>"000000000",
128106=>"101000010",
128107=>"000111101",
128108=>"000000111",
128109=>"101000000",
128110=>"000000000",
128111=>"001000011",
128112=>"000000011",
128113=>"001000001",
128114=>"011000000",
128115=>"000000000",
128116=>"011011001",
128117=>"000000000",
128118=>"111111101",
128119=>"000010011",
128120=>"111101000",
128121=>"110010111",
128122=>"000100000",
128123=>"001100111",
128124=>"111100000",
128125=>"000010000",
128126=>"000011011",
128127=>"101101100",
128128=>"100000000",
128129=>"000111010",
128130=>"000000011",
128131=>"000001010",
128132=>"111100000",
128133=>"000100010",
128134=>"010001011",
128135=>"000001001",
128136=>"111111110",
128137=>"011000000",
128138=>"000000011",
128139=>"000010000",
128140=>"000010010",
128141=>"000000110",
128142=>"100010111",
128143=>"110000000",
128144=>"100001001",
128145=>"110110111",
128146=>"101101100",
128147=>"100101000",
128148=>"100110100",
128149=>"111000000",
128150=>"110000000",
128151=>"000000011",
128152=>"000000000",
128153=>"000100011",
128154=>"111100000",
128155=>"011000000",
128156=>"011000111",
128157=>"111100000",
128158=>"001111111",
128159=>"000001111",
128160=>"001001011",
128161=>"101000011",
128162=>"000011111",
128163=>"000100111",
128164=>"011011000",
128165=>"010111111",
128166=>"001010011",
128167=>"010101001",
128168=>"111000100",
128169=>"000010011",
128170=>"111111100",
128171=>"111000000",
128172=>"000010011",
128173=>"111100000",
128174=>"110000001",
128175=>"000111111",
128176=>"000000100",
128177=>"000100011",
128178=>"111100100",
128179=>"000100000",
128180=>"010011011",
128181=>"111011111",
128182=>"000111010",
128183=>"111001000",
128184=>"011011000",
128185=>"000100011",
128186=>"111000101",
128187=>"111111111",
128188=>"011011010",
128189=>"111010000",
128190=>"000011110",
128191=>"000010011",
128192=>"101100100",
128193=>"101100100",
128194=>"111101111",
128195=>"000100000",
128196=>"000000000",
128197=>"111100101",
128198=>"000000011",
128199=>"111100100",
128200=>"111111000",
128201=>"100011000",
128202=>"110111001",
128203=>"000011010",
128204=>"011000110",
128205=>"110111001",
128206=>"111101101",
128207=>"011111111",
128208=>"011000100",
128209=>"010000100",
128210=>"010000000",
128211=>"001010111",
128212=>"101100101",
128213=>"000100111",
128214=>"111100000",
128215=>"001000000",
128216=>"000111011",
128217=>"000100111",
128218=>"100111111",
128219=>"100100000",
128220=>"110011001",
128221=>"111011101",
128222=>"000111111",
128223=>"011000000",
128224=>"111111000",
128225=>"000000100",
128226=>"101000111",
128227=>"011001011",
128228=>"001000000",
128229=>"000110010",
128230=>"101101000",
128231=>"000110100",
128232=>"000000000",
128233=>"011000000",
128234=>"111110101",
128235=>"011011000",
128236=>"000111000",
128237=>"111000000",
128238=>"000001001",
128239=>"010101101",
128240=>"011111101",
128241=>"101001011",
128242=>"011011000",
128243=>"001111101",
128244=>"010001001",
128245=>"011101000",
128246=>"010000100",
128247=>"001001000",
128248=>"111101000",
128249=>"000101100",
128250=>"000011000",
128251=>"000111001",
128252=>"011000000",
128253=>"101000001",
128254=>"000110111",
128255=>"111100011",
128256=>"001001001",
128257=>"101111111",
128258=>"100101111",
128259=>"001111111",
128260=>"111110011",
128261=>"000000001",
128262=>"100100110",
128263=>"111111101",
128264=>"000000110",
128265=>"000000000",
128266=>"111011000",
128267=>"101101000",
128268=>"101011110",
128269=>"000000000",
128270=>"110100100",
128271=>"111110000",
128272=>"101000111",
128273=>"111011111",
128274=>"001110111",
128275=>"111011000",
128276=>"000111110",
128277=>"101111111",
128278=>"001001111",
128279=>"010111101",
128280=>"000000000",
128281=>"101001111",
128282=>"000000000",
128283=>"000000100",
128284=>"101101000",
128285=>"011011111",
128286=>"111000000",
128287=>"000001111",
128288=>"110000101",
128289=>"000000001",
128290=>"000111001",
128291=>"000000111",
128292=>"000000000",
128293=>"110011001",
128294=>"110011010",
128295=>"000001101",
128296=>"101111000",
128297=>"010111000",
128298=>"111101101",
128299=>"000000011",
128300=>"111111010",
128301=>"001111111",
128302=>"000000011",
128303=>"110100111",
128304=>"111001000",
128305=>"000111110",
128306=>"000111101",
128307=>"000000000",
128308=>"111111101",
128309=>"101000000",
128310=>"110110110",
128311=>"010000001",
128312=>"000111111",
128313=>"000001000",
128314=>"101111111",
128315=>"000111001",
128316=>"111001001",
128317=>"000011000",
128318=>"000000111",
128319=>"010111001",
128320=>"000000000",
128321=>"111111110",
128322=>"110111000",
128323=>"010001001",
128324=>"000000000",
128325=>"000001000",
128326=>"111111000",
128327=>"101000110",
128328=>"111011001",
128329=>"001000001",
128330=>"000101011",
128331=>"110000000",
128332=>"010110111",
128333=>"001000010",
128334=>"111111110",
128335=>"101110111",
128336=>"111110111",
128337=>"011111100",
128338=>"111000111",
128339=>"000100111",
128340=>"000000010",
128341=>"100111110",
128342=>"011111100",
128343=>"000000000",
128344=>"000000111",
128345=>"100110111",
128346=>"111000000",
128347=>"111000000",
128348=>"001000000",
128349=>"001000111",
128350=>"011010010",
128351=>"010100100",
128352=>"111111000",
128353=>"100001000",
128354=>"000000011",
128355=>"011110110",
128356=>"011010001",
128357=>"000101101",
128358=>"000000111",
128359=>"000010110",
128360=>"000101000",
128361=>"011000101",
128362=>"111110000",
128363=>"000000000",
128364=>"001000100",
128365=>"110000111",
128366=>"110000000",
128367=>"111001000",
128368=>"011011001",
128369=>"001100101",
128370=>"111011001",
128371=>"001000100",
128372=>"011111110",
128373=>"000111111",
128374=>"111111000",
128375=>"011000000",
128376=>"101001110",
128377=>"000000111",
128378=>"000000000",
128379=>"000111111",
128380=>"000010011",
128381=>"100000000",
128382=>"010001111",
128383=>"000000011",
128384=>"000000000",
128385=>"011011000",
128386=>"010010111",
128387=>"010001110",
128388=>"001100111",
128389=>"000000000",
128390=>"001110000",
128391=>"110000000",
128392=>"111101000",
128393=>"000000011",
128394=>"000000111",
128395=>"000001111",
128396=>"000000001",
128397=>"010111101",
128398=>"111111111",
128399=>"000000011",
128400=>"100100110",
128401=>"000001000",
128402=>"010111001",
128403=>"000001000",
128404=>"000001001",
128405=>"111001101",
128406=>"111010000",
128407=>"011011010",
128408=>"111101000",
128409=>"000111000",
128410=>"111011010",
128411=>"000111100",
128412=>"011111000",
128413=>"000000000",
128414=>"110101100",
128415=>"000010110",
128416=>"101111000",
128417=>"100110111",
128418=>"011000000",
128419=>"001001101",
128420=>"001011011",
128421=>"001000001",
128422=>"111111101",
128423=>"010010001",
128424=>"000111111",
128425=>"111111111",
128426=>"101000111",
128427=>"000000110",
128428=>"111010000",
128429=>"001101111",
128430=>"000000111",
128431=>"000000001",
128432=>"111101101",
128433=>"011001000",
128434=>"010100111",
128435=>"100010011",
128436=>"111100110",
128437=>"111001101",
128438=>"011000001",
128439=>"001000111",
128440=>"110100100",
128441=>"011100100",
128442=>"111111110",
128443=>"001101001",
128444=>"111000011",
128445=>"010011000",
128446=>"100100100",
128447=>"001000001",
128448=>"000000110",
128449=>"100000000",
128450=>"010111100",
128451=>"001001000",
128452=>"000000111",
128453=>"110001111",
128454=>"100101111",
128455=>"010111111",
128456=>"111111000",
128457=>"000000100",
128458=>"111011111",
128459=>"111111001",
128460=>"010100101",
128461=>"011010100",
128462=>"111000110",
128463=>"000111110",
128464=>"000010000",
128465=>"111110010",
128466=>"101101101",
128467=>"111101100",
128468=>"111001111",
128469=>"100110000",
128470=>"000101111",
128471=>"110111000",
128472=>"001111001",
128473=>"101000111",
128474=>"101100000",
128475=>"000000101",
128476=>"001110111",
128477=>"000010111",
128478=>"001001111",
128479=>"001011111",
128480=>"000000000",
128481=>"001000010",
128482=>"101111111",
128483=>"111011000",
128484=>"001101001",
128485=>"001000001",
128486=>"111110000",
128487=>"000010110",
128488=>"011110100",
128489=>"000111011",
128490=>"111111000",
128491=>"111000000",
128492=>"000000000",
128493=>"000000111",
128494=>"000010000",
128495=>"111100010",
128496=>"111111000",
128497=>"010001011",
128498=>"110101111",
128499=>"111111111",
128500=>"101101111",
128501=>"000000100",
128502=>"000000101",
128503=>"000110100",
128504=>"111101001",
128505=>"111111101",
128506=>"100000000",
128507=>"110101111",
128508=>"110110000",
128509=>"111000000",
128510=>"001111100",
128511=>"110111000",
128512=>"110110110",
128513=>"101101010",
128514=>"000000000",
128515=>"111010100",
128516=>"111100001",
128517=>"111111000",
128518=>"011111011",
128519=>"010001100",
128520=>"111111100",
128521=>"001000000",
128522=>"000001111",
128523=>"101101000",
128524=>"100100101",
128525=>"000000010",
128526=>"011010110",
128527=>"111101000",
128528=>"011111000",
128529=>"000011011",
128530=>"101101110",
128531=>"010000100",
128532=>"111111111",
128533=>"101001001",
128534=>"011111011",
128535=>"110000010",
128536=>"111000101",
128537=>"001000101",
128538=>"100000011",
128539=>"101011010",
128540=>"000110000",
128541=>"111110000",
128542=>"100000101",
128543=>"100000100",
128544=>"011011000",
128545=>"111100000",
128546=>"111000101",
128547=>"011111111",
128548=>"000001101",
128549=>"100101010",
128550=>"111100100",
128551=>"000000111",
128552=>"111111000",
128553=>"100100111",
128554=>"101101010",
128555=>"110000000",
128556=>"001111111",
128557=>"010111111",
128558=>"011001100",
128559=>"000010010",
128560=>"100111101",
128561=>"111111011",
128562=>"000000111",
128563=>"111011111",
128564=>"011000000",
128565=>"100111011",
128566=>"010000000",
128567=>"000000100",
128568=>"001000000",
128569=>"100101101",
128570=>"111110100",
128571=>"101100110",
128572=>"100001101",
128573=>"100111010",
128574=>"001000000",
128575=>"100110111",
128576=>"011000000",
128577=>"010000111",
128578=>"000111101",
128579=>"011011110",
128580=>"100100100",
128581=>"100111000",
128582=>"010010000",
128583=>"010101011",
128584=>"111101001",
128585=>"011010000",
128586=>"111100000",
128587=>"000100000",
128588=>"100100000",
128589=>"000100100",
128590=>"011011110",
128591=>"010101111",
128592=>"000100001",
128593=>"010011010",
128594=>"011101010",
128595=>"011100101",
128596=>"111100000",
128597=>"100111100",
128598=>"010000100",
128599=>"111111011",
128600=>"111101111",
128601=>"111111111",
128602=>"011011111",
128603=>"010000101",
128604=>"000010000",
128605=>"101101001",
128606=>"100100111",
128607=>"110110001",
128608=>"000011110",
128609=>"000000000",
128610=>"111000101",
128611=>"111110100",
128612=>"000010000",
128613=>"011011101",
128614=>"110110001",
128615=>"011011000",
128616=>"001011110",
128617=>"100100000",
128618=>"000000011",
128619=>"111111111",
128620=>"111100110",
128621=>"000011111",
128622=>"001000000",
128623=>"100000000",
128624=>"111110000",
128625=>"100000111",
128626=>"011010110",
128627=>"000011101",
128628=>"000000110",
128629=>"000000000",
128630=>"100000000",
128631=>"000101111",
128632=>"000100111",
128633=>"001100101",
128634=>"101001000",
128635=>"100010111",
128636=>"010110001",
128637=>"010010000",
128638=>"010010010",
128639=>"111011010",
128640=>"000010111",
128641=>"010000000",
128642=>"011010000",
128643=>"111011101",
128644=>"010000001",
128645=>"110000111",
128646=>"011001011",
128647=>"100000001",
128648=>"001011000",
128649=>"000000000",
128650=>"011011011",
128651=>"111101111",
128652=>"000011000",
128653=>"100100001",
128654=>"111111110",
128655=>"110100000",
128656=>"110011001",
128657=>"110110111",
128658=>"111001010",
128659=>"111011000",
128660=>"111101011",
128661=>"101111000",
128662=>"000101000",
128663=>"101100000",
128664=>"001101001",
128665=>"100000111",
128666=>"001111111",
128667=>"000000000",
128668=>"000000100",
128669=>"100000000",
128670=>"000000110",
128671=>"111111000",
128672=>"110011001",
128673=>"111011100",
128674=>"111101111",
128675=>"000000111",
128676=>"000000111",
128677=>"011011110",
128678=>"111001001",
128679=>"000100000",
128680=>"100111111",
128681=>"000101100",
128682=>"111111111",
128683=>"111111010",
128684=>"001000000",
128685=>"000000000",
128686=>"110110010",
128687=>"000000000",
128688=>"000000000",
128689=>"001100110",
128690=>"000000000",
128691=>"000110100",
128692=>"111111111",
128693=>"000011111",
128694=>"000011000",
128695=>"101100111",
128696=>"100110101",
128697=>"011101100",
128698=>"010101100",
128699=>"001111111",
128700=>"111011011",
128701=>"111111011",
128702=>"010011001",
128703=>"100010011",
128704=>"000000000",
128705=>"111110010",
128706=>"111000011",
128707=>"111100011",
128708=>"000000111",
128709=>"111111101",
128710=>"000000000",
128711=>"000000110",
128712=>"100111000",
128713=>"000001100",
128714=>"000000010",
128715=>"111101000",
128716=>"000011011",
128717=>"010011111",
128718=>"011011011",
128719=>"000000010",
128720=>"010010000",
128721=>"010011011",
128722=>"111111000",
128723=>"111100000",
128724=>"000000100",
128725=>"001011101",
128726=>"011111111",
128727=>"010000000",
128728=>"000000100",
128729=>"000000000",
128730=>"000001000",
128731=>"101000101",
128732=>"011010000",
128733=>"000000101",
128734=>"000000000",
128735=>"000010000",
128736=>"000000000",
128737=>"100100111",
128738=>"101101001",
128739=>"110111100",
128740=>"000111000",
128741=>"111111111",
128742=>"100000000",
128743=>"011111101",
128744=>"100111101",
128745=>"100000000",
128746=>"100110010",
128747=>"011011111",
128748=>"011111111",
128749=>"100000101",
128750=>"000000000",
128751=>"000000100",
128752=>"000010000",
128753=>"111111011",
128754=>"000000000",
128755=>"011011011",
128756=>"000111000",
128757=>"111111000",
128758=>"000100000",
128759=>"000000001",
128760=>"000000000",
128761=>"110000000",
128762=>"010111111",
128763=>"011011000",
128764=>"000101000",
128765=>"111010100",
128766=>"000001111",
128767=>"000100100",
128768=>"100110011",
128769=>"011000010",
128770=>"100101111",
128771=>"111010010",
128772=>"001001101",
128773=>"110000001",
128774=>"001011101",
128775=>"000011111",
128776=>"100110010",
128777=>"001001000",
128778=>"100100000",
128779=>"100100100",
128780=>"100100110",
128781=>"111110000",
128782=>"001101101",
128783=>"000010010",
128784=>"110111001",
128785=>"001111001",
128786=>"100000000",
128787=>"000000011",
128788=>"011001010",
128789=>"111110110",
128790=>"001010000",
128791=>"000111110",
128792=>"011000000",
128793=>"001001001",
128794=>"000011000",
128795=>"001011111",
128796=>"100101101",
128797=>"011010000",
128798=>"100000101",
128799=>"100110110",
128800=>"111000111",
128801=>"110110100",
128802=>"000010100",
128803=>"000100100",
128804=>"011111111",
128805=>"111110010",
128806=>"011000001",
128807=>"000111011",
128808=>"001011010",
128809=>"010000111",
128810=>"000010110",
128811=>"101100000",
128812=>"111100010",
128813=>"011000000",
128814=>"001100111",
128815=>"100010000",
128816=>"011000001",
128817=>"101100100",
128818=>"000011011",
128819=>"001011011",
128820=>"110100000",
128821=>"011010000",
128822=>"000010110",
128823=>"000011111",
128824=>"110100100",
128825=>"011011111",
128826=>"001001100",
128827=>"011111111",
128828=>"100000001",
128829=>"010110100",
128830=>"100100000",
128831=>"011110010",
128832=>"100100111",
128833=>"111100011",
128834=>"101111111",
128835=>"100100111",
128836=>"111100000",
128837=>"000000111",
128838=>"000001011",
128839=>"011111111",
128840=>"100110110",
128841=>"000010000",
128842=>"110100111",
128843=>"100100110",
128844=>"100100110",
128845=>"111111101",
128846=>"100110110",
128847=>"111111011",
128848=>"100000111",
128849=>"110100000",
128850=>"011011111",
128851=>"001000000",
128852=>"011101110",
128853=>"110000110",
128854=>"100001101",
128855=>"001001101",
128856=>"111000000",
128857=>"001000000",
128858=>"000000110",
128859=>"001111111",
128860=>"000000001",
128861=>"000000000",
128862=>"111111111",
128863=>"000000101",
128864=>"000000000",
128865=>"111000000",
128866=>"100100110",
128867=>"111111111",
128868=>"110010010",
128869=>"011101100",
128870=>"011010011",
128871=>"011000011",
128872=>"001100111",
128873=>"001011011",
128874=>"000011011",
128875=>"100100000",
128876=>"000000111",
128877=>"011011000",
128878=>"000001001",
128879=>"000011011",
128880=>"011011100",
128881=>"001111101",
128882=>"100110001",
128883=>"011111000",
128884=>"001011010",
128885=>"100100000",
128886=>"100011101",
128887=>"110100111",
128888=>"100100110",
128889=>"000011111",
128890=>"001111110",
128891=>"011110110",
128892=>"100001001",
128893=>"110100100",
128894=>"100100100",
128895=>"100100100",
128896=>"100100010",
128897=>"110100110",
128898=>"000001011",
128899=>"001010000",
128900=>"000111011",
128901=>"010000000",
128902=>"101001011",
128903=>"100100100",
128904=>"011101011",
128905=>"011011010",
128906=>"001001000",
128907=>"000001111",
128908=>"100111000",
128909=>"101111000",
128910=>"011100100",
128911=>"001011000",
128912=>"001011000",
128913=>"110110000",
128914=>"100110000",
128915=>"110110001",
128916=>"010010000",
128917=>"100100111",
128918=>"000001000",
128919=>"111110110",
128920=>"000100100",
128921=>"110110100",
128922=>"110100100",
128923=>"000101111",
128924=>"011111101",
128925=>"100110111",
128926=>"000000110",
128927=>"100000000",
128928=>"001000100",
128929=>"111101011",
128930=>"100000110",
128931=>"100000001",
128932=>"000000111",
128933=>"111001011",
128934=>"010010000",
128935=>"000000011",
128936=>"001011011",
128937=>"000000000",
128938=>"110110111",
128939=>"100100100",
128940=>"110100000",
128941=>"110100001",
128942=>"110000111",
128943=>"000001000",
128944=>"100000011",
128945=>"000001001",
128946=>"110100100",
128947=>"100100001",
128948=>"001010000",
128949=>"011101100",
128950=>"000001001",
128951=>"010111001",
128952=>"110110110",
128953=>"101111000",
128954=>"111111000",
128955=>"100100110",
128956=>"011011001",
128957=>"100100110",
128958=>"001001111",
128959=>"001011001",
128960=>"111110111",
128961=>"000001001",
128962=>"001111011",
128963=>"101111010",
128964=>"011011100",
128965=>"100110111",
128966=>"111011000",
128967=>"110100010",
128968=>"000001001",
128969=>"100110110",
128970=>"011011001",
128971=>"001111101",
128972=>"011011010",
128973=>"010110110",
128974=>"100110111",
128975=>"100110110",
128976=>"001111111",
128977=>"110110000",
128978=>"000001001",
128979=>"011000000",
128980=>"110100111",
128981=>"000000010",
128982=>"100101111",
128983=>"000000001",
128984=>"000110111",
128985=>"000010000",
128986=>"111110100",
128987=>"001011001",
128988=>"100100111",
128989=>"111011000",
128990=>"010011011",
128991=>"110111001",
128992=>"100110110",
128993=>"101000111",
128994=>"000000110",
128995=>"111101011",
128996=>"011011000",
128997=>"100000011",
128998=>"011011011",
128999=>"001001111",
129000=>"001000111",
129001=>"011000010",
129002=>"000001001",
129003=>"000001001",
129004=>"110110111",
129005=>"011010000",
129006=>"100000000",
129007=>"100001000",
129008=>"001111111",
129009=>"000001110",
129010=>"000011111",
129011=>"111100000",
129012=>"011000010",
129013=>"000011010",
129014=>"001100001",
129015=>"011100101",
129016=>"100100110",
129017=>"010000011",
129018=>"111111101",
129019=>"011011010",
129020=>"011000000",
129021=>"000000001",
129022=>"011111111",
129023=>"111101101",
129024=>"100110110",
129025=>"000010000",
129026=>"011000000",
129027=>"001100100",
129028=>"000000001",
129029=>"000010001",
129030=>"111001110",
129031=>"000000000",
129032=>"000000000",
129033=>"000100111",
129034=>"100111111",
129035=>"000010111",
129036=>"011111011",
129037=>"101000111",
129038=>"011110110",
129039=>"101010000",
129040=>"000011111",
129041=>"111110110",
129042=>"111011011",
129043=>"000000001",
129044=>"001100111",
129045=>"000011000",
129046=>"111111001",
129047=>"101101101",
129048=>"000000101",
129049=>"000000001",
129050=>"000111111",
129051=>"111100100",
129052=>"111010101",
129053=>"000111111",
129054=>"000010011",
129055=>"100111111",
129056=>"111101101",
129057=>"000111010",
129058=>"111100111",
129059=>"000111101",
129060=>"001001010",
129061=>"000011010",
129062=>"000000000",
129063=>"000000000",
129064=>"010101110",
129065=>"111101010",
129066=>"111110111",
129067=>"111111111",
129068=>"001111111",
129069=>"000111001",
129070=>"011111000",
129071=>"111111101",
129072=>"000100100",
129073=>"000111000",
129074=>"111101101",
129075=>"111111011",
129076=>"010000110",
129077=>"000000000",
129078=>"010110110",
129079=>"000010110",
129080=>"000110111",
129081=>"101000100",
129082=>"000000000",
129083=>"111111111",
129084=>"101111111",
129085=>"111111111",
129086=>"101000111",
129087=>"001100111",
129088=>"000111010",
129089=>"000111010",
129090=>"111010110",
129091=>"110111110",
129092=>"000100111",
129093=>"000111111",
129094=>"101000100",
129095=>"001111000",
129096=>"001011111",
129097=>"000000010",
129098=>"001011000",
129099=>"010010111",
129100=>"111111100",
129101=>"100001011",
129102=>"001100110",
129103=>"000111010",
129104=>"111111100",
129105=>"010111100",
129106=>"000000001",
129107=>"000010011",
129108=>"000000000",
129109=>"011111110",
129110=>"000110100",
129111=>"010101000",
129112=>"010000011",
129113=>"111000010",
129114=>"110011111",
129115=>"101110111",
129116=>"001100100",
129117=>"100100100",
129118=>"000000000",
129119=>"011001011",
129120=>"111111111",
129121=>"110110110",
129122=>"000111011",
129123=>"111101001",
129124=>"000000110",
129125=>"111100000",
129126=>"000000000",
129127=>"100101110",
129128=>"000100100",
129129=>"111001011",
129130=>"010100000",
129131=>"000010100",
129132=>"101000000",
129133=>"100000110",
129134=>"000000000",
129135=>"000110011",
129136=>"011011111",
129137=>"010000000",
129138=>"000011111",
129139=>"100111111",
129140=>"101110110",
129141=>"010010110",
129142=>"100000111",
129143=>"000000011",
129144=>"011000110",
129145=>"100000000",
129146=>"010110111",
129147=>"000100111",
129148=>"010001000",
129149=>"001011010",
129150=>"000111010",
129151=>"110100110",
129152=>"001111111",
129153=>"010010010",
129154=>"000000000",
129155=>"000111011",
129156=>"001111111",
129157=>"111111101",
129158=>"100110111",
129159=>"111110000",
129160=>"101110101",
129161=>"111001001",
129162=>"000000000",
129163=>"011110000",
129164=>"001101100",
129165=>"000000000",
129166=>"000000101",
129167=>"001000001",
129168=>"011011011",
129169=>"010110010",
129170=>"101000111",
129171=>"010001001",
129172=>"000100100",
129173=>"111100000",
129174=>"011010010",
129175=>"110111111",
129176=>"111101111",
129177=>"010000010",
129178=>"011011010",
129179=>"010011010",
129180=>"110100000",
129181=>"100010011",
129182=>"111101101",
129183=>"111010001",
129184=>"111011001",
129185=>"110110000",
129186=>"011111011",
129187=>"011000000",
129188=>"100000000",
129189=>"011011111",
129190=>"001011011",
129191=>"101000110",
129192=>"011011111",
129193=>"111101100",
129194=>"000000010",
129195=>"101110101",
129196=>"011110011",
129197=>"000101101",
129198=>"101010000",
129199=>"110111011",
129200=>"011011000",
129201=>"111001100",
129202=>"000100111",
129203=>"111011011",
129204=>"000011110",
129205=>"000101010",
129206=>"010011100",
129207=>"000100110",
129208=>"100100000",
129209=>"001001001",
129210=>"000000000",
129211=>"000101111",
129212=>"101111111",
129213=>"100010110",
129214=>"110100110",
129215=>"100101000",
129216=>"111001000",
129217=>"000111010",
129218=>"001100000",
129219=>"111001101",
129220=>"101101101",
129221=>"010001111",
129222=>"111100000",
129223=>"100111011",
129224=>"000000000",
129225=>"111010111",
129226=>"101001001",
129227=>"000000000",
129228=>"000000010",
129229=>"100000000",
129230=>"000110110",
129231=>"000111011",
129232=>"101100111",
129233=>"111111111",
129234=>"101001000",
129235=>"101001111",
129236=>"010010010",
129237=>"001001000",
129238=>"111111011",
129239=>"000110111",
129240=>"000000100",
129241=>"000001001",
129242=>"111111001",
129243=>"111000101",
129244=>"110111110",
129245=>"111111100",
129246=>"000000000",
129247=>"100110111",
129248=>"000001001",
129249=>"000100010",
129250=>"000000000",
129251=>"000011000",
129252=>"011000101",
129253=>"101100000",
129254=>"110000001",
129255=>"000000010",
129256=>"011111100",
129257=>"001000000",
129258=>"001000111",
129259=>"000100000",
129260=>"011000000",
129261=>"000001001",
129262=>"110111101",
129263=>"000000000",
129264=>"010010000",
129265=>"011100110",
129266=>"011010111",
129267=>"000000111",
129268=>"001011011",
129269=>"011011000",
129270=>"111011011",
129271=>"101010010",
129272=>"000000000",
129273=>"111111111",
129274=>"101100111",
129275=>"100010100",
129276=>"101000101",
129277=>"101101110",
129278=>"100100100",
129279=>"111111111",
129280=>"011001000",
129281=>"110110110",
129282=>"001100011",
129283=>"100010110",
129284=>"001011111",
129285=>"100010010",
129286=>"111011001",
129287=>"010111001",
129288=>"000000010",
129289=>"100110100",
129290=>"111100001",
129291=>"010001111",
129292=>"111110110",
129293=>"111000000",
129294=>"101011101",
129295=>"011101111",
129296=>"110010010",
129297=>"100110000",
129298=>"001001001",
129299=>"000110110",
129300=>"001111101",
129301=>"100111110",
129302=>"111001011",
129303=>"001111001",
129304=>"101001001",
129305=>"101101001",
129306=>"111111110",
129307=>"110110110",
129308=>"001001001",
129309=>"111000011",
129310=>"110100110",
129311=>"001000001",
129312=>"001100100",
129313=>"101001101",
129314=>"011011000",
129315=>"100110110",
129316=>"001011011",
129317=>"001001011",
129318=>"110110110",
129319=>"110110100",
129320=>"001011001",
129321=>"000000000",
129322=>"110110100",
129323=>"110011110",
129324=>"101111111",
129325=>"001110111",
129326=>"110000010",
129327=>"001001011",
129328=>"111001101",
129329=>"001101001",
129330=>"110101111",
129331=>"110010100",
129332=>"100010100",
129333=>"010110000",
129334=>"100110110",
129335=>"110110100",
129336=>"110100000",
129337=>"100000001",
129338=>"001001001",
129339=>"110010100",
129340=>"100111100",
129341=>"001001011",
129342=>"100010010",
129343=>"010000000",
129344=>"110101111",
129345=>"111110110",
129346=>"111111001",
129347=>"111110100",
129348=>"001001011",
129349=>"010000000",
129350=>"001111111",
129351=>"111000000",
129352=>"111011110",
129353=>"000111110",
129354=>"100010000",
129355=>"000000100",
129356=>"110110110",
129357=>"011001001",
129358=>"001001000",
129359=>"011001111",
129360=>"011010001",
129361=>"000001000",
129362=>"110111111",
129363=>"111001001",
129364=>"000000011",
129365=>"110110110",
129366=>"011001001",
129367=>"100000000",
129368=>"100000010",
129369=>"001011111",
129370=>"000100101",
129371=>"101000100",
129372=>"110110110",
129373=>"001001011",
129374=>"110110110",
129375=>"110110111",
129376=>"110110110",
129377=>"100110110",
129378=>"101110111",
129379=>"001001111",
129380=>"001000000",
129381=>"101010100",
129382=>"100001000",
129383=>"110000000",
129384=>"110110100",
129385=>"010100101",
129386=>"110110111",
129387=>"010110111",
129388=>"011011110",
129389=>"001101001",
129390=>"000000110",
129391=>"011011110",
129392=>"011101011",
129393=>"110110111",
129394=>"110100100",
129395=>"001011011",
129396=>"110110110",
129397=>"001100000",
129398=>"100100111",
129399=>"110110110",
129400=>"110110010",
129401=>"001001111",
129402=>"001001100",
129403=>"001001001",
129404=>"010010010",
129405=>"100000000",
129406=>"110000001",
129407=>"110000001",
129408=>"010000000",
129409=>"000000110",
129410=>"110110110",
129411=>"000010110",
129412=>"111000100",
129413=>"001101011",
129414=>"001011010",
129415=>"000100001",
129416=>"001011011",
129417=>"010110110",
129418=>"011111001",
129419=>"000110111",
129420=>"011011001",
129421=>"100100111",
129422=>"111101101",
129423=>"010000110",
129424=>"101001001",
129425=>"001101111",
129426=>"011010111",
129427=>"110101110",
129428=>"000101010",
129429=>"100110110",
129430=>"001111101",
129431=>"001011111",
129432=>"001011100",
129433=>"111000111",
129434=>"101001101",
129435=>"010000010",
129436=>"000111100",
129437=>"110110100",
129438=>"110110110",
129439=>"001000000",
129440=>"001001001",
129441=>"001001010",
129442=>"011010001",
129443=>"101111111",
129444=>"110000111",
129445=>"000001000",
129446=>"010001011",
129447=>"101101011",
129448=>"110010010",
129449=>"000110110",
129450=>"001001000",
129451=>"000010010",
129452=>"011001000",
129453=>"011011110",
129454=>"000010010",
129455=>"000000000",
129456=>"011111000",
129457=>"111110010",
129458=>"001001001",
129459=>"000000000",
129460=>"001110000",
129461=>"111111111",
129462=>"111111000",
129463=>"001011111",
129464=>"011001001",
129465=>"111001111",
129466=>"111101001",
129467=>"110111000",
129468=>"000000000",
129469=>"001011011",
129470=>"011111111",
129471=>"110000001",
129472=>"001011011",
129473=>"110110110",
129474=>"010111111",
129475=>"011011000",
129476=>"001001001",
129477=>"000000111",
129478=>"101111111",
129479=>"101101101",
129480=>"010001001",
129481=>"011001000",
129482=>"110101100",
129483=>"110010110",
129484=>"001011011",
129485=>"111111111",
129486=>"110110100",
129487=>"111110000",
129488=>"001001001",
129489=>"010001000",
129490=>"110011011",
129491=>"001001001",
129492=>"101100111",
129493=>"100110101",
129494=>"100101110",
129495=>"110110110",
129496=>"000001011",
129497=>"010010110",
129498=>"001001000",
129499=>"001111001",
129500=>"111111000",
129501=>"111011001",
129502=>"011001001",
129503=>"110110110",
129504=>"000010010",
129505=>"000000100",
129506=>"110000000",
129507=>"001101001",
129508=>"011110110",
129509=>"110011011",
129510=>"011000000",
129511=>"111101110",
129512=>"111000110",
129513=>"111010010",
129514=>"101101001",
129515=>"001001001",
129516=>"000110110",
129517=>"010111111",
129518=>"001001011",
129519=>"001000100",
129520=>"010100111",
129521=>"111011001",
129522=>"110010100",
129523=>"111111000",
129524=>"000001111",
129525=>"100100111",
129526=>"000100110",
129527=>"010110000",
129528=>"100110111",
129529=>"100101110",
129530=>"101101001",
129531=>"111011101",
129532=>"011011011",
129533=>"001001001",
129534=>"001001101",
129535=>"001011000",
129536=>"001001101",
129537=>"100111111",
129538=>"000000100",
129539=>"000000110",
129540=>"001001000",
129541=>"000100000",
129542=>"000000111",
129543=>"011000000",
129544=>"010100111",
129545=>"111111100",
129546=>"000000000",
129547=>"000100111",
129548=>"100000111",
129549=>"000101111",
129550=>"000000011",
129551=>"100111111",
129552=>"111110000",
129553=>"101000000",
129554=>"111101111",
129555=>"111001000",
129556=>"011111111",
129557=>"100000000",
129558=>"011011001",
129559=>"000111111",
129560=>"000000011",
129561=>"001101001",
129562=>"000000010",
129563=>"011011000",
129564=>"000000010",
129565=>"000100000",
129566=>"100100111",
129567=>"111010000",
129568=>"000000101",
129569=>"110101111",
129570=>"111111001",
129571=>"010000000",
129572=>"011011011",
129573=>"000001001",
129574=>"011111000",
129575=>"010011101",
129576=>"111111000",
129577=>"111111101",
129578=>"100110100",
129579=>"011000000",
129580=>"110100110",
129581=>"100111111",
129582=>"101101101",
129583=>"100100000",
129584=>"000100111",
129585=>"011010100",
129586=>"100110111",
129587=>"111000000",
129588=>"000000000",
129589=>"111101000",
129590=>"011011011",
129591=>"101111111",
129592=>"001000100",
129593=>"000000101",
129594=>"100001011",
129595=>"010111000",
129596=>"110011111",
129597=>"110111110",
129598=>"000100111",
129599=>"110111010",
129600=>"011000101",
129601=>"100001010",
129602=>"110000101",
129603=>"010010100",
129604=>"111100000",
129605=>"100100110",
129606=>"000100101",
129607=>"011001011",
129608=>"001010101",
129609=>"000000101",
129610=>"000000000",
129611=>"100100110",
129612=>"100000000",
129613=>"110100100",
129614=>"111011000",
129615=>"101101111",
129616=>"100000001",
129617=>"010001000",
129618=>"000101110",
129619=>"001000000",
129620=>"000000000",
129621=>"110011011",
129622=>"101110011",
129623=>"000000010",
129624=>"111111110",
129625=>"110000111",
129626=>"011111100",
129627=>"111110000",
129628=>"000000011",
129629=>"000000111",
129630=>"011011000",
129631=>"011010001",
129632=>"111111011",
129633=>"110101101",
129634=>"000000111",
129635=>"110101100",
129636=>"100000011",
129637=>"111101000",
129638=>"000000011",
129639=>"011000000",
129640=>"111111111",
129641=>"111000100",
129642=>"111000000",
129643=>"000000001",
129644=>"111011111",
129645=>"000000011",
129646=>"111111001",
129647=>"001001111",
129648=>"101111000",
129649=>"100111111",
129650=>"000010110",
129651=>"011000000",
129652=>"000000111",
129653=>"100000000",
129654=>"001000100",
129655=>"001000001",
129656=>"000100000",
129657=>"011000110",
129658=>"111111111",
129659=>"101100000",
129660=>"111110011",
129661=>"100100000",
129662=>"010010001",
129663=>"000000100",
129664=>"111111000",
129665=>"100001110",
129666=>"111000011",
129667=>"111001100",
129668=>"101100000",
129669=>"101101110",
129670=>"100000000",
129671=>"010100000",
129672=>"100100110",
129673=>"000000000",
129674=>"000000000",
129675=>"111000011",
129676=>"000110000",
129677=>"000000000",
129678=>"100000111",
129679=>"000000000",
129680=>"110011011",
129681=>"111111111",
129682=>"000110010",
129683=>"101100101",
129684=>"100100100",
129685=>"000100000",
129686=>"000111111",
129687=>"001001010",
129688=>"000001111",
129689=>"000000111",
129690=>"101100111",
129691=>"000100111",
129692=>"111100101",
129693=>"111100001",
129694=>"000111011",
129695=>"011010011",
129696=>"100111111",
129697=>"000010110",
129698=>"111001000",
129699=>"000000101",
129700=>"100101110",
129701=>"011001100",
129702=>"110110000",
129703=>"110100000",
129704=>"100101111",
129705=>"100011010",
129706=>"111011010",
129707=>"010110110",
129708=>"111100010",
129709=>"000000101",
129710=>"011001001",
129711=>"011000011",
129712=>"000100011",
129713=>"110000001",
129714=>"000000010",
129715=>"110010111",
129716=>"001000101",
129717=>"000000111",
129718=>"111110100",
129719=>"100100001",
129720=>"011100001",
129721=>"001111110",
129722=>"001111001",
129723=>"100000000",
129724=>"000000000",
129725=>"111111111",
129726=>"111101001",
129727=>"010011100",
129728=>"100000101",
129729=>"100000111",
129730=>"000010011",
129731=>"000000011",
129732=>"000101111",
129733=>"101101111",
129734=>"110100110",
129735=>"011000000",
129736=>"111111111",
129737=>"011011010",
129738=>"101111111",
129739=>"100101111",
129740=>"001100110",
129741=>"111111000",
129742=>"101010011",
129743=>"011111111",
129744=>"010000000",
129745=>"110000100",
129746=>"111101101",
129747=>"111111011",
129748=>"011000000",
129749=>"101100110",
129750=>"000000111",
129751=>"000101111",
129752=>"011010000",
129753=>"101100110",
129754=>"111101111",
129755=>"000000100",
129756=>"111011100",
129757=>"111000010",
129758=>"110100011",
129759=>"000000000",
129760=>"000010010",
129761=>"000100101",
129762=>"010010000",
129763=>"000010110",
129764=>"100000000",
129765=>"111011100",
129766=>"001000000",
129767=>"001100101",
129768=>"111100000",
129769=>"001001001",
129770=>"100100000",
129771=>"100000101",
129772=>"111111000",
129773=>"111111000",
129774=>"100000000",
129775=>"101011111",
129776=>"111111000",
129777=>"110101111",
129778=>"101000000",
129779=>"110000100",
129780=>"000100100",
129781=>"010000001",
129782=>"000000000",
129783=>"011001111",
129784=>"000011111",
129785=>"111100110",
129786=>"100000010",
129787=>"000101101",
129788=>"110110111",
129789=>"101000000",
129790=>"000000001",
129791=>"000000000",
129792=>"100101101",
129793=>"111000010",
129794=>"010010000",
129795=>"100000000",
129796=>"111111110",
129797=>"111101101",
129798=>"101111110",
129799=>"110100000",
129800=>"111110111",
129801=>"000000100",
129802=>"100100011",
129803=>"000000000",
129804=>"111000100",
129805=>"000001101",
129806=>"000100011",
129807=>"111101111",
129808=>"000110111",
129809=>"000000011",
129810=>"000000011",
129811=>"111000100",
129812=>"000010000",
129813=>"111110111",
129814=>"111111011",
129815=>"101111011",
129816=>"101000011",
129817=>"000000001",
129818=>"111000011",
129819=>"000000000",
129820=>"101100000",
129821=>"111111111",
129822=>"000001110",
129823=>"000000001",
129824=>"111011000",
129825=>"000000000",
129826=>"110000101",
129827=>"101000111",
129828=>"000110010",
129829=>"001001000",
129830=>"110010010",
129831=>"000000000",
129832=>"111111010",
129833=>"000000011",
129834=>"000000101",
129835=>"110001000",
129836=>"010010001",
129837=>"111000111",
129838=>"110000101",
129839=>"000000000",
129840=>"111011000",
129841=>"011101111",
129842=>"011011011",
129843=>"000110100",
129844=>"100101111",
129845=>"101101111",
129846=>"010011011",
129847=>"000100001",
129848=>"110101100",
129849=>"000000001",
129850=>"011000000",
129851=>"010000000",
129852=>"001000001",
129853=>"111111111",
129854=>"101000001",
129855=>"111101101",
129856=>"110100010",
129857=>"111000010",
129858=>"000100100",
129859=>"100001101",
129860=>"101100100",
129861=>"000000001",
129862=>"101101111",
129863=>"111001101",
129864=>"001110010",
129865=>"100000000",
129866=>"101100000",
129867=>"101010010",
129868=>"010000000",
129869=>"100100111",
129870=>"101011111",
129871=>"000100000",
129872=>"100101101",
129873=>"111111000",
129874=>"100000000",
129875=>"110001000",
129876=>"111111000",
129877=>"100111111",
129878=>"000011011",
129879=>"000000100",
129880=>"001000101",
129881=>"000000001",
129882=>"011101011",
129883=>"010011111",
129884=>"011000100",
129885=>"010110100",
129886=>"000111010",
129887=>"101000110",
129888=>"111100101",
129889=>"000000000",
129890=>"100000100",
129891=>"011011001",
129892=>"001001001",
129893=>"000010111",
129894=>"000000000",
129895=>"100111011",
129896=>"000000101",
129897=>"100111010",
129898=>"111010010",
129899=>"000000000",
129900=>"000000000",
129901=>"000111011",
129902=>"000000000",
129903=>"000000111",
129904=>"100100110",
129905=>"000000010",
129906=>"110010110",
129907=>"000001010",
129908=>"111110000",
129909=>"000101101",
129910=>"111000101",
129911=>"000000000",
129912=>"111111000",
129913=>"100101010",
129914=>"000110111",
129915=>"111101111",
129916=>"001111110",
129917=>"011011001",
129918=>"011011111",
129919=>"101000101",
129920=>"000000101",
129921=>"000000000",
129922=>"000000110",
129923=>"000000100",
129924=>"000101000",
129925=>"110011000",
129926=>"100100010",
129927=>"000000000",
129928=>"000000000",
129929=>"000000100",
129930=>"100111010",
129931=>"001101010",
129932=>"000111101",
129933=>"111100101",
129934=>"111101000",
129935=>"000000101",
129936=>"101000000",
129937=>"111111111",
129938=>"011011101",
129939=>"111111100",
129940=>"000100000",
129941=>"101101110",
129942=>"101000000",
129943=>"011111101",
129944=>"111101101",
129945=>"111011011",
129946=>"111010000",
129947=>"010000000",
129948=>"101000000",
129949=>"000100000",
129950=>"111111110",
129951=>"101100101",
129952=>"110111011",
129953=>"011011111",
129954=>"111000001",
129955=>"000000000",
129956=>"000010111",
129957=>"011100001",
129958=>"010010000",
129959=>"011100000",
129960=>"000101110",
129961=>"111001100",
129962=>"111000100",
129963=>"101000100",
129964=>"000001001",
129965=>"111000000",
129966=>"011111111",
129967=>"000000101",
129968=>"111000101",
129969=>"000000100",
129970=>"011101101",
129971=>"000100110",
129972=>"011001000",
129973=>"111100111",
129974=>"000000100",
129975=>"000011100",
129976=>"000100100",
129977=>"001001011",
129978=>"011111111",
129979=>"011011000",
129980=>"100111000",
129981=>"000000000",
129982=>"111100111",
129983=>"000111111",
129984=>"000100100",
129985=>"000000000",
129986=>"000111011",
129987=>"010000100",
129988=>"000000001",
129989=>"011000010",
129990=>"000000000",
129991=>"111000000",
129992=>"111101111",
129993=>"000000000",
129994=>"000101111",
129995=>"100000000",
129996=>"111111011",
129997=>"110100001",
129998=>"100000000",
129999=>"000111011",
130000=>"000010010",
130001=>"100001000",
130002=>"000000000",
130003=>"001111011",
130004=>"000000000",
130005=>"101101001",
130006=>"111000000",
130007=>"011111011",
130008=>"111011111",
130009=>"000010111",
130010=>"011110111",
130011=>"111110000",
130012=>"111111110",
130013=>"001111100",
130014=>"000000100",
130015=>"000110110",
130016=>"010000010",
130017=>"000000011",
130018=>"111111111",
130019=>"001101110",
130020=>"001011010",
130021=>"000100101",
130022=>"000000100",
130023=>"100110100",
130024=>"011011000",
130025=>"111111100",
130026=>"001011111",
130027=>"101000100",
130028=>"001000110",
130029=>"000100000",
130030=>"111111001",
130031=>"111000001",
130032=>"000000010",
130033=>"110100001",
130034=>"100101100",
130035=>"110110101",
130036=>"001111011",
130037=>"110011110",
130038=>"000000001",
130039=>"000111111",
130040=>"000100010",
130041=>"011010110",
130042=>"111000111",
130043=>"000110011",
130044=>"111011011",
130045=>"100010111",
130046=>"111010000",
130047=>"100000100",
130048=>"100101000",
130049=>"000000100",
130050=>"111000001",
130051=>"011000000",
130052=>"010111011",
130053=>"000000111",
130054=>"111111000",
130055=>"110111111",
130056=>"100110110",
130057=>"010000001",
130058=>"100000001",
130059=>"100100101",
130060=>"000110010",
130061=>"000010111",
130062=>"000001100",
130063=>"111111000",
130064=>"010000000",
130065=>"010000000",
130066=>"110111000",
130067=>"000000111",
130068=>"111000111",
130069=>"111000000",
130070=>"111101100",
130071=>"110111011",
130072=>"010111010",
130073=>"001000000",
130074=>"111000000",
130075=>"000000010",
130076=>"010000010",
130077=>"001101000",
130078=>"000000000",
130079=>"001001000",
130080=>"111111001",
130081=>"101010010",
130082=>"000101101",
130083=>"001111001",
130084=>"010011001",
130085=>"111000111",
130086=>"111101000",
130087=>"011011000",
130088=>"111100000",
130089=>"010000001",
130090=>"101101000",
130091=>"000000000",
130092=>"010111101",
130093=>"111000111",
130094=>"100111001",
130095=>"000110110",
130096=>"111000110",
130097=>"100111011",
130098=>"101101000",
130099=>"000000100",
130100=>"001001000",
130101=>"001101101",
130102=>"000100000",
130103=>"010000001",
130104=>"110110100",
130105=>"001001000",
130106=>"000101101",
130107=>"000010100",
130108=>"001110111",
130109=>"010111111",
130110=>"101001101",
130111=>"111011111",
130112=>"000101111",
130113=>"010111101",
130114=>"010010001",
130115=>"010111001",
130116=>"111101000",
130117=>"101000001",
130118=>"010110111",
130119=>"000111101",
130120=>"011001101",
130121=>"101010010",
130122=>"000001011",
130123=>"111001000",
130124=>"111101001",
130125=>"011011011",
130126=>"110111110",
130127=>"101111010",
130128=>"111100000",
130129=>"110111111",
130130=>"111101001",
130131=>"000001000",
130132=>"000000000",
130133=>"011000000",
130134=>"100100000",
130135=>"010000000",
130136=>"111011000",
130137=>"000110001",
130138=>"111111000",
130139=>"110110111",
130140=>"110111001",
130141=>"100110100",
130142=>"010011110",
130143=>"000000001",
130144=>"101100000",
130145=>"110100000",
130146=>"000010010",
130147=>"111111001",
130148=>"000000000",
130149=>"000001101",
130150=>"000000111",
130151=>"001001100",
130152=>"110000010",
130153=>"000111111",
130154=>"111111101",
130155=>"010111001",
130156=>"111111001",
130157=>"011100110",
130158=>"000000011",
130159=>"110000110",
130160=>"011110110",
130161=>"010111111",
130162=>"010000000",
130163=>"000000001",
130164=>"000001110",
130165=>"111001101",
130166=>"101000010",
130167=>"101111001",
130168=>"010111110",
130169=>"101110101",
130170=>"101101000",
130171=>"000000111",
130172=>"001000100",
130173=>"010000001",
130174=>"011110100",
130175=>"111000000",
130176=>"000011011",
130177=>"011111000",
130178=>"010110110",
130179=>"000111111",
130180=>"001010111",
130181=>"011011101",
130182=>"110111111",
130183=>"111000000",
130184=>"100011011",
130185=>"111000111",
130186=>"111100100",
130187=>"010000111",
130188=>"000000001",
130189=>"111111101",
130190=>"011000001",
130191=>"100001000",
130192=>"001111110",
130193=>"000011111",
130194=>"000000101",
130195=>"101100000",
130196=>"111000110",
130197=>"000110001",
130198=>"111111111",
130199=>"100111100",
130200=>"101100001",
130201=>"000101000",
130202=>"000000011",
130203=>"000010010",
130204=>"011101000",
130205=>"110110110",
130206=>"011001000",
130207=>"111101001",
130208=>"011101111",
130209=>"111101011",
130210=>"000111101",
130211=>"111100000",
130212=>"000000001",
130213=>"010000011",
130214=>"111011001",
130215=>"000000000",
130216=>"000000000",
130217=>"111000000",
130218=>"000010110",
130219=>"111001001",
130220=>"110101110",
130221=>"111101100",
130222=>"101011001",
130223=>"111000000",
130224=>"100111111",
130225=>"110110000",
130226=>"110100000",
130227=>"000000100",
130228=>"101111110",
130229=>"001001011",
130230=>"111101100",
130231=>"001011010",
130232=>"100011011",
130233=>"111000001",
130234=>"000111110",
130235=>"011010010",
130236=>"001001011",
130237=>"111111111",
130238=>"000000011",
130239=>"000110111",
130240=>"111100100",
130241=>"000000000",
130242=>"110011010",
130243=>"001011011",
130244=>"111000101",
130245=>"111001010",
130246=>"000111111",
130247=>"000010010",
130248=>"100110000",
130249=>"000000000",
130250=>"010101000",
130251=>"111101101",
130252=>"011111111",
130253=>"100001001",
130254=>"111111110",
130255=>"111001010",
130256=>"000000111",
130257=>"011001001",
130258=>"111000010",
130259=>"111111100",
130260=>"000010111",
130261=>"010011011",
130262=>"000000000",
130263=>"111111111",
130264=>"000000101",
130265=>"111100111",
130266=>"000100101",
130267=>"110000111",
130268=>"100101001",
130269=>"111101010",
130270=>"111101100",
130271=>"001000000",
130272=>"111110111",
130273=>"001111010",
130274=>"001000000",
130275=>"111000000",
130276=>"010000000",
130277=>"000000101",
130278=>"100000000",
130279=>"111111100",
130280=>"000111111",
130281=>"111111101",
130282=>"011100100",
130283=>"001000000",
130284=>"101111000",
130285=>"111100001",
130286=>"110000101",
130287=>"000000000",
130288=>"111101100",
130289=>"100100100",
130290=>"101001000",
130291=>"000010110",
130292=>"001101000",
130293=>"010111101",
130294=>"111000000",
130295=>"000000010",
130296=>"111111000",
130297=>"010110111",
130298=>"100000000",
130299=>"111101111",
130300=>"111111000",
130301=>"000010000",
130302=>"101111110",
130303=>"110000000",
130304=>"001000000",
130305=>"000000111",
130306=>"000100100",
130307=>"000011001",
130308=>"011000100",
130309=>"111000000",
130310=>"000000011",
130311=>"100110110",
130312=>"000000001",
130313=>"000011001",
130314=>"011111010",
130315=>"000011000",
130316=>"000100101",
130317=>"000000010",
130318=>"001011001",
130319=>"110111010",
130320=>"010011011",
130321=>"010011011",
130322=>"000100111",
130323=>"011100111",
130324=>"000100000",
130325=>"100100101",
130326=>"111001010",
130327=>"001000011",
130328=>"011000011",
130329=>"100100111",
130330=>"010000110",
130331=>"011011000",
130332=>"000000001",
130333=>"101101100",
130334=>"011000000",
130335=>"000100100",
130336=>"000000000",
130337=>"010000111",
130338=>"101010011",
130339=>"111101010",
130340=>"010100000",
130341=>"011001001",
130342=>"100100110",
130343=>"000111010",
130344=>"010100101",
130345=>"011111011",
130346=>"100010000",
130347=>"111110111",
130348=>"011011011",
130349=>"111100000",
130350=>"101101100",
130351=>"110100000",
130352=>"010000011",
130353=>"111111111",
130354=>"100100010",
130355=>"000111111",
130356=>"011111000",
130357=>"011111101",
130358=>"110000001",
130359=>"000100000",
130360=>"000001000",
130361=>"000000110",
130362=>"100100111",
130363=>"000010110",
130364=>"110111000",
130365=>"100100110",
130366=>"000000000",
130367=>"001001101",
130368=>"111111011",
130369=>"011001000",
130370=>"100001010",
130371=>"001011000",
130372=>"000000000",
130373=>"001000000",
130374=>"000100011",
130375=>"011111001",
130376=>"100101101",
130377=>"010001111",
130378=>"101100000",
130379=>"000000111",
130380=>"010011010",
130381=>"110011111",
130382=>"100110110",
130383=>"010010011",
130384=>"100100100",
130385=>"010000011",
130386=>"111011101",
130387=>"001000000",
130388=>"000010000",
130389=>"110100001",
130390=>"010001000",
130391=>"000010000",
130392=>"000101001",
130393=>"110010010",
130394=>"010110000",
130395=>"110110110",
130396=>"101100101",
130397=>"000000000",
130398=>"011011010",
130399=>"110011000",
130400=>"101001001",
130401=>"010101111",
130402=>"101001101",
130403=>"001011000",
130404=>"000000000",
130405=>"000001000",
130406=>"000100010",
130407=>"100101101",
130408=>"000011010",
130409=>"000100100",
130410=>"111011010",
130411=>"011011101",
130412=>"000101000",
130413=>"111111000",
130414=>"100100111",
130415=>"011011111",
130416=>"110001001",
130417=>"000010011",
130418=>"001100110",
130419=>"101000000",
130420=>"000000011",
130421=>"100100010",
130422=>"000111111",
130423=>"111000000",
130424=>"011000100",
130425=>"111000000",
130426=>"000001011",
130427=>"111100101",
130428=>"000110010",
130429=>"110000000",
130430=>"100100111",
130431=>"100001100",
130432=>"011010000",
130433=>"011011000",
130434=>"000000111",
130435=>"111101100",
130436=>"100000100",
130437=>"100111100",
130438=>"011110100",
130439=>"000001100",
130440=>"110000100",
130441=>"000111111",
130442=>"000000000",
130443=>"011000110",
130444=>"100100000",
130445=>"101100101",
130446=>"111011010",
130447=>"100001001",
130448=>"011001101",
130449=>"000010011",
130450=>"000000000",
130451=>"100000011",
130452=>"100111011",
130453=>"000000000",
130454=>"111011011",
130455=>"101001000",
130456=>"011011000",
130457=>"110101111",
130458=>"100000010",
130459=>"011010000",
130460=>"100100000",
130461=>"011011010",
130462=>"000111110",
130463=>"100101100",
130464=>"001001110",
130465=>"010011010",
130466=>"100100000",
130467=>"000000010",
130468=>"010100111",
130469=>"000000000",
130470=>"010011101",
130471=>"000000000",
130472=>"011010111",
130473=>"011111011",
130474=>"110100101",
130475=>"000000000",
130476=>"111111000",
130477=>"100000000",
130478=>"100101001",
130479=>"000000000",
130480=>"100100010",
130481=>"000110110",
130482=>"000100000",
130483=>"000100000",
130484=>"111110100",
130485=>"101111111",
130486=>"111100100",
130487=>"001011001",
130488=>"101101100",
130489=>"101111111",
130490=>"011001000",
130491=>"011000000",
130492=>"000101100",
130493=>"111111111",
130494=>"110110010",
130495=>"100111111",
130496=>"000100111",
130497=>"000000000",
130498=>"000000101",
130499=>"100100100",
130500=>"000000010",
130501=>"010010000",
130502=>"011000001",
130503=>"000001111",
130504=>"101101011",
130505=>"111000000",
130506=>"000000100",
130507=>"101011010",
130508=>"100001111",
130509=>"000001011",
130510=>"000110000",
130511=>"100011111",
130512=>"000110111",
130513=>"110110100",
130514=>"000110011",
130515=>"010111010",
130516=>"000100111",
130517=>"100101100",
130518=>"000111011",
130519=>"000001011",
130520=>"100101111",
130521=>"111100100",
130522=>"010100000",
130523=>"100100110",
130524=>"111011011",
130525=>"011111100",
130526=>"111111111",
130527=>"010011001",
130528=>"000000100",
130529=>"000000011",
130530=>"111100111",
130531=>"000101001",
130532=>"000100000",
130533=>"000001111",
130534=>"000000011",
130535=>"001000100",
130536=>"100100000",
130537=>"100100111",
130538=>"111111110",
130539=>"001100111",
130540=>"001000000",
130541=>"000010111",
130542=>"000100000",
130543=>"101111100",
130544=>"011010011",
130545=>"111011101",
130546=>"000010111",
130547=>"101011101",
130548=>"110110000",
130549=>"111111111",
130550=>"100110000",
130551=>"011011101",
130552=>"000000101",
130553=>"000101011",
130554=>"110100100",
130555=>"011111111",
130556=>"111011000",
130557=>"011111000",
130558=>"111110000",
130559=>"111010000",
130560=>"011100100",
130561=>"011000010",
130562=>"100101101",
130563=>"000000000",
130564=>"111011000",
130565=>"000001110",
130566=>"100100111",
130567=>"000000010",
130568=>"000000010",
130569=>"000000110",
130570=>"110110010",
130571=>"111000101",
130572=>"111111000",
130573=>"111101100",
130574=>"010000000",
130575=>"001101111",
130576=>"110000010",
130577=>"111111000",
130578=>"101001101",
130579=>"110011001",
130580=>"101000101",
130581=>"100000000",
130582=>"011111110",
130583=>"111010000",
130584=>"111110000",
130585=>"110110011",
130586=>"000011011",
130587=>"011000000",
130588=>"011011001",
130589=>"111110110",
130590=>"001000011",
130591=>"000110101",
130592=>"101101111",
130593=>"010110111",
130594=>"011100111",
130595=>"111000000",
130596=>"001001011",
130597=>"110110100",
130598=>"000010010",
130599=>"111111010",
130600=>"000111111",
130601=>"000001011",
130602=>"010011111",
130603=>"000000000",
130604=>"011011011",
130605=>"111111001",
130606=>"011000000",
130607=>"111111111",
130608=>"111111001",
130609=>"011111111",
130610=>"000000010",
130611=>"010010010",
130612=>"010100111",
130613=>"000000000",
130614=>"011000100",
130615=>"010011111",
130616=>"001011010",
130617=>"010111111",
130618=>"000000100",
130619=>"001000010",
130620=>"110101000",
130621=>"110111111",
130622=>"010000011",
130623=>"001111111",
130624=>"000000111",
130625=>"111111000",
130626=>"101101111",
130627=>"110001101",
130628=>"001101001",
130629=>"000111111",
130630=>"110000010",
130631=>"100101100",
130632=>"000000000",
130633=>"111101111",
130634=>"010000011",
130635=>"000010111",
130636=>"000010010",
130637=>"011001000",
130638=>"100110111",
130639=>"111111111",
130640=>"100100111",
130641=>"110111000",
130642=>"000000000",
130643=>"001011000",
130644=>"010000111",
130645=>"110111000",
130646=>"100110110",
130647=>"111100100",
130648=>"000000000",
130649=>"010011100",
130650=>"000010110",
130651=>"100100111",
130652=>"011101111",
130653=>"001001001",
130654=>"000010010",
130655=>"010100101",
130656=>"111100111",
130657=>"111111001",
130658=>"111000000",
130659=>"000100110",
130660=>"100001010",
130661=>"000111101",
130662=>"000100000",
130663=>"000000000",
130664=>"101111011",
130665=>"000000010",
130666=>"110000111",
130667=>"100010110",
130668=>"000010000",
130669=>"101111111",
130670=>"010000001",
130671=>"111111010",
130672=>"001001011",
130673=>"000000000",
130674=>"111000011",
130675=>"101110111",
130676=>"000100001",
130677=>"000010000",
130678=>"000001000",
130679=>"001000110",
130680=>"101000000",
130681=>"000000000",
130682=>"111111111",
130683=>"111101000",
130684=>"001001110",
130685=>"100001010",
130686=>"111101111",
130687=>"000101111",
130688=>"011000101",
130689=>"001010000",
130690=>"010000000",
130691=>"010010110",
130692=>"000000010",
130693=>"111101001",
130694=>"111111001",
130695=>"001001001",
130696=>"100110011",
130697=>"000000000",
130698=>"000110110",
130699=>"100101111",
130700=>"000000000",
130701=>"000000000",
130702=>"000000001",
130703=>"000000011",
130704=>"100111011",
130705=>"110010001",
130706=>"001000001",
130707=>"010111011",
130708=>"011010000",
130709=>"010110111",
130710=>"011111000",
130711=>"000000100",
130712=>"000000000",
130713=>"000000000",
130714=>"110111111",
130715=>"111000000",
130716=>"000010011",
130717=>"000000010",
130718=>"000100010",
130719=>"101001000",
130720=>"001101101",
130721=>"110000100",
130722=>"111101101",
130723=>"111111111",
130724=>"110011010",
130725=>"100111111",
130726=>"111110011",
130727=>"000011011",
130728=>"110010000",
130729=>"000000010",
130730=>"000101111",
130731=>"110111111",
130732=>"010110000",
130733=>"000100111",
130734=>"110110110",
130735=>"001000111",
130736=>"111111011",
130737=>"000110110",
130738=>"111100101",
130739=>"100110010",
130740=>"111111110",
130741=>"110010000",
130742=>"111011000",
130743=>"011001001",
130744=>"001000000",
130745=>"010010110",
130746=>"010000000",
130747=>"010001001",
130748=>"101000000",
130749=>"000000000",
130750=>"001111011",
130751=>"000000000",
130752=>"101000111",
130753=>"000011111",
130754=>"010010010",
130755=>"011111110",
130756=>"000010101",
130757=>"110110010",
130758=>"011011000",
130759=>"000000000",
130760=>"111111111",
130761=>"010010001",
130762=>"100111010",
130763=>"111111101",
130764=>"111100111",
130765=>"111000000",
130766=>"000101101",
130767=>"100010110",
130768=>"100110100",
130769=>"100100111",
130770=>"000110001",
130771=>"010001111",
130772=>"111000111",
130773=>"000110110",
130774=>"011111001",
130775=>"111111001",
130776=>"111111000",
130777=>"111111001",
130778=>"110111111",
130779=>"000000010",
130780=>"001101000",
130781=>"001010000",
130782=>"101010000",
130783=>"000000010",
130784=>"111111000",
130785=>"010100110",
130786=>"111000001",
130787=>"111111010",
130788=>"110000011",
130789=>"000000000",
130790=>"101011000",
130791=>"001001011",
130792=>"111000001",
130793=>"000000011",
130794=>"000011011",
130795=>"111101101",
130796=>"010111101",
130797=>"011010111",
130798=>"100000000",
130799=>"111001000",
130800=>"110111001",
130801=>"011011110",
130802=>"111000110",
130803=>"101011011",
130804=>"111011001",
130805=>"000000111",
130806=>"101101111",
130807=>"111111101",
130808=>"111011000",
130809=>"000101001",
130810=>"010001111",
130811=>"101110110",
130812=>"111111111",
130813=>"111110011",
130814=>"000000011",
130815=>"000010010",
130816=>"011010011",
130817=>"000000110",
130818=>"100110101",
130819=>"000101111",
130820=>"000000000",
130821=>"000001010",
130822=>"111000111",
130823=>"011111111",
130824=>"100101111",
130825=>"000000101",
130826=>"110011011",
130827=>"100000001",
130828=>"000010000",
130829=>"000100111",
130830=>"001111111",
130831=>"110000110",
130832=>"000000000",
130833=>"000000000",
130834=>"111111111",
130835=>"001001010",
130836=>"011111000",
130837=>"001000000",
130838=>"010001110",
130839=>"010010111",
130840=>"000001101",
130841=>"111111111",
130842=>"000100100",
130843=>"111111111",
130844=>"100111111",
130845=>"101101111",
130846=>"111111110",
130847=>"000000000",
130848=>"000000000",
130849=>"010001001",
130850=>"000000101",
130851=>"000100001",
130852=>"110011011",
130853=>"000010110",
130854=>"000000000",
130855=>"010111111",
130856=>"000000111",
130857=>"111111111",
130858=>"111110111",
130859=>"000000000",
130860=>"011011011",
130861=>"000001111",
130862=>"001100000",
130863=>"011110001",
130864=>"100011000",
130865=>"110011011",
130866=>"000000101",
130867=>"111001000",
130868=>"101000000",
130869=>"110010010",
130870=>"100000010",
130871=>"111111110",
130872=>"111111011",
130873=>"011011111",
130874=>"111100111",
130875=>"000000000",
130876=>"111101011",
130877=>"011111111",
130878=>"000000100",
130879=>"000111100",
130880=>"000000000",
130881=>"011111111",
130882=>"111111111",
130883=>"111101010",
130884=>"111110010",
130885=>"000000000",
130886=>"101000000",
130887=>"010000000",
130888=>"111001111",
130889=>"010010000",
130890=>"010111111",
130891=>"000001000",
130892=>"011011000",
130893=>"000100011",
130894=>"111111011",
130895=>"101101101",
130896=>"001000000",
130897=>"011111111",
130898=>"010111111",
130899=>"111101011",
130900=>"011011011",
130901=>"110001000",
130902=>"110000100",
130903=>"000111111",
130904=>"100000010",
130905=>"111110110",
130906=>"110000000",
130907=>"001110111",
130908=>"111111000",
130909=>"010001011",
130910=>"000000000",
130911=>"011111101",
130912=>"111101011",
130913=>"110001101",
130914=>"000100000",
130915=>"110100010",
130916=>"100100110",
130917=>"111111111",
130918=>"111001000",
130919=>"111101111",
130920=>"111111110",
130921=>"000000000",
130922=>"110111111",
130923=>"011010010",
130924=>"110111001",
130925=>"101100000",
130926=>"000000000",
130927=>"111011000",
130928=>"111111011",
130929=>"011000100",
130930=>"000000010",
130931=>"111101111",
130932=>"010000000",
130933=>"101100000",
130934=>"111111111",
130935=>"000111010",
130936=>"000000000",
130937=>"111111000",
130938=>"000101101",
130939=>"000000010",
130940=>"100100001",
130941=>"111111000",
130942=>"000000000",
130943=>"111111010",
130944=>"111111000",
130945=>"010111000",
130946=>"000001111",
130947=>"000000001",
130948=>"101011111",
130949=>"110011111",
130950=>"110110111",
130951=>"111011001",
130952=>"001111011",
130953=>"101000000",
130954=>"110100110",
130955=>"111111000",
130956=>"000000000",
130957=>"000000000",
130958=>"011010000",
130959=>"111000100",
130960=>"001011111",
130961=>"001011000",
130962=>"101000000",
130963=>"111000010",
130964=>"010100100",
130965=>"010111111",
130966=>"111111010",
130967=>"101001110",
130968=>"000000001",
130969=>"111100101",
130970=>"101100100",
130971=>"000000000",
130972=>"111000100",
130973=>"111111111",
130974=>"111111111",
130975=>"000010011",
130976=>"011010001",
130977=>"110100100",
130978=>"111111011",
130979=>"111101111",
130980=>"110010001",
130981=>"110110110",
130982=>"000000111",
130983=>"100000000",
130984=>"000000011",
130985=>"000000111",
130986=>"111111100",
130987=>"000100100",
130988=>"111001011",
130989=>"111111111",
130990=>"001011011",
130991=>"111001111",
130992=>"000000000",
130993=>"111111001",
130994=>"111100110",
130995=>"110011001",
130996=>"000001001",
130997=>"101101110",
130998=>"000001001",
130999=>"000100000",
131000=>"110110101",
131001=>"110110101",
131002=>"110000000",
131003=>"111010011",
131004=>"111000000",
131005=>"000011000",
131006=>"000010100",
131007=>"101000000",
131008=>"000000000",
131009=>"000000000",
131010=>"011011111",
131011=>"110100010",
131012=>"000001100",
131013=>"011001001",
131014=>"000011010",
131015=>"000100110",
131016=>"101111000",
131017=>"011111010",
131018=>"010010001",
131019=>"000011010",
131020=>"000010000",
131021=>"001101100",
131022=>"111100001",
131023=>"110100100",
131024=>"111101111",
131025=>"100100011",
131026=>"010010111",
131027=>"010010001",
131028=>"100100111",
131029=>"100110000",
131030=>"010111001",
131031=>"000101111",
131032=>"000000010",
131033=>"111011101",
131034=>"100110010",
131035=>"100000000",
131036=>"000100001",
131037=>"000000010",
131038=>"011111010",
131039=>"000001000",
131040=>"010010100",
131041=>"111100100",
131042=>"001010110",
131043=>"100110010",
131044=>"000000100",
131045=>"100000000",
131046=>"000010010",
131047=>"011011111",
131048=>"010011111",
131049=>"100000011",
131050=>"001110110",
131051=>"000100100",
131052=>"011111111",
131053=>"010000001",
131054=>"001101001",
131055=>"101100000",
131056=>"100111010",
131057=>"100110000",
131058=>"111111111",
131059=>"000010010",
131060=>"110101111",
131061=>"000000000",
131062=>"111000000",
131063=>"111111111",
131064=>"000000100",
131065=>"111111111",
131066=>"010010000",
131067=>"010111010",
131068=>"100000100",
131069=>"000000000",
131070=>"110000110",
131071=>"001111111");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;
