LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L2BNROM IS
    PORT (
        coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); -- Instruction bus
        address : IN unsigned(4 DOWNTO 0));
END L2BNROM;

ARCHITECTURE RTL OF L2BNROM IS

    TYPE ROM_mem IS ARRAY (0 TO 31) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem :=
    (0 => "1101100010111110" & "0010111100110111",
    1 => "0100110011010100" & "0001101000100110",
    2 => "0001001000010111" & "0100011110001111",
    3 => "0000111010101000" & "0011101010101000",
    4 => "0001000100101000" & "0100010111010010",
    5 => "0000011100101111" & "0001111000001010",
    6 => "0111111111010010" & "0010010100110010",
    7 => "0100101110011101" & "0001110110110010",
    8 => "1111110100011011" & "0011010011000100",
    9 => "0011001011110101" & "0010001011001001",
    10 => "0001101110101100" & "0011100101001110",
    11 => "1111111000010010" & "0001100010100000",
    12 => "1100001001000000" & "0000111111011010",
    13 => "0001110011001001" & "0100000000011100",
    14 => "0100001011101011" & "0011001000111100",
    15 => "0011100110101111" & "0011101011010101",
    16 => "0001110001000000" & "0100011101110100",
    17 => "0110000001001101" & "0010100011010110",
    18 => "0001001000101000" & "0011000100010000",
    19 => "0010101010010000" & "0010110101000101",
    20 => "0000101100101001" & "0010000101100110",
    21 => "0100010101011011" & "0011010000010010",
    22 => "0010001000010001" & "0011000000000011",
    23 => "0010001010100010" & "0010010111011000",
    24 => "0001101010100100" & "0100010001010010",
    25 => "0010000111101000" & "0011100100111001",
    26 => "0100101111010110" & "0011011111010011",
    27 => "0001111110111100" & "0100000000001001",
    28 => "0010011001100001" & "0010110101010111",
    29 => "0011110111001100" & "0010110011110100",
    30 => "1111000000110110" & "0011100000101111",
    31 => "0001101010101010" & "0010111000101011");
BEGIN
    coefs <= ROM_content(to_integer(address));
END RTL;