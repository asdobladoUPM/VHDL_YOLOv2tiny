LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L1WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(1) DOWNTO 0));
END L1WROM;

ARCHITECTURE RTL OF L1WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 47) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0 => "111000000",
  1 => "110000100",
  2 => "111110100",
  3 => "011011111",
  4 => "101011101",
  5 => "111111101",
  6 => "111111111",
  7 => "111111111",
  8 => "000000000",
  9 => "111111111",
  10 => "000000000",
  11 => "001000100",
  12 => "000011111",
  13 => "000111111",
  14 => "000011111",
  15 => "110100100",
  16 => "000011111",
  17 => "001001011",
  18 => "110010000",
  19 => "110010000",
  20 => "111010000",
  21 => "000000110",
  22 => "101101010",
  23 => "101001010",
  24 => "111101101",
  25 => "111101101",
  26 => "000000101",
  27 => "011011011",
  28 => "011011011",
  29 => "011011011",
  30 => "111110000",
  31 => "111110000",
  32 => "111110000",
  33 => "100100100",
  34 => "100100100",
  35 => "100100100",
  36 => "000000000",
  37 => "111111111",
  38 => "111111111",
  39 => "111000111",
  40 => "111000111",
  41 => "111000111",
  42 => "000001111",
  43 => "000011111",
  44 => "000111111",
  45 => "001101000",
  46 => "000000000",
  47 => "111111111");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;