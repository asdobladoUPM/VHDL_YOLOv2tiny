LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L5BNROM IS
    PORT (
        coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); -- Instruction bus
        address : IN unsigned(9 DOWNTO 0));
END L5BNROM;

ARCHITECTURE RTL OF L5BNROM IS

    TYPE ROM_mem IS ARRAY (0 TO 1023) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem :=
    (0=>"0010000111011100"&"0010000100010011",
1=>"0000111000100011"&"0010001101010101",
2=>"0010100000101011"&"0001111101111000",
3=>"0001001111000001"&"0010000100101000",
4=>"0001000001011010"&"0010010001101111",
5=>"0001101101111011"&"0010001101000001",
6=>"0000101011000110"&"0001110001110011",
7=>"0001101101010001"&"0010010000100101",
8=>"0001101010010100"&"0010001101101111",
9=>"0010100100010100"&"0010100010101101",
10=>"0000111100011011"&"0010001010011010",
11=>"0001100001101011"&"0010001001100101",
12=>"0001011000011011"&"0010010010010101",
13=>"0000110011101111"&"0001111001011000",
14=>"0010011111100101"&"0010000111001100",
15=>"0001100100000001"&"0010010010101101",
16=>"0010000001000010"&"0010010101101010",
17=>"0001000010101111"&"0010010101011111",
18=>"0001111110101100"&"0010010110111101",
19=>"0010000100110000"&"0010010101100011",
20=>"0001010100101110"&"0010101000011001",
21=>"0010000011011010"&"0010001001111110",
22=>"0001100010010111"&"0010001001011010",
23=>"0001010111010110"&"0010001010101001",
24=>"0001110110000010"&"0010001101100111",
25=>"0000010000111011"&"0010000110110101",
26=>"0001111111010101"&"0010001100111001",
27=>"0010001010011100"&"0010000000111101",
28=>"0000111101010100"&"0001110011001010",
29=>"0000111100010101"&"0010000101100011",
30=>"0000111110110000"&"0010001001100101",
31=>"1111010110001101"&"0010000101110101",
32=>"0000110011001011"&"0010011100100111",
33=>"0001000011001011"&"0010000001001110",
34=>"0000011001000000"&"0010010100101101",
35=>"0000000110111100"&"0001110111011011",
36=>"0000010011001111"&"0001111101111100",
37=>"0010100010110000"&"0010010000110110",
38=>"0001100011000001"&"0010001101100011",
39=>"0000100001001010"&"0010000011010011",
40=>"0001001101101100"&"0010001011011000",
41=>"0001101111011100"&"0010001111111001",
42=>"0001000111010001"&"0010010001011011",
43=>"0001001110001000"&"0010001100001111",
44=>"0010101100111110"&"0010000011011100",
45=>"0000101010000100"&"0001011111000010",
46=>"0010000110011111"&"0001110101100101",
47=>"0010100001110110"&"0010001000010101",
48=>"0010101111011011"&"0001111100101011",
49=>"0001111000010101"&"0010001110001000",
50=>"0001011010010111"&"0010011100001010",
51=>"0001111011101111"&"0010001011101010",
52=>"0001011101101010"&"0001100100110100",
53=>"0001000111001110"&"0010010101100101",
54=>"0010001111100010"&"0001100101100111",
55=>"0001011100011111"&"0010001100000101",
56=>"0001001011111001"&"0010100010111110",
57=>"0010000010101100"&"0010001011000111",
58=>"0001100100010000"&"0010001100100011",
59=>"0001000111000111"&"0010001100001101",
60=>"0010010101101111"&"0010001000011010",
61=>"0000110011111001"&"0001110101110001",
62=>"0001010100100110"&"0010010001010010",
63=>"0010001001110110"&"0010000100101001",
64=>"0010010001001101"&"0010001001110110",
65=>"0001000101000110"&"0001111110101000",
66=>"0010010001000111"&"0010001110111010",
67=>"0001011111000111"&"0001011011100110",
68=>"0001111000101011"&"0010000111000001",
69=>"0011001110001101"&"0010001101100000",
70=>"0001010111000111"&"0010010101110101",
71=>"0000110001001111"&"0010010111010101",
72=>"0000101101000010"&"0010010110000101",
73=>"0001011111010001"&"0010010101001000",
74=>"0001000000001100"&"0010001010110000",
75=>"0001101110100010"&"0001111101010111",
76=>"0001010001001111"&"0010011001111100",
77=>"0000010100101001"&"0010011000111100",
78=>"0001101011100001"&"0010001101100011",
79=>"0010001001100111"&"0001110001101010",
80=>"0010011100101011"&"0010011010011000",
81=>"0001110100110101"&"0010001010010110",
82=>"0000000101010010"&"0010001111000010",
83=>"0000101001100110"&"0010010000110001",
84=>"0000111110011011"&"0010011110011000",
85=>"0001010110100100"&"0010001101110010",
86=>"0001000111100111"&"0010011011011100",
87=>"0010000111001010"&"0001111010111001",
88=>"0001010001100001"&"0010010010111110",
89=>"0001010101010101"&"0010001110101001",
90=>"0000111011001011"&"0010000010101001",
91=>"0001001001111001"&"0010001000001001",
92=>"0010000001110001"&"0010010010011111",
93=>"0010001000001110"&"0010001011111010",
94=>"0000101111001000"&"0010001000010110",
95=>"1111111101011001"&"0010011101111111",
96=>"0000101001101100"&"0010011101110111",
97=>"0000110110010010"&"0010010001110011",
98=>"0001100111000000"&"0010010100111011",
99=>"0001010001110101"&"0010010111100110",
100=>"0001011101010110"&"0010011100101100",
101=>"0001000101000001"&"0010000001101000",
102=>"0000111111011011"&"0010000110101010",
103=>"0010011111001101"&"0010000110010001",
104=>"0001101101001010"&"0010001000000110",
105=>"0001001110001101"&"0010010110110111",
106=>"0010000011010010"&"0010000111100011",
107=>"0011011001000011"&"0010001010110111",
108=>"0000111110110100"&"0010011110101010",
109=>"0001000110011001"&"0010011101001100",
110=>"0001110100010010"&"0010000111101010",
111=>"0000011000000101"&"0010000011010110",
112=>"0010001111101110"&"0010010010001011",
113=>"0010000010100101"&"0010000000001001",
114=>"0010010110011111"&"0010010000001111",
115=>"0000010000111100"&"0010001111011111",
116=>"0000111000100101"&"0001111100111001",
117=>"0000010100111100"&"0010001011001111",
118=>"0001111011011000"&"0010011010111110",
119=>"0000000110100100"&"0010001101001010",
120=>"0000010111101010"&"0010011011100110",
121=>"0010110111101110"&"0010000101101100",
122=>"0010001111000001"&"0010010000000000",
123=>"1111111010010110"&"0010001000111000",
124=>"0001011101001011"&"0010000110111100",
125=>"0000100010111010"&"0001110011110010",
126=>"0001111110100001"&"0001111001001111",
127=>"0000100101100011"&"0010001010110001",
128=>"0001110100011011"&"0010000011011011",
129=>"0001110011011100"&"0010010110111000",
130=>"0000101011100101"&"0010000111101111",
131=>"0010000100000101"&"0010011100101001",
132=>"0000111100110000"&"0010000101011000",
133=>"0011110101010101"&"0010000100111001",
134=>"0010010100110110"&"0001110110001011",
135=>"0000100010000111"&"0010010011010011",
136=>"0010110000001011"&"0010010011001000",
137=>"0001011010010010"&"0010001000000001",
138=>"0000010010101000"&"0010000110110101",
139=>"0001100100000001"&"0010011101100100",
140=>"0001001001111011"&"0010011101111001",
141=>"0001010101111110"&"0001101000011101",
142=>"0001001101011010"&"0010001111111101",
143=>"1111110010001000"&"0010000101100000",
144=>"1110010010011110"&"0001101110110100",
145=>"0001011011001101"&"0010000011000000",
146=>"0001110111000000"&"0001111011101100",
147=>"0000001010001100"&"0010000011011001",
148=>"0001101100111011"&"0010001111010100",
149=>"0001111110111001"&"0010010101100000",
150=>"0001101101011101"&"0010011100101010",
151=>"0001110001110100"&"0010001001101111",
152=>"0001111001101001"&"0010011010111011",
153=>"0001110000100011"&"0010011011101001",
154=>"0010000101011010"&"0010011000000101",
155=>"0000110010100110"&"0010010111010000",
156=>"0010000000101111"&"0001111001110001",
157=>"0001100100111100"&"0010000110101111",
158=>"0001011100010101"&"0001101100000011",
159=>"0000110111010110"&"0010011010110000",
160=>"0001010101111100"&"0010001111000000",
161=>"0001010001101000"&"0010000110011100",
162=>"0001000100110110"&"0010001100100111",
163=>"0001100011100110"&"0010000001100010",
164=>"0001111111001100"&"0001110111110011",
165=>"0001000010000110"&"0010010110101010",
166=>"0001001001101010"&"0010011010010111",
167=>"0001010001101100"&"0010000111100111",
168=>"0000110011101101"&"0010010100100011",
169=>"1110101001101000"&"0001011010011111",
170=>"0000110011111111"&"0010001000010010",
171=>"0000011101011011"&"0010001111110100",
172=>"0001101110000010"&"0010001000111111",
173=>"0000101001101110"&"0010000110110101",
174=>"0001111110110001"&"0010001001000011",
175=>"0001001010101000"&"0010000110000010",
176=>"0010000011001001"&"0010011110100000",
177=>"0010001000001000"&"0010010010011100",
178=>"0001110000011101"&"0010001100100101",
179=>"0000001000101000"&"0010011000110011",
180=>"0000110011111101"&"0010001111010110",
181=>"0001110100011000"&"0010001111110000",
182=>"0000100111000111"&"0010011010111011",
183=>"0000100110001010"&"0010100001101001",
184=>"0010110110111110"&"0010011110010000",
185=>"0000101110100100"&"0001110101111110",
186=>"0001000101000111"&"0010001010000111",
187=>"0000100010011100"&"0010010011100101",
188=>"1110110100000010"&"0001111110010101",
189=>"0010000111001111"&"0001011110110110",
190=>"1111110111101000"&"0010000111101111",
191=>"0001010111000010"&"0010010010010001",
192=>"0010010101111000"&"0010001001011010",
193=>"0000111111101111"&"0001101011010011",
194=>"0001100001101100"&"0010000101101111",
195=>"0001110111001101"&"0010001010001010",
196=>"0001011010001011"&"0010000100011000",
197=>"0001100011101110"&"0010010101000000",
198=>"0001000110111001"&"0010011001011100",
199=>"0010010001000101"&"0010010001010111",
200=>"0000000011100110"&"0010000011011111",
201=>"0010110001100010"&"0010001100101100",
202=>"0000010111001111"&"0001111000100111",
203=>"1110111000010000"&"0010000100111111",
204=>"0001101111110000"&"0010010111000011",
205=>"0001010001001000"&"0010000011111011",
206=>"0001001111011001"&"0001111000110001",
207=>"1111011010010100"&"0010010010100110",
208=>"0010011000101110"&"0010001111101100",
209=>"0001110001000011"&"0010011110100000",
210=>"0010001100010111"&"0001100111111100",
211=>"0001011101001000"&"0010010000010011",
212=>"0001011100010011"&"0001100001111001",
213=>"0000110001001100"&"0010011100100001",
214=>"0001110010101010"&"0001111101111110",
215=>"0010001011010000"&"0010001110110101",
216=>"0000100001010100"&"0010001111111011",
217=>"0001011011111000"&"0001111110100010",
218=>"0010011100000110"&"0010000011100000",
219=>"0010000010100011"&"0010011111110100",
220=>"0001101100101010"&"0010010110001001",
221=>"0001100111111001"&"0010011011111010",
222=>"0001111001101101"&"0010011001000001",
223=>"0001001101010010"&"0010010011101100",
224=>"0001111001010001"&"0010000001100001",
225=>"0001010111101100"&"0010011010000011",
226=>"0000011110111101"&"0010001110011110",
227=>"0010011101111101"&"0010000111111011",
228=>"0001000010100101"&"0010001000001011",
229=>"0000001111110110"&"0010011001100010",
230=>"0001101011010000"&"0010010100101011",
231=>"0000001101110011"&"0010011000001000",
232=>"0001101010000111"&"0001100100100110",
233=>"0000010101101000"&"0010010100100010",
234=>"0001100111101001"&"0010001111100000",
235=>"0001000010010011"&"0001101001001011",
236=>"0010010010000000"&"0001100011100100",
237=>"0000110101100001"&"0010001101111010",
238=>"0001001011010011"&"0010010011010010",
239=>"0010011111000101"&"0001101000001011",
240=>"0000000101100101"&"0010100001000100",
241=>"0000000111010000"&"0010011100011110",
242=>"0001101101000000"&"0010010101000101",
243=>"0001000000000110"&"0010000110000100",
244=>"0010011111110111"&"0010010010001011",
245=>"0001101010001010"&"0010001111111001",
246=>"0001101101110000"&"0001111101100011",
247=>"0010000001111111"&"0010010010110101",
248=>"0000000000011000"&"0010001001100011",
249=>"0001011010100000"&"0001111000101011",
250=>"0000011101100001"&"0010010100100100",
251=>"0001111101100101"&"0001111011010110",
252=>"0001011100001101"&"0010001111001100",
253=>"0001011100101010"&"0010000001010101",
254=>"0001010001110011"&"0001111110001010",
255=>"0000011011011001"&"0001111101010011",
256=>"0000111100010101"&"0001111101000101",
257=>"0001100101011010"&"0010010101111101",
258=>"0001110111010111"&"0010001111011001",
259=>"0001100011100100"&"0010010001101000",
260=>"0011010000111111"&"0001110010110010",
261=>"0001011000001100"&"0010010001000100",
262=>"0000110010001010"&"0010010000111100",
263=>"0000100010000000"&"0010011000001011",
264=>"0001000010000000"&"0010000111001011",
265=>"0001110100010000"&"0010010100101011",
266=>"0010011000000111"&"0010001101000110",
267=>"0001111000001001"&"0010000110101110",
268=>"0010111011010110"&"0010001010010000",
269=>"0000001111110111"&"0010011000000110",
270=>"0001000001000101"&"0001111010101101",
271=>"0000101001111001"&"0010001100011111",
272=>"0000011110011110"&"0010010101101011",
273=>"0000110001111110"&"0010010111010111",
274=>"0001111000101010"&"0010001000110010",
275=>"0001000110101001"&"0010010010111000",
276=>"0000111111011101"&"0010001101100111",
277=>"0000101101100010"&"0001101011000111",
278=>"0001111110101010"&"0010000111000111",
279=>"0001101001010010"&"0010010000111111",
280=>"0010001000110010"&"0010010010111100",
281=>"1111000000110010"&"0001101001100010",
282=>"0000001010011010"&"0001100111100000",
283=>"0010000110010010"&"0001111010011000",
284=>"0000100000011000"&"0010000110000110",
285=>"1111110001111010"&"0001111100011000",
286=>"0001011001110111"&"0010001110010010",
287=>"0001101010011101"&"0010001111010000",
288=>"0000110101110010"&"0001111000001001",
289=>"0011000011100111"&"0010011000011111",
290=>"0010010111110101"&"0001110010111010",
291=>"1111110000011110"&"0001110110000101",
292=>"0000111101011110"&"0010010101000001",
293=>"0010111111000101"&"0010001110010111",
294=>"0001001011011011"&"0001111111011100",
295=>"0001001101010000"&"0001110110101111",
296=>"0001100001000000"&"0010001000001001",
297=>"0001011101110000"&"0010000010101101",
298=>"0000100111110111"&"0010001100000100",
299=>"0001110010100001"&"0010010101010000",
300=>"0000111111011011"&"0010010110001001",
301=>"0010001011111010"&"0001101011001101",
302=>"1110111100001011"&"0001111110111010",
303=>"1111101010011001"&"0010001101100110",
304=>"0011000001101000"&"0010000111110001",
305=>"0001110100100111"&"0001111001011000",
306=>"1111110010011101"&"0010000011011010",
307=>"0001010110100101"&"0010010101101011",
308=>"0001011111010111"&"0010010011000111",
309=>"1111010010111010"&"0001110100001000",
310=>"0000111101111100"&"0010010011001001",
311=>"0001111011111111"&"0010000111111011",
312=>"0001001101001110"&"0010010110011110",
313=>"1111111010110100"&"0010011011111010",
314=>"0000000100001110"&"0001010100100100",
315=>"0001101110011101"&"0010000011001100",
316=>"0000100000110001"&"0001111111000010",
317=>"0000101001010100"&"0010011011011001",
318=>"0000001011010011"&"0010011110111111",
319=>"0001111110001110"&"0001111100111101",
320=>"0001100111110100"&"0001100101010111",
321=>"0000010010011101"&"0010010101100000",
322=>"0001010111100111"&"0001110110100001",
323=>"0000101001100101"&"0001110010111100",
324=>"0000011100101100"&"0001101110001111",
325=>"0000001001111100"&"0001111111111110",
326=>"0001010010000110"&"0010011000100001",
327=>"0010000001110110"&"0010100001010001",
328=>"0001100010111110"&"0010010110011111",
329=>"0001100001110010"&"0010010000111010",
330=>"1101110110101111"&"0010000110001011",
331=>"0001110111101110"&"0010001001110010",
332=>"0010010110110001"&"0010011001110001",
333=>"0001100111100010"&"0010000110001010",
334=>"0010010111000101"&"0010000001100100",
335=>"0000010101100100"&"0010010000000011",
336=>"0001010110100111"&"0010000100101110",
337=>"0001001111110010"&"0010001110010101",
338=>"0010010011001101"&"0010000001100011",
339=>"0010001010000010"&"0010011000011010",
340=>"0010000000100101"&"0010010011111101",
341=>"0000100011010001"&"0001111001001110",
342=>"0001110101100111"&"0010010010100010",
343=>"1111110001111110"&"0010000111000101",
344=>"0001001000011101"&"0010001101001011",
345=>"0001010111010101"&"0001101000011011",
346=>"0010101101100000"&"0001111001001010",
347=>"0001000111010110"&"0010010101000111",
348=>"0010000100000101"&"0010001100010001",
349=>"0001011101010111"&"0001111100001100",
350=>"0001010001011000"&"0001110111100011",
351=>"0000111110001000"&"0010011110111101",
352=>"0001011000001110"&"0010011100101100",
353=>"0010000000101011"&"0010000001100111",
354=>"0001110000010111"&"0010010010000001",
355=>"1111100101110011"&"0010010111000111",
356=>"0001011001101111"&"0001111011101011",
357=>"0001010011011010"&"0010001000111111",
358=>"0000110110010110"&"0001101100110101",
359=>"1111111001000010"&"0001110011010001",
360=>"0001001100001111"&"0001111001010110",
361=>"0001100111100011"&"0001111111001110",
362=>"0000101101111010"&"0001100101011101",
363=>"0000000110010011"&"0010011101000100",
364=>"0001101010110100"&"0010011010000010",
365=>"0000010111100100"&"0001111111100101",
366=>"0001000001000111"&"0010010100101101",
367=>"0001010000011110"&"0010000111111011",
368=>"0010011101011010"&"0001110110110100",
369=>"0001001001111101"&"0010001010111010",
370=>"0010011100000000"&"0010010010111001",
371=>"0001010001110110"&"0010001110100101",
372=>"0000111100111011"&"0010010110110111",
373=>"0001100011101101"&"0010011010110101",
374=>"0010010010000100"&"0010000000011111",
375=>"0001101000000101"&"0001110011111110",
376=>"0001100000001101"&"0010010010100101",
377=>"1111110001010111"&"0010001101111110",
378=>"0001011000111010"&"0010010101000100",
379=>"1110011111101011"&"0001101100010111",
380=>"0001101101100110"&"0010001001101001",
381=>"0000111000000101"&"0010011000101111",
382=>"0000011011010010"&"0001111110110011",
383=>"0000000101011100"&"0010010101110011",
384=>"0000101101111100"&"0010010111110001",
385=>"0000110000001111"&"0010001100010010",
386=>"0000110110101110"&"0001111001010101",
387=>"0001000111101000"&"0010000010010011",
388=>"0000111010001001"&"0010000111011001",
389=>"0010001111011110"&"0010010011001001",
390=>"1111110100100100"&"0001111100101110",
391=>"0001011000110100"&"0001110100111100",
392=>"0001001101101110"&"0001101010111101",
393=>"0000111111000010"&"0010011010101000",
394=>"0000111011000110"&"0010011001111010",
395=>"1101100100011100"&"0001000010000000",
396=>"0001010000101111"&"0010001101011110",
397=>"0001110011011101"&"0010000110000011",
398=>"0010001000010001"&"0010011100000111",
399=>"1111100111011010"&"0010001001000111",
400=>"0001111110011011"&"0001110001100111",
401=>"0000110111101110"&"0010010101001100",
402=>"0001001100010011"&"0010000101110101",
403=>"0001010110001000"&"0010000110110110",
404=>"0000100001101001"&"0010000111010000",
405=>"0001100110010110"&"0010000100001111",
406=>"0001110011110001"&"0010001000111001",
407=>"0001100010101101"&"0010011000100010",
408=>"0000000001110001"&"0001101001111101",
409=>"0010010101010111"&"0010010010111110",
410=>"1111001001100100"&"0001101101100100",
411=>"0001010001010111"&"0001111110000100",
412=>"1111101001001111"&"0001101111101101",
413=>"0001011011111001"&"0010010010101001",
414=>"0010000110000001"&"0010000010011011",
415=>"0001011010100100"&"0010100010101000",
416=>"0001001011010101"&"0010011001110110",
417=>"0000101010101110"&"0010000111111110",
418=>"0010110011111101"&"0010010000001101",
419=>"0000110000010101"&"0010100001011001",
420=>"1110011001101001"&"0001001110010011",
421=>"0010000010111111"&"0010011011011101",
422=>"0010000110001001"&"0010001010111011",
423=>"1111100010101001"&"0001011111111111",
424=>"0001001010001111"&"0010001010110011",
425=>"0001111010111100"&"0010010010000010",
426=>"0001101111100111"&"0010011001010111",
427=>"0000001111101100"&"0010000111011100",
428=>"0001010000100001"&"0010011011110000",
429=>"0000100110011000"&"0010010000111101",
430=>"0011000111000100"&"0010001100010001",
431=>"0010000010110111"&"0010000100010001",
432=>"0000000111010000"&"0010000000101000",
433=>"1111111100000100"&"0010100001001101",
434=>"0000110111000010"&"0001110010110000",
435=>"0010111010001100"&"0010000001110101",
436=>"0000001011011110"&"0010001110010100",
437=>"1111011111010011"&"0010010110101001",
438=>"0000101000101000"&"0010001110110101",
439=>"0000110100101001"&"0010000010111100",
440=>"1111110001111011"&"0001111000001111",
441=>"0000100100111110"&"0001111011110010",
442=>"0001000001000000"&"0010000100001100",
443=>"0001101011111010"&"0010001010010001",
444=>"0001101011110110"&"0001111010000000",
445=>"0000111010000001"&"0010011011111100",
446=>"0010001010001001"&"0010010100110001",
447=>"0001101000101001"&"0001101110101010",
448=>"0000111011010101"&"0010011011010110",
449=>"0000101100110101"&"0010100000101011",
450=>"0001100011111111"&"0010010001100000",
451=>"0001101100011010"&"0010010110110101",
452=>"0001000101000000"&"0010000110100011",
453=>"0001101110100101"&"0010010001101010",
454=>"0000101001111011"&"0010001110111010",
455=>"1111111100001000"&"0010001100101110",
456=>"0010001001010111"&"0010001110010011",
457=>"0000010110001101"&"0010000110011001",
458=>"0001100101100010"&"0010011100111011",
459=>"0000100000111110"&"0010000010110001",
460=>"1110101110011011"&"0001100000110101",
461=>"0010000100100001"&"0001111001110101",
462=>"0000101110101110"&"0001110101110011",
463=>"1111111111101101"&"0001111000110101",
464=>"1111001011011111"&"0010000101110000",
465=>"0001101111011000"&"0010001000110111",
466=>"0010110001000000"&"0010000011010010",
467=>"0001101000111011"&"0010010111001111",
468=>"0000111011010010"&"0001111010000101",
469=>"0001001110100011"&"0010010110010000",
470=>"0000010000000100"&"0010010110100100",
471=>"0000101011100000"&"0010011111011100",
472=>"0001001010111011"&"0001101110001010",
473=>"0000010111100110"&"0010001100011011",
474=>"1111110111000000"&"0001100110001001",
475=>"0000011011010011"&"0001111111001111",
476=>"0001000001111011"&"0010011111011010",
477=>"0001100100000001"&"0010010101001010",
478=>"0000011101101010"&"0010001011011100",
479=>"0000001101011010"&"0010100000101111",
480=>"0001011100011101"&"0010001100001000",
481=>"0001101100110001"&"0010010000010101",
482=>"0001001001110100"&"0001111111011001",
483=>"0000110111011101"&"0001011011100111",
484=>"0000001001100001"&"0001011100010000",
485=>"0000011110100010"&"0010001101100100",
486=>"1111010001111000"&"0010000000010100",
487=>"0011000011011101"&"0001110111001000",
488=>"0000111101011010"&"0010001101000000",
489=>"0000011000001011"&"0001111001111000",
490=>"0000010110000111"&"0001110111101011",
491=>"0001100010000010"&"0010011010010001",
492=>"0000010100000100"&"0001101010110001",
493=>"0000100011111100"&"0010011010001100",
494=>"0010001110101110"&"0010010000101010",
495=>"0001010000010100"&"0010010001000110",
496=>"0001111111110010"&"0001111111100010",
497=>"0001110011110000"&"0010011001110111",
498=>"0001100010010101"&"0010000011100011",
499=>"0001110100000001"&"0010001101111110",
500=>"0001100001110100"&"0010001101111111",
501=>"0001110101000110"&"0010001001110101",
502=>"0000110111100101"&"0010001011011000",
503=>"0000111101000011"&"0010000001110010",
504=>"0010000001111011"&"0010010000101010",
505=>"0001100101011001"&"0010011000011100",
506=>"0000100100011110"&"0001111110001101",
507=>"0001001011100000"&"0010001011011010",
508=>"0001000111000101"&"0001110110110010",
509=>"0001110101100001"&"0010010110110010",
510=>"0001000011001101"&"0010010111100100",
511=>"0001110011001100"&"0010000100000001",
512=>"0001011010001000"&"0001111101101101",
513=>"0001111101000101"&"0010000110011000",
514=>"0010110011111100"&"0010010010011000",
515=>"0010101100111001"&"0010001010100100",
516=>"0001000000001110"&"0010011111000011",
517=>"1100110110001101"&"0001010011000100",
518=>"0000111011110110"&"0010011100110011",
519=>"0001000000110011"&"0001111111110000",
520=>"0000111000001110"&"0001111010111000",
521=>"0001101111001011"&"0010011001010101",
522=>"0000100001100111"&"0001111100100101",
523=>"0010101110111011"&"0001111110101100",
524=>"0010000001001000"&"0010011010100010",
525=>"0001110100111010"&"0010000011001010",
526=>"0000110010111010"&"0010100000001100",
527=>"0000101111000000"&"0010011111110011",
528=>"0000101111111001"&"0010011000100001",
529=>"0001100110100100"&"0010011110111001",
530=>"0000111100101101"&"0010010010011110",
531=>"0001100100000011"&"0010000100110100",
532=>"0001001010100011"&"0010010100011000",
533=>"0000101100001100"&"0001101010011011",
534=>"0001011001000110"&"0010001010101011",
535=>"0000101011000101"&"0010001010001010",
536=>"1111011011101000"&"0010001101100101",
537=>"0001000000001001"&"0010101000101011",
538=>"1111010010111011"&"0001110110101000",
539=>"0000101011011110"&"0001100010100011",
540=>"0001010011000001"&"0001110101000000",
541=>"0001011101110101"&"0010010111101001",
542=>"0001001100010010"&"0010001000110011",
543=>"1111111110110000"&"0010011000101111",
544=>"0001000010001011"&"0010010000111000",
545=>"1111111000110011"&"0001111010000001",
546=>"0010100111010101"&"0010010001111011",
547=>"0001111001001001"&"0010011011000010",
548=>"0000101101010101"&"0010000100000110",
549=>"0001010111111100"&"0010011101000100",
550=>"0000101111101001"&"0001101010110111",
551=>"0001101100110111"&"0010011010011011",
552=>"0000010011110011"&"0010011001111110",
553=>"0010111101000011"&"0010000100000001",
554=>"0000001001110010"&"0010010110010000",
555=>"0000010110100101"&"0010010000100101",
556=>"0001010000111011"&"0010010111100001",
557=>"0001101011010110"&"0010100000000110",
558=>"0000101100100101"&"0010001101110011",
559=>"0010100000010100"&"0010000110111110",
560=>"0001000110110000"&"0010010111101110",
561=>"0000101110000100"&"0010001010110011",
562=>"0001110111010011"&"0001101101100101",
563=>"0010111111011101"&"0001111010101100",
564=>"0000111100101010"&"0010101001101011",
565=>"0000100101010100"&"0010011010101110",
566=>"0010000101010010"&"0010000100101101",
567=>"0001110101101010"&"0010001100011110",
568=>"0001011001011010"&"0010010001111010",
569=>"0000100100100001"&"0001110100001101",
570=>"0001110110100110"&"0001111101000101",
571=>"0010000011011111"&"0010010001001010",
572=>"0000011110110111"&"0001110001110010",
573=>"0000111110011111"&"0010001101110001",
574=>"0000001101100010"&"0001111110010101",
575=>"1111001101110110"&"0001101001011001",
576=>"0010000011000110"&"0010001111011101",
577=>"0000011111000001"&"0010001100011101",
578=>"0010011001000010"&"0010001110000000",
579=>"0010000101010111"&"0010001011010110",
580=>"0001011101000111"&"0010001011001110",
581=>"0000101010010010"&"0010010100110100",
582=>"0000101000100011"&"0010010011010111",
583=>"0001010001010110"&"0010011000010010",
584=>"0001101100001111"&"0010011100011010",
585=>"1101010101001011"&"0001001011111001",
586=>"0000101000010011"&"0010001100000011",
587=>"0000110101101111"&"0010011010100011",
588=>"1101110000011010"&"0001110111111010",
589=>"0001000110101010"&"0010010100100011",
590=>"0001011111100001"&"0010010000110011",
591=>"0000111110110010"&"0010010111001000",
592=>"1110111001011010"&"0001110111111011",
593=>"0001001111100100"&"0010010111010010",
594=>"0001001111111110"&"0010000111101000",
595=>"0001011010110101"&"0001110101101111",
596=>"0001111110000000"&"0010001010000110",
597=>"0001001101100101"&"0010000111111001",
598=>"0010101110110111"&"0010001111100111",
599=>"1110101011110001"&"0001101110000111",
600=>"0000110110001111"&"0010011011110101",
601=>"0010011010011100"&"0010010100011011",
602=>"0010100111010001"&"0001111001101011",
603=>"0000011010111001"&"0010010111101111",
604=>"0000110101110001"&"0010011111001011",
605=>"1110010101101100"&"0001010101101010",
606=>"0000100100001010"&"0010011000010101",
607=>"0000011101000101"&"0001110101001111",
608=>"0000101101101110"&"0010001111001010",
609=>"0001110001101111"&"0010010011001111",
610=>"0001000100000001"&"0010001110100100",
611=>"0000101100101100"&"0010100001110011",
612=>"0010001111000001"&"0010010101111111",
613=>"0001001110011011"&"0010001000110001",
614=>"0010100101101100"&"0001101110111100",
615=>"0001100001110001"&"0010010110000101",
616=>"0001001001100000"&"0010010101000011",
617=>"0001011000010001"&"0010010001000101",
618=>"0001100110111011"&"0001101110110100",
619=>"0001010011101101"&"0010010000011100",
620=>"0010001111010001"&"0010001111100101",
621=>"0001010111110000"&"0010010101001010",
622=>"0001001010011011"&"0010010111101101",
623=>"0000101100110001"&"0010100000100111",
624=>"0010001010111000"&"0010010011101100",
625=>"0001111110110110"&"0010000001111011",
626=>"0001011011001000"&"0010000100110100",
627=>"0000100101000011"&"0010000011011101",
628=>"0001011101011010"&"0001101110110110",
629=>"0000010011100110"&"0001111100000000",
630=>"0000101011010100"&"0010001001001100",
631=>"0000101111110111"&"0010011110110101",
632=>"0001100010000000"&"0010001111101110",
633=>"0000011110001111"&"0001110010111000",
634=>"0010001101110011"&"0010010101110000",
635=>"0001101000111110"&"0010001000001100",
636=>"0010000111000010"&"0001110010100010",
637=>"0011001110110110"&"0010001000100111",
638=>"0000100001001110"&"0010011001000010",
639=>"0000110010100000"&"0001111001010100",
640=>"0010001000010011"&"0010000000100101",
641=>"0001001000101101"&"0001111111110011",
642=>"0000010111111110"&"0010011010100111",
643=>"1111111101011011"&"0010001010010000",
644=>"1111111100010000"&"0010001100110100",
645=>"0001100111110011"&"0010010011001110",
646=>"1111101101111010"&"0010000110101100",
647=>"0001110010011001"&"0010010110101010",
648=>"0001100110100011"&"0010000111000011",
649=>"0000000010110011"&"0001111000000011",
650=>"0001011101100000"&"0010100100111101",
651=>"0000111111101011"&"0010011010010110",
652=>"0001011111101101"&"0001101101001000",
653=>"0001101010011110"&"0001111101001111",
654=>"0010000110101100"&"0010000111100011",
655=>"0001110000110001"&"0010000001001101",
656=>"1111111010111100"&"0001111001111011",
657=>"0001001101001001"&"0010011010011110",
658=>"0010001101100101"&"0010010101001011",
659=>"0010011010111111"&"0001100101111111",
660=>"0001110010001010"&"0010010001110111",
661=>"0000101110110000"&"0010001111111110",
662=>"0010110000101001"&"0001110110011010",
663=>"0000111000110101"&"0010011010000111",
664=>"0010110011001001"&"0010001100000111",
665=>"0001101111000110"&"0010100010100001",
666=>"0001101010000010"&"0010010001010000",
667=>"0001000100010100"&"0001111111111010",
668=>"0010010101110101"&"0010010111011010",
669=>"0001011100111101"&"0010001100010000",
670=>"0001011110000101"&"0010000010001000",
671=>"0000110100110011"&"0001111011110001",
672=>"0010011011011110"&"0001110100110001",
673=>"0001110111111101"&"0010001111010110",
674=>"0000110011000001"&"0010010011001010",
675=>"0000010001001010"&"0010000000000100",
676=>"0010011110111100"&"0010010101001000",
677=>"0001111110101010"&"0010011001011000",
678=>"0001101011100010"&"0010000111110110",
679=>"0000001101010101"&"0010000110111010",
680=>"0001001111010111"&"0010001110000100",
681=>"0001101000110100"&"0010010001011101",
682=>"0001011111001101"&"0010000100111000",
683=>"0000000110001100"&"0001101000101000",
684=>"0000111010000011"&"0001110100101101",
685=>"0001011001101110"&"0010001011000110",
686=>"1111101011011010"&"0001011000100000",
687=>"0010001111100000"&"0010010100100110",
688=>"0000100101000101"&"0010000110101110",
689=>"0000111100000011"&"0010001111111101",
690=>"0001100100111000"&"0010010010001101",
691=>"1111101011001011"&"0001100100001011",
692=>"0010111000111110"&"0010001000111011",
693=>"0000101101110111"&"0010011011011101",
694=>"0010011100101100"&"0010001111011100",
695=>"0001110101111011"&"0010001111000110",
696=>"0010100010011101"&"0010000110101010",
697=>"0011010000000110"&"0001111110111110",
698=>"0000001100101100"&"0001100010010011",
699=>"1111101001111011"&"0001111100111011",
700=>"0000110101001000"&"0010001111101110",
701=>"0000110010101000"&"0010001101111111",
702=>"0001010010100010"&"0010000111001100",
703=>"0000110111010001"&"0001101001000010",
704=>"0001100111010000"&"0001111100001111",
705=>"0001110011001011"&"0010011011010000",
706=>"0010000101110111"&"0010010011000111",
707=>"0000001001010001"&"0001100111111011",
708=>"0000101111010100"&"0010000100000100",
709=>"0001010010101000"&"0010001111000111",
710=>"0001011001010100"&"0010001001001101",
711=>"0010000111101100"&"0010010100101010",
712=>"0000011000010011"&"0010010011100100",
713=>"0000101110010011"&"0010011111110000",
714=>"0001010010010100"&"0010011011110011",
715=>"0000001110110100"&"0010001011001001",
716=>"0001100010000111"&"0010001101100100",
717=>"0010011110001111"&"0010010110000100",
718=>"0010010010001001"&"0001110010111101",
719=>"0001101010100010"&"0010000011011010",
720=>"0001011110000010"&"0001101101111110",
721=>"0001100000110101"&"0010001000100101",
722=>"0010011101101010"&"0010001110111101",
723=>"0000110100111100"&"0010100110010000",
724=>"0001001101000101"&"0010001101101010",
725=>"0000111010000111"&"0010001101101010",
726=>"0000100111001001"&"0001101011110010",
727=>"1111110001100000"&"0001111011000111",
728=>"0001101111100011"&"0010010101100001",
729=>"0000110111110101"&"0010001100001110",
730=>"0001000000000110"&"0010000011011011",
731=>"0000100110000111"&"0010010001101000",
732=>"0001001101001101"&"0010001000001010",
733=>"0001100111101000"&"0001110111001100",
734=>"0001011100111001"&"0010001011010000",
735=>"0000001100000010"&"0010000110111111",
736=>"0010000110111001"&"0010011000100111",
737=>"0001100101100110"&"0010000101111100",
738=>"0000100110111000"&"0010011111000010",
739=>"0000100000010110"&"0010001100001010",
740=>"1111101111100111"&"0001111110000100",
741=>"0001001001110000"&"0010001000111010",
742=>"0000110101011010"&"0010011010111000",
743=>"0001011110001000"&"0010011010010110",
744=>"0010011100011100"&"0001111001110101",
745=>"0000110001110110"&"0010000111011110",
746=>"0001100010000111"&"0010011000101001",
747=>"0010001010100111"&"0010011011011101",
748=>"0010001100100000"&"0001110100111001",
749=>"0000011101101000"&"0010011100101101",
750=>"0000010100000110"&"0010001011101001",
751=>"0000110000011111"&"0010010011101010",
752=>"0000101010101001"&"0010001110101101",
753=>"0010000011011011"&"0010001011000010",
754=>"0000110111111111"&"0010000011000111",
755=>"0001011010010101"&"0001110011001011",
756=>"0001000001100110"&"0010011100011001",
757=>"1111110010111011"&"0010010010110001",
758=>"0001011100100110"&"0001110010110001",
759=>"0001100101111001"&"0010010011101000",
760=>"0000110111111101"&"0010001100100100",
761=>"0000110110100001"&"0010000000101001",
762=>"0001101000100000"&"0001111001000111",
763=>"0001100011000100"&"0010010011011010",
764=>"1111111100001111"&"0001110000011010",
765=>"0010011011111101"&"0010011010110111",
766=>"0001100100001111"&"0010011101110011",
767=>"0010010110000101"&"0001111011010111",
768=>"0000011110000110"&"0010010100110100",
769=>"0001101100011011"&"0010000100011110",
770=>"0000001110100100"&"0001111110000100",
771=>"0010011001100000"&"0010011101001011",
772=>"0000000010101110"&"0010010101011010",
773=>"0010011110110001"&"0001110001110000",
774=>"0001001011000110"&"0001111011110000",
775=>"0001000110111101"&"0010000110010100",
776=>"0000111011011100"&"0010100001010010",
777=>"0001111000100010"&"0010001100101101",
778=>"0010001010011111"&"0010001001111000",
779=>"0010010011100000"&"0010001111101001",
780=>"0001011000011010"&"0010001011100111",
781=>"0000011011010011"&"0010001111010000",
782=>"0000101110010011"&"0010001100101101",
783=>"0010000111100011"&"0001111011110010",
784=>"0001000000011011"&"0010000110110011",
785=>"0001100011110010"&"0010010110101011",
786=>"0010000010100000"&"0010001110100011",
787=>"0001100100001100"&"0010001000010101",
788=>"0000000010110110"&"0001111011110100",
789=>"0000110101111001"&"0010000101101100",
790=>"0000101010100011"&"0010011011111101",
791=>"0001010000000101"&"0010001000101011",
792=>"0001001000010000"&"0010010001100110",
793=>"0001011011100100"&"0010010010010011",
794=>"0000110001101111"&"0010001110111001",
795=>"1111101110110110"&"0010010001101010",
796=>"0010000101110000"&"0010010111010100",
797=>"0000110111101100"&"0010010010000111",
798=>"0000001010001001"&"0010011000110101",
799=>"0001001000111100"&"0001110010110110",
800=>"0000110001000100"&"0010010010101101",
801=>"0001010001001101"&"0010011001101000",
802=>"0001010111100111"&"0001111101011111",
803=>"1111011011001010"&"0001110001000011",
804=>"0001110101011010"&"0010000111010001",
805=>"0001010001110100"&"0010011101001110",
806=>"0001010001000001"&"0010010001000010",
807=>"0000100101101001"&"0010011000010101",
808=>"0001100011101011"&"0010000111100101",
809=>"0000110101010001"&"0010010100011101",
810=>"0001111000101000"&"0010010001101100",
811=>"0000110100000000"&"0010001100101000",
812=>"0010001001011000"&"0010001101011000",
813=>"0000010111010111"&"0001110101110011",
814=>"1111010001100000"&"0010000010100101",
815=>"0001101110110011"&"0010000100100110",
816=>"0001110000010111"&"0010010110010011",
817=>"0010100011100000"&"0010001011110110",
818=>"0000011001001100"&"0010010001101011",
819=>"0000010011001011"&"0010001100101101",
820=>"0001101001101110"&"0001110010101010",
821=>"0001011111111100"&"0010011000100001",
822=>"0001000111101100"&"0001111010100010",
823=>"0001010101010001"&"0010000001001001",
824=>"0001011100000111"&"0010010000111101",
825=>"0001110001100011"&"0001110000100111",
826=>"0001110100101011"&"0010000011101010",
827=>"0000100011100001"&"0010100000110100",
828=>"0001000110110111"&"0010010101110111",
829=>"0000001100111101"&"0001101000101010",
830=>"0010000110100111"&"0010011111111000",
831=>"0001010010110000"&"0001111101100110",
832=>"0001101001010001"&"0010010101101101",
833=>"0001001001001001"&"0010010001111010",
834=>"0001000001010101"&"0001111110110010",
835=>"0001101101110110"&"0010011011110110",
836=>"0001000111100110"&"0010010111101100",
837=>"0000110000100011"&"0001111010011010",
838=>"0000110100011111"&"0010010001101010",
839=>"1111101100101101"&"0010010001000001",
840=>"0000101101101000"&"0010010101101100",
841=>"1111110101000010"&"0001101100010100",
842=>"0001100001011101"&"0010001000000000",
843=>"0010011010100010"&"0010010100011001",
844=>"0010010100010100"&"0001101110101011",
845=>"0010011100111011"&"0010000100101010",
846=>"0010010111001001"&"0010010101111011",
847=>"0001010101001010"&"0010010100110111",
848=>"0010010011111010"&"0010001100000001",
849=>"0001011001111100"&"0001111001000011",
850=>"0010100010110001"&"0010010000101101",
851=>"0000101110110110"&"0010010010110101",
852=>"0001001111001100"&"0001111010110101",
853=>"0000111110101111"&"0001110100001111",
854=>"1111101101101001"&"0001101100101000",
855=>"0001101100110000"&"0010011101111001",
856=>"0001001110110110"&"0010011111100001",
857=>"0001101110101111"&"0010000010011010",
858=>"0010011010110011"&"0001110111111100",
859=>"0001100011010111"&"0010010110110011",
860=>"0001111011110100"&"0001111010001010",
861=>"0001010101100010"&"0010011010011010",
862=>"0000110000101101"&"0010010001001111",
863=>"0000111101110001"&"0010011101011101",
864=>"0001011001111111"&"0010011010011100",
865=>"0000011111011110"&"0010010011010101",
866=>"0000111111001001"&"0010011011101000",
867=>"0000011011101100"&"0010000000011001",
868=>"0010010100111011"&"0010000001110100",
869=>"0000101100101011"&"0001110010000110",
870=>"0000111000111100"&"0010001110011101",
871=>"0001101011110101"&"0010001100110001",
872=>"0000111000011110"&"0010010000111001",
873=>"0010001001111101"&"0010010101011000",
874=>"0010000111000010"&"0001111100010110",
875=>"0000100111011010"&"0010010010110110",
876=>"0010000000001010"&"0001110100110000",
877=>"0000001111110101"&"0010000000100100",
878=>"0001011110010011"&"0010010111011011",
879=>"1111100110010101"&"0010010100001011",
880=>"0000111011111110"&"0010001000100010",
881=>"0001001100111100"&"0010011000110000",
882=>"0001100100111110"&"0001110000110101",
883=>"0000010011101011"&"0010011011110011",
884=>"0001110110101010"&"0001111001000110",
885=>"0000100100100101"&"0010011101100100",
886=>"0001101101001100"&"0010010001011010",
887=>"0001101111010110"&"0010000110100010",
888=>"1110111101101101"&"0010000110100010",
889=>"0010011010100011"&"0010001111010000",
890=>"0001111111101010"&"0010001111101100",
891=>"0001011100110100"&"0001111111001000",
892=>"0000110110100001"&"0010011011010111",
893=>"0001101001101100"&"0010001111000111",
894=>"0000110000010111"&"0010100100001001",
895=>"0000100101000011"&"0010000101101011",
896=>"0010000110101111"&"0001110010000001",
897=>"0000100110101011"&"0010010001100011",
898=>"0001100010100101"&"0001110110001011",
899=>"0001111110100010"&"0010010001011101",
900=>"0010010000011001"&"0010001111101011",
901=>"0010100010110110"&"0010010001111000",
902=>"1111101111001111"&"0010000111101110",
903=>"0001110010010110"&"0010011100111111",
904=>"1111100100110110"&"0010000110000011",
905=>"0001111111110100"&"0010011000010100",
906=>"0001100000100111"&"0001110101001001",
907=>"0001000111110000"&"0010000101000010",
908=>"0000111111101001"&"0010010011110001",
909=>"1110110110111101"&"0001100100101000",
910=>"0000001110011110"&"0010011001111000",
911=>"0001101000011110"&"0001101010111101",
912=>"0001001100010101"&"0001100010100110",
913=>"0000010110000010"&"0010100011100111",
914=>"0000000101000111"&"0010011010101111",
915=>"0001101011110000"&"0001110110001010",
916=>"0000101000110101"&"0010000111000010",
917=>"0000000110100101"&"0010010001010101",
918=>"0001011011000010"&"0001110101110110",
919=>"0001111001111100"&"0010010100100110",
920=>"0000110110101101"&"0010000010110010",
921=>"0000010000101011"&"0010000001100011",
922=>"0001011100010101"&"0010010111100100",
923=>"0001101001110111"&"0010010110111001",
924=>"0001001100000011"&"0010010000010111",
925=>"0000011010110100"&"0010000011101111",
926=>"0000111011001111"&"0010010001000010",
927=>"0001110010011010"&"0001110001111001",
928=>"0001100011000100"&"0010100111100010",
929=>"0001011100000101"&"0001110001010110",
930=>"0000110101111100"&"0010010111001000",
931=>"0010010101111000"&"0001110110100110",
932=>"0001001000010011"&"0001110100010010",
933=>"0000000111001101"&"0001110011110111",
934=>"0000111110110100"&"0010010101110000",
935=>"0000001011100111"&"0010010000100001",
936=>"0001110100011100"&"0001110111111000",
937=>"0001110101001110"&"0010001111100110",
938=>"0000011100011100"&"0010010010110111",
939=>"0010000110010101"&"0001111101110110",
940=>"0001100110000101"&"0010001110011000",
941=>"0001010110010000"&"0010001101001011",
942=>"0010001000011011"&"0010000110111010",
943=>"0001010100100100"&"0010000001001000",
944=>"0011010011000011"&"0010001010001110",
945=>"1111100101010011"&"0001101100010001",
946=>"0001011000100011"&"0010011101100100",
947=>"0001000111010011"&"0010011001010000",
948=>"0001110111010001"&"0001111010101100",
949=>"0000010111100011"&"0010011000111000",
950=>"0000111010100100"&"0010010011001100",
951=>"0010011110011100"&"0010001010000000",
952=>"0001000001111000"&"0010000111110101",
953=>"0001111100100000"&"0001110001101101",
954=>"0001100110001110"&"0001111010000101",
955=>"0000110010111110"&"0001110000000110",
956=>"0001100101011101"&"0010010101100101",
957=>"0000101010100001"&"0010100001001010",
958=>"0001111100110110"&"0001111100011101",
959=>"0001111001111111"&"0010001000001111",
960=>"0000000101001011"&"0010001100101000",
961=>"0001111010010101"&"0010001011111000",
962=>"0001100100110010"&"0010000010011110",
963=>"0000011111001010"&"0010001101101100",
964=>"0000100111101001"&"0001111000011101",
965=>"0010010111010011"&"0010001100010100",
966=>"1111001110110111"&"0010001011011111",
967=>"0001110011111101"&"0001110010110010",
968=>"1111101011100111"&"0010000110000011",
969=>"1111110110111001"&"0010000001000101",
970=>"0001000010001100"&"0010010000110101",
971=>"0001000001001001"&"0010000111000001",
972=>"0000111011111111"&"0010000000100110",
973=>"1111111101100000"&"0010010110001001",
974=>"0001110100010110"&"0010011001110110",
975=>"0000110010011011"&"0001111001110100",
976=>"0000101001100110"&"0001010101110000",
977=>"0001001011011000"&"0010011100000010",
978=>"0000011010110111"&"0010011010100000",
979=>"0001011101011000"&"0010000111011111",
980=>"0001011010111010"&"0010000111110110",
981=>"0001000000110011"&"0010010101010000",
982=>"0001011100111110"&"0010000110000111",
983=>"0001011010111101"&"0010001101111010",
984=>"0010001110001001"&"0001110111100111",
985=>"0000010000001111"&"0010010110100010",
986=>"0001010010100110"&"0010001000000010",
987=>"0010000000100110"&"0010010101000101",
988=>"0000000100000000"&"0001110101001111",
989=>"0000101010111001"&"0010010001011111",
990=>"0001011100101100"&"0001111111101101",
991=>"0001011111100010"&"0010011011000010",
992=>"0010110110101010"&"0010001011110111",
993=>"0001010100010101"&"0010001010101001",
994=>"0011011001011010"&"0010001111111000",
995=>"0010011000000111"&"0001111011011110",
996=>"1110101001100001"&"0001110000111110",
997=>"1101111000010111"&"0001111000010010",
998=>"0000111111001100"&"0010010111010110",
999=>"0001000111100000"&"0010010001000001",
1000=>"0001010111111111"&"0010000001001011",
1001=>"0001101111001101"&"0001111011111001",
1002=>"0010010111001011"&"0010010101000001",
1003=>"0000110110100010"&"0010100100001011",
1004=>"0001101110110010"&"0010000100010101",
1005=>"0001110101111111"&"0010000100110000",
1006=>"0000001111000000"&"0010010000000110",
1007=>"0010010111000001"&"0010001011010110",
1008=>"0000110000111000"&"0001111110101001",
1009=>"0010100000111110"&"0010000101110001",
1010=>"0000101011010101"&"0010010011101000",
1011=>"0010011011101101"&"0010000011000010",
1012=>"0001110100001101"&"0001110111011011",
1013=>"0001111110110110"&"0010001101110101",
1014=>"0010010010011110"&"0010010010110001",
1015=>"0000101110100110"&"0010000010111100",
1016=>"0000111111010000"&"0010001001100100",
1017=>"0000010100101100"&"0001110000100100",
1018=>"0001001011000010"&"0010011001110110",
1019=>"0001110010001001"&"0010001100101100",
1020=>"0001010100011111"&"0010000101011110",
1021=>"0010110011010001"&"0010010010000101",
1022=>"0001000110100000"&"0010010111100010",
1023=>"0001000011011000"&"0001111111011101");
    
BEGIN
    coefs <= ROM_content(to_integer(address));
END RTL;