LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L4WROM IS
    PORT (
        weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
        address : IN unsigned(weightsbitsAddress(4) DOWNTO 0));
END L4WROM;

ARCHITECTURE RTL OF L4WROM IS

    TYPE ROM_mem IS ARRAY (0 TO 8191) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem := (0=>"001001001",
    1=>"111000111",
    2=>"000000000",
    3=>"110100000",
    4=>"110110100",
    5=>"010010110",
    6=>"101001011",
    7=>"100000100",
    8=>"100110100",
    9=>"101101101",
    10=>"011011001",
    11=>"001000100",
    12=>"101101111",
    13=>"000110100",
    14=>"111000001",
    15=>"011001000",
    16=>"101111101",
    17=>"110110110",
    18=>"000000000",
    19=>"000100111",
    20=>"100100100",
    21=>"000001001",
    22=>"010111111",
    23=>"011011011",
    24=>"010111110",
    25=>"100101001",
    26=>"110110111",
    27=>"101000001",
    28=>"011011100",
    29=>"011110100",
    30=>"100100000",
    31=>"001110101",
    32=>"010010010",
    33=>"001011001",
    34=>"011000111",
    35=>"011001010",
    36=>"111100110",
    37=>"001001000",
    38=>"110110100",
    39=>"001001000",
    40=>"011111011",
    41=>"001001001",
    42=>"000100010",
    43=>"000001011",
    44=>"100100100",
    45=>"100000001",
    46=>"000111111",
    47=>"100010111",
    48=>"010110000",
    49=>"110000001",
    50=>"001000011",
    51=>"011110010",
    52=>"001001101",
    53=>"111100000",
    54=>"100100101",
    55=>"111000000",
    56=>"111001011",
    57=>"011001110",
    58=>"100000000",
    59=>"000110000",
    60=>"011011111",
    61=>"100000000",
    62=>"000000000",
    63=>"101001001",
    64=>"111111000",
    65=>"111111111",
    66=>"111111011",
    67=>"100000011",
    68=>"100101101",
    69=>"000000110",
    70=>"001111011",
    71=>"001110100",
    72=>"000000000",
    73=>"000111000",
    74=>"100110000",
    75=>"101111000",
    76=>"101111000",
    77=>"111111111",
    78=>"001101101",
    79=>"000000000",
    80=>"111010010",
    81=>"000000101",
    82=>"000000000",
    83=>"001001001",
    84=>"001000100",
    85=>"000000000",
    86=>"111101111",
    87=>"111000111",
    88=>"110111010",
    89=>"111111111",
    90=>"000000011",
    91=>"111101101",
    92=>"010011111",
    93=>"111111000",
    94=>"110110110",
    95=>"111000011",
    96=>"000000000",
    97=>"010000001",
    98=>"110110110",
    99=>"000000000",
    100=>"001000110",
    101=>"000011001",
    102=>"010000011",
    103=>"000000000",
    104=>"111111111",
    105=>"000000100",
    106=>"101100110",
    107=>"010000011",
    108=>"111111101",
    109=>"110101010",
    110=>"000010111",
    111=>"111111111",
    112=>"011000110",
    113=>"010000010",
    114=>"000000100",
    115=>"100111110",
    116=>"111101111",
    117=>"101101000",
    118=>"101101101",
    119=>"000111101",
    120=>"010000011",
    121=>"110001001",
    122=>"000000000",
    123=>"101111000",
    124=>"000000001",
    125=>"000000000",
    126=>"000000000",
    127=>"111000000",
    128=>"001001001",
    129=>"011111111",
    130=>"111111111",
    131=>"010111110",
    132=>"010110110",
    133=>"000000100",
    134=>"111111111",
    135=>"101101101",
    136=>"011001010",
    137=>"000010000",
    138=>"010011000",
    139=>"111001001",
    140=>"111111111",
    141=>"000000000",
    142=>"111100100",
    143=>"110111110",
    144=>"000000000",
    145=>"010111010",
    146=>"011001100",
    147=>"000000000",
    148=>"000000100",
    149=>"000101000",
    150=>"001000101",
    151=>"000000011",
    152=>"001000001",
    153=>"000110000",
    154=>"000000001",
    155=>"010101000",
    156=>"101000100",
    157=>"010111000",
    158=>"111111111",
    159=>"101101100",
    160=>"001000001",
    161=>"110110011",
    162=>"000000000",
    163=>"001000101",
    164=>"000000000",
    165=>"101101101",
    166=>"010110010",
    167=>"000010000",
    168=>"111111111",
    169=>"000000000",
    170=>"001100100",
    171=>"110110101",
    172=>"000100000",
    173=>"101001001",
    174=>"001001001",
    175=>"010110010",
    176=>"100100110",
    177=>"000000000",
    178=>"000000000",
    179=>"000000000",
    180=>"111111010",
    181=>"101001001",
    182=>"000000001",
    183=>"000101000",
    184=>"110011010",
    185=>"000001000",
    186=>"100101101",
    187=>"100101000",
    188=>"001000101",
    189=>"101000001",
    190=>"010010001",
    191=>"111010000",
    192=>"101011111",
    193=>"100110111",
    194=>"001111001",
    195=>"010110010",
    196=>"110010000",
    197=>"111110000",
    198=>"111001111",
    199=>"100111011",
    200=>"111011000",
    201=>"101101101",
    202=>"011110000",
    203=>"000110110",
    204=>"111111100",
    205=>"000000100",
    206=>"011001001",
    207=>"000110010",
    208=>"111000011",
    209=>"110111010",
    210=>"011111100",
    211=>"100010011",
    212=>"001000000",
    213=>"000000101",
    214=>"101001111",
    215=>"110110000",
    216=>"000000000",
    217=>"011000111",
    218=>"110000001",
    219=>"001001011",
    220=>"000111110",
    221=>"010000110",
    222=>"011110111",
    223=>"001000001",
    224=>"000001100",
    225=>"000110010",
    226=>"000100000",
    227=>"110000000",
    228=>"111101100",
    229=>"000111111",
    230=>"001011010",
    231=>"011111110",
    232=>"101101110",
    233=>"000000111",
    234=>"011000101",
    235=>"111000000",
    236=>"001101101",
    237=>"111111110",
    238=>"101001111",
    239=>"011001001",
    240=>"001000111",
    241=>"000100101",
    242=>"011111110",
    243=>"001001111",
    244=>"000000111",
    245=>"001000101",
    246=>"100010111",
    247=>"000110000",
    248=>"000001011",
    249=>"000100111",
    250=>"111111110",
    251=>"100000000",
    252=>"110110110",
    253=>"000010000",
    254=>"101111100",
    255=>"001000000",
    256=>"001001100",
    257=>"100000000",
    258=>"100100000",
    259=>"011001001",
    260=>"101111111",
    261=>"011001001",
    262=>"110110111",
    263=>"001001000",
    264=>"000000000",
    265=>"100100110",
    266=>"011001000",
    267=>"110110011",
    268=>"001001111",
    269=>"011000001",
    270=>"000010000",
    271=>"100110110",
    272=>"001001000",
    273=>"101101111",
    274=>"100011001",
    275=>"011110001",
    276=>"110011011",
    277=>"100110110",
    278=>"011011001",
    279=>"011001001",
    280=>"011001001",
    281=>"100100110",
    282=>"011001001",
    283=>"001101100",
    284=>"110001101",
    285=>"101100111",
    286=>"111010011",
    287=>"100100100",
    288=>"011011001",
    289=>"001101101",
    290=>"110011001",
    291=>"011001000",
    292=>"010011001",
    293=>"011011001",
    294=>"000101100",
    295=>"100001010",
    296=>"010010010",
    297=>"100100110",
    298=>"000110100",
    299=>"000001000",
    300=>"110010011",
    301=>"011011001",
    302=>"011011001",
    303=>"000010000",
    304=>"100111111",
    305=>"100110111",
    306=>"111011001",
    307=>"100000001",
    308=>"111001100",
    309=>"000001000",
    310=>"111111101",
    311=>"011001001",
    312=>"100010011",
    313=>"100110111",
    314=>"000011001",
    315=>"000011001",
    316=>"011011001",
    317=>"011011001",
    318=>"001110111",
    319=>"000000000",
    320=>"000100011",
    321=>"110000111",
    322=>"111101100",
    323=>"010101111",
    324=>"011000100",
    325=>"001100110",
    326=>"010110010",
    327=>"100101001",
    328=>"011111010",
    329=>"000111001",
    330=>"100000011",
    331=>"001111100",
    332=>"111111111",
    333=>"111111110",
    334=>"001111100",
    335=>"000000001",
    336=>"110010010",
    337=>"110000000",
    338=>"011011101",
    339=>"010000000",
    340=>"001000100",
    341=>"000000001",
    342=>"111000110",
    343=>"110000010",
    344=>"101001001",
    345=>"111010110",
    346=>"110001011",
    347=>"101000011",
    348=>"101101010",
    349=>"001000000",
    350=>"111111111",
    351=>"001000101",
    352=>"101101101",
    353=>"111000100",
    354=>"111000000",
    355=>"100000101",
    356=>"000000110",
    357=>"001101100",
    358=>"101000011",
    359=>"010000101",
    360=>"101111100",
    361=>"000111010",
    362=>"011010111",
    363=>"000000001",
    364=>"100111000",
    365=>"100001011",
    366=>"101101101",
    367=>"100110000",
    368=>"100101000",
    369=>"000000000",
    370=>"011011100",
    371=>"000110100",
    372=>"000110011",
    373=>"000100001",
    374=>"000011011",
    375=>"100000101",
    376=>"110100110",
    377=>"000111100",
    378=>"010110001",
    379=>"000101011",
    380=>"111000111",
    381=>"001001000",
    382=>"111101011",
    383=>"110000000",
    384=>"001001001",
    385=>"000000000",
    386=>"011111010",
    387=>"000110111",
    388=>"001011001",
    389=>"110100100",
    390=>"000000011",
    391=>"100000000",
    392=>"001011001",
    393=>"011111111",
    394=>"100110100",
    395=>"100100100",
    396=>"100111000",
    397=>"110111111",
    398=>"001001101",
    399=>"101111111",
    400=>"111011111",
    401=>"001001001",
    402=>"001000000",
    403=>"000001001",
    404=>"001001100",
    405=>"000010000",
    406=>"111101111",
    407=>"111100111",
    408=>"010011011",
    409=>"010010011",
    410=>"111001011",
    411=>"101101011",
    412=>"000000011",
    413=>"010000010",
    414=>"010000100",
    415=>"000101101",
    416=>"001001001",
    417=>"100110100",
    418=>"110100110",
    419=>"011001111",
    420=>"010111110",
    421=>"001000100",
    422=>"001011011",
    423=>"001000000",
    424=>"000101000",
    425=>"101100100",
    426=>"011001100",
    427=>"110100000",
    428=>"000000100",
    429=>"110110110",
    430=>"000101110",
    431=>"100100001",
    432=>"110110110",
    433=>"010010011",
    434=>"001001010",
    435=>"110110111",
    436=>"000101000",
    437=>"001001001",
    438=>"001100100",
    439=>"010010010",
    440=>"101000011",
    441=>"100100011",
    442=>"100100000",
    443=>"100100100",
    444=>"100100100",
    445=>"101100100",
    446=>"000010010",
    447=>"101001101",
    448=>"000000000",
    449=>"111111111",
    450=>"000000000",
    451=>"111111110",
    452=>"111111111",
    453=>"011100110",
    454=>"100001000",
    455=>"000111000",
    456=>"111111100",
    457=>"000111010",
    458=>"111101111",
    459=>"001001001",
    460=>"000111010",
    461=>"111111011",
    462=>"101000100",
    463=>"000001000",
    464=>"111011000",
    465=>"111111001",
    466=>"000000000",
    467=>"000000000",
    468=>"000000110",
    469=>"000000000",
    470=>"000000010",
    471=>"101111111",
    472=>"011011010",
    473=>"011010000",
    474=>"100110111",
    475=>"010000010",
    476=>"111101111",
    477=>"110111010",
    478=>"011001111",
    479=>"001001010",
    480=>"110000001",
    481=>"111111111",
    482=>"001010111",
    483=>"110110110",
    484=>"000110000",
    485=>"000001101",
    486=>"111111011",
    487=>"000000000",
    488=>"000000000",
    489=>"110110000",
    490=>"011111110",
    491=>"111110011",
    492=>"000000000",
    493=>"100000000",
    494=>"000000001",
    495=>"110000000",
    496=>"110000000",
    497=>"111111111",
    498=>"110000000",
    499=>"011010010",
    500=>"000111111",
    501=>"000000001",
    502=>"000000000",
    503=>"111101111",
    504=>"111011011",
    505=>"000100011",
    506=>"000000000",
    507=>"000000000",
    508=>"001000101",
    509=>"111111111",
    510=>"000000000",
    511=>"111001101",
    512=>"000100100",
    513=>"110100100",
    514=>"011011010",
    515=>"111111101",
    516=>"001001000",
    517=>"010010000",
    518=>"000100111",
    519=>"001001011",
    520=>"011011011",
    521=>"011011011",
    522=>"011011011",
    523=>"001001100",
    524=>"101101101",
    525=>"001110110",
    526=>"010011100",
    527=>"011011001",
    528=>"001110100",
    529=>"110110110",
    530=>"000010110",
    531=>"000000000",
    532=>"000001100",
    533=>"000100101",
    534=>"100100100",
    535=>"110100101",
    536=>"100100100",
    537=>"100100100",
    538=>"100101111",
    539=>"001011111",
    540=>"100110100",
    541=>"111001001",
    542=>"110110010",
    543=>"001001100",
    544=>"011011011",
    545=>"001001001",
    546=>"011011001",
    547=>"001000000",
    548=>"001011000",
    549=>"010001001",
    550=>"010011111",
    551=>"100110110",
    552=>"001011011",
    553=>"000010100",
    554=>"110110001",
    555=>"010110110",
    556=>"000100101",
    557=>"000111101",
    558=>"001001011",
    559=>"101100100",
    560=>"010101100",
    561=>"000000000",
    562=>"111111001",
    563=>"001000100",
    564=>"000100000",
    565=>"000001000",
    566=>"101011101",
    567=>"011011010",
    568=>"100100100",
    569=>"001001000",
    570=>"110100100",
    571=>"000001000",
    572=>"100100100",
    573=>"111100000",
    574=>"001001000",
    575=>"101001001",
    576=>"000100100",
    577=>"001001001",
    578=>"001000110",
    579=>"100110110",
    580=>"000011111",
    581=>"100100110",
    582=>"011011001",
    583=>"000110011",
    584=>"000111101",
    585=>"000100111",
    586=>"010111011",
    587=>"001000111",
    588=>"001101101",
    589=>"100010011",
    590=>"001001111",
    591=>"110111010",
    592=>"100010001",
    593=>"111011000",
    594=>"011001100",
    595=>"011011001",
    596=>"000000101",
    597=>"000011000",
    598=>"111011000",
    599=>"010011000",
    600=>"001001101",
    601=>"011001101",
    602=>"011011000",
    603=>"000011000",
    604=>"011010000",
    605=>"001000111",
    606=>"000100100",
    607=>"100000110",
    608=>"011010011",
    609=>"101101111",
    610=>"001000100",
    611=>"000000111",
    612=>"101110001",
    613=>"001000111",
    614=>"010011001",
    615=>"111001001",
    616=>"000100111",
    617=>"000000000",
    618=>"001101100",
    619=>"111001001",
    620=>"100010001",
    621=>"100110000",
    622=>"100110111",
    623=>"100010011",
    624=>"110010001",
    625=>"111011011",
    626=>"101001101",
    627=>"100011001",
    628=>"000011011",
    629=>"100111110",
    630=>"100100101",
    631=>"110011001",
    632=>"110011001",
    633=>"000110110",
    634=>"100111011",
    635=>"100110111",
    636=>"110011000",
    637=>"000011001",
    638=>"100110111",
    639=>"011011000",
    640=>"000100101",
    641=>"011010110",
    642=>"011101011",
    643=>"000101111",
    644=>"000110111",
    645=>"011000100",
    646=>"100000000",
    647=>"000110101",
    648=>"011001000",
    649=>"010110011",
    650=>"010010110",
    651=>"010000000",
    652=>"111110010",
    653=>"111000101",
    654=>"110000000",
    655=>"010111000",
    656=>"000000101",
    657=>"010110000",
    658=>"100110110",
    659=>"010101101",
    660=>"001000100",
    661=>"000000000",
    662=>"100000011",
    663=>"001100000",
    664=>"100100111",
    665=>"111000011",
    666=>"101001001",
    667=>"111100000",
    668=>"100000011",
    669=>"000010000",
    670=>"000000000",
    671=>"000000000",
    672=>"000000111",
    673=>"111011000",
    674=>"000111111",
    675=>"100000000",
    676=>"000000111",
    677=>"100100101",
    678=>"011010000",
    679=>"111111111",
    680=>"000111111",
    681=>"110000011",
    682=>"100111101",
    683=>"100000000",
    684=>"001100111",
    685=>"111010100",
    686=>"101000111",
    687=>"111100101",
    688=>"111111111",
    689=>"100100000",
    690=>"110100100",
    691=>"110111010",
    692=>"000000011",
    693=>"101001101",
    694=>"001100101",
    695=>"111111000",
    696=>"100001000",
    697=>"011001110",
    698=>"000001001",
    699=>"000000100",
    700=>"010100000",
    701=>"001010001",
    702=>"011111001",
    703=>"100100111",
    704=>"111001000",
    705=>"000100101",
    706=>"111000000",
    707=>"111110010",
    708=>"100110001",
    709=>"000110001",
    710=>"011000001",
    711=>"111001100",
    712=>"000100111",
    713=>"111011000",
    714=>"001011100",
    715=>"100111001",
    716=>"111101110",
    717=>"000101110",
    718=>"000110011",
    719=>"010000111",
    720=>"001100110",
    721=>"000110111",
    722=>"000000111",
    723=>"001000100",
    724=>"100011001",
    725=>"000110011",
    726=>"000110111",
    727=>"100110001",
    728=>"011101000",
    729=>"000110001",
    730=>"011100100",
    731=>"111011000",
    732=>"000000111",
    733=>"011100011",
    734=>"100111000",
    735=>"100110001",
    736=>"110001100",
    737=>"000110111",
    738=>"100111001",
    739=>"001000100",
    740=>"000110001",
    741=>"011000111",
    742=>"011001000",
    743=>"000100011",
    744=>"111001000",
    745=>"111010001",
    746=>"100111011",
    747=>"100100000",
    748=>"111000000",
    749=>"101100000",
    750=>"111001100",
    751=>"000010011",
    752=>"111100111",
    753=>"000000110",
    754=>"000100011",
    755=>"000110111",
    756=>"111110110",
    757=>"111010000",
    758=>"100110001",
    759=>"111011001",
    760=>"100110001",
    761=>"111001001",
    762=>"100011100",
    763=>"111000000",
    764=>"000110111",
    765=>"010011111",
    766=>"111111001",
    767=>"000100011",
    768=>"000000001",
    769=>"000000000",
    770=>"000000000",
    771=>"000111000",
    772=>"111111011",
    773=>"100011001",
    774=>"100001100",
    775=>"001011010",
    776=>"111111111",
    777=>"100010010",
    778=>"111111110",
    779=>"100011001",
    780=>"010111010",
    781=>"000000000",
    782=>"001111011",
    783=>"111111111",
    784=>"000000000",
    785=>"111111111",
    786=>"111101111",
    787=>"000011101",
    788=>"111101111",
    789=>"010011000",
    790=>"000000000",
    791=>"001001011",
    792=>"000000000",
    793=>"000000100",
    794=>"001111100",
    795=>"010011100",
    796=>"011011010",
    797=>"100001001",
    798=>"100000000",
    799=>"000000000",
    800=>"111111111",
    801=>"100110011",
    802=>"000000000",
    803=>"100000110",
    804=>"111111111",
    805=>"100110001",
    806=>"011111100",
    807=>"111111111",
    808=>"000000000",
    809=>"000000000",
    810=>"100011001",
    811=>"000000010",
    812=>"000000000",
    813=>"011010100",
    814=>"111111111",
    815=>"000000000",
    816=>"010111000",
    817=>"010111101",
    818=>"100010000",
    819=>"010100010",
    820=>"110110100",
    821=>"011011110",
    822=>"000000010",
    823=>"100101101",
    824=>"101011111",
    825=>"011110000",
    826=>"111101111",
    827=>"111011110",
    828=>"111111111",
    829=>"010000001",
    830=>"111110111",
    831=>"000111011",
    832=>"010111000",
    833=>"000010000",
    834=>"011010000",
    835=>"010111010",
    836=>"000111100",
    837=>"011111010",
    838=>"000111010",
    839=>"100111001",
    840=>"011011010",
    841=>"000111000",
    842=>"010011010",
    843=>"000011010",
    844=>"111111111",
    845=>"100001110",
    846=>"000111000",
    847=>"010111010",
    848=>"010010010",
    849=>"010011010",
    850=>"001011110",
    851=>"010110000",
    852=>"011111000",
    853=>"010010010",
    854=>"101001101",
    855=>"010111010",
    856=>"001000001",
    857=>"010011000",
    858=>"110111000",
    859=>"010011010",
    860=>"010010010",
    861=>"000000000",
    862=>"000111010",
    863=>"010111010",
    864=>"010111010",
    865=>"010110010",
    866=>"111011000",
    867=>"101100100",
    868=>"010111010",
    869=>"010111110",
    870=>"010110010",
    871=>"011010010",
    872=>"000111000",
    873=>"010111010",
    874=>"010011010",
    875=>"000000011",
    876=>"000111000",
    877=>"110111010",
    878=>"111101100",
    879=>"001111011",
    880=>"000111010",
    881=>"010011010",
    882=>"111111010",
    883=>"000011010",
    884=>"010011010",
    885=>"000110000",
    886=>"010111010",
    887=>"001100000",
    888=>"010010000",
    889=>"010111000",
    890=>"000011010",
    891=>"010110010",
    892=>"000101001",
    893=>"101101001",
    894=>"110010010",
    895=>"010000000",
    896=>"011111001",
    897=>"110110100",
    898=>"011011000",
    899=>"001011111",
    900=>"001001000",
    901=>"100100100",
    902=>"100110100",
    903=>"001011011",
    904=>"111111110",
    905=>"000101111",
    906=>"001011111",
    907=>"111100000",
    908=>"001001111",
    909=>"010000000",
    910=>"111100000",
    911=>"111011000",
    912=>"100100100",
    913=>"001001111",
    914=>"110111001",
    915=>"000100100",
    916=>"111100100",
    917=>"110100100",
    918=>"100001111",
    919=>"100100100",
    920=>"101100001",
    921=>"001001011",
    922=>"000010110",
    923=>"000100111",
    924=>"110100100",
    925=>"001001011",
    926=>"110110100",
    927=>"110100000",
    928=>"100000010",
    929=>"011000000",
    930=>"000100000",
    931=>"011000001",
    932=>"000010100",
    933=>"111011001",
    934=>"110001111",
    935=>"110110000",
    936=>"011110100",
    937=>"110110100",
    938=>"010100001",
    939=>"001110110",
    940=>"111000100",
    941=>"000110110",
    942=>"011001011",
    943=>"000000000",
    944=>"001001011",
    945=>"110100000",
    946=>"110100100",
    947=>"000100000",
    948=>"100100100",
    949=>"000001001",
    950=>"011111100",
    951=>"111011110",
    952=>"100100110",
    953=>"101101001",
    954=>"101011000",
    955=>"011011011",
    956=>"111001110",
    957=>"101001011",
    958=>"001110110",
    959=>"110110000",
    960=>"100000000",
    961=>"101101101",
    962=>"011101011",
    963=>"001111100",
    964=>"000000000",
    965=>"010100001",
    966=>"111111011",
    967=>"000000000",
    968=>"111000001",
    969=>"111111001",
    970=>"001111111",
    971=>"100000001",
    972=>"111101101",
    973=>"110111111",
    974=>"100000000",
    975=>"000000010",
    976=>"000101011",
    977=>"000111100",
    978=>"000000000",
    979=>"011101111",
    980=>"000000000",
    981=>"110000001",
    982=>"100111111",
    983=>"011111111",
    984=>"110100001",
    985=>"110100011",
    986=>"001111110",
    987=>"101111111",
    988=>"101101111",
    989=>"001111110",
    990=>"110100001",
    991=>"110000001",
    992=>"111001001",
    993=>"010000001",
    994=>"100000001",
    995=>"000000001",
    996=>"001001001",
    997=>"100000000",
    998=>"101111111",
    999=>"110100111",
    1000=>"110000011",
    1001=>"110000000",
    1002=>"100000101",
    1003=>"011110101",
    1004=>"100000000",
    1005=>"101110101",
    1006=>"100000001",
    1007=>"010011111",
    1008=>"000001110",
    1009=>"100001110",
    1010=>"000000000",
    1011=>"111111111",
    1012=>"100111111",
    1013=>"110000001",
    1014=>"111000011",
    1015=>"110000000",
    1016=>"110111111",
    1017=>"000000101",
    1018=>"000000001",
    1019=>"111111011",
    1020=>"000000000",
    1021=>"000000001",
    1022=>"111010100",
    1023=>"101000001",
    1024=>"000110110",
    1025=>"010000000",
    1026=>"111111111",
    1027=>"111111010",
    1028=>"000100110",
    1029=>"110111111",
    1030=>"000000000",
    1031=>"000000000",
    1032=>"111100110",
    1033=>"111110010",
    1034=>"111111010",
    1035=>"100111111",
    1036=>"110111010",
    1037=>"010000110",
    1038=>"001000110",
    1039=>"000000000",
    1040=>"001111011",
    1041=>"000111011",
    1042=>"011000000",
    1043=>"000000000",
    1044=>"011100110",
    1045=>"000000000",
    1046=>"101001011",
    1047=>"011001011",
    1048=>"011101111",
    1049=>"000111011",
    1050=>"000000000",
    1051=>"010001000",
    1052=>"001011001",
    1053=>"100010000",
    1054=>"111111111",
    1055=>"111111011",
    1056=>"011001000",
    1057=>"001001000",
    1058=>"010011111",
    1059=>"000000100",
    1060=>"111101111",
    1061=>"111111111",
    1062=>"010111111",
    1063=>"001000000",
    1064=>"001111101",
    1065=>"000000000",
    1066=>"110111101",
    1067=>"000000001",
    1068=>"000000100",
    1069=>"000010000",
    1070=>"111001100",
    1071=>"111111111",
    1072=>"000000101",
    1073=>"000001001",
    1074=>"111111011",
    1075=>"000000011",
    1076=>"000100000",
    1077=>"000000111",
    1078=>"010010001",
    1079=>"011000100",
    1080=>"001001000",
    1081=>"010111010",
    1082=>"000100101",
    1083=>"011101100",
    1084=>"001000000",
    1085=>"111111111",
    1086=>"000000000",
    1087=>"000110111",
    1088=>"111011000",
    1089=>"000001100",
    1090=>"011111111",
    1091=>"000000101",
    1092=>"000010110",
    1093=>"110011000",
    1094=>"101001011",
    1095=>"010010110",
    1096=>"000011011",
    1097=>"101001000",
    1098=>"010000000",
    1099=>"010011001",
    1100=>"111111110",
    1101=>"000100110",
    1102=>"000100110",
    1103=>"000000001",
    1104=>"100110010",
    1105=>"000000000",
    1106=>"101101101",
    1107=>"010110000",
    1108=>"111101111",
    1109=>"000000000",
    1110=>"111101010",
    1111=>"001111011",
    1112=>"000110111",
    1113=>"000000010",
    1114=>"111110011",
    1115=>"001000111",
    1116=>"101000000",
    1117=>"110110010",
    1118=>"001101011",
    1119=>"001101111",
    1120=>"110110010",
    1121=>"000011010",
    1122=>"111111111",
    1123=>"010110000",
    1124=>"111110000",
    1125=>"110110110",
    1126=>"000010000",
    1127=>"011000110",
    1128=>"101101111",
    1129=>"000000000",
    1130=>"110011000",
    1131=>"001101001",
    1132=>"100111011",
    1133=>"110110100",
    1134=>"010010010",
    1135=>"001001111",
    1136=>"100100000",
    1137=>"000000011",
    1138=>"100111111",
    1139=>"111111011",
    1140=>"111111111",
    1141=>"110001011",
    1142=>"100100110",
    1143=>"000000000",
    1144=>"111011000",
    1145=>"001100000",
    1146=>"111101101",
    1147=>"011101111",
    1148=>"010110010",
    1149=>"100100001",
    1150=>"000100001",
    1151=>"111000001",
    1152=>"111000000",
    1153=>"100001111",
    1154=>"111111101",
    1155=>"011011011",
    1156=>"010000000",
    1157=>"110011001",
    1158=>"111111101",
    1159=>"000010110",
    1160=>"110110011",
    1161=>"100001111",
    1162=>"000011011",
    1163=>"011011111",
    1164=>"101101100",
    1165=>"111001101",
    1166=>"011011011",
    1167=>"001101100",
    1168=>"010000001",
    1169=>"111101111",
    1170=>"000010001",
    1171=>"001011011",
    1172=>"011001001",
    1173=>"001001000",
    1174=>"100100100",
    1175=>"100110001",
    1176=>"100100110",
    1177=>"001011111",
    1178=>"111101110",
    1179=>"011011000",
    1180=>"000110000",
    1181=>"100100000",
    1182=>"110001001",
    1183=>"110000010",
    1184=>"100110100",
    1185=>"111111011",
    1186=>"001100110",
    1187=>"110110000",
    1188=>"100100000",
    1189=>"110110110",
    1190=>"100100010",
    1191=>"011010100",
    1192=>"000001000",
    1193=>"111011011",
    1194=>"011011011",
    1195=>"000100110",
    1196=>"000011011",
    1197=>"000000000",
    1198=>"001100110",
    1199=>"001101111",
    1200=>"100100010",
    1201=>"010011001",
    1202=>"100100110",
    1203=>"111110111",
    1204=>"110110011",
    1205=>"111111111",
    1206=>"011000000",
    1207=>"011000000",
    1208=>"001001110",
    1209=>"001011000",
    1210=>"000000000",
    1211=>"000000000",
    1212=>"000100100",
    1213=>"100100000",
    1214=>"011011010",
    1215=>"001001001",
    1216=>"110100100",
    1217=>"011011111",
    1218=>"000011111",
    1219=>"110100100",
    1220=>"010100100",
    1221=>"001001000",
    1222=>"011111110",
    1223=>"110110100",
    1224=>"000010000",
    1225=>"001011011",
    1226=>"110110111",
    1227=>"100001100",
    1228=>"101100101",
    1229=>"111010000",
    1230=>"000000110",
    1231=>"001011111",
    1232=>"111110000",
    1233=>"001011011",
    1234=>"000000100",
    1235=>"101100100",
    1236=>"100000000",
    1237=>"000001001",
    1238=>"111110100",
    1239=>"111001000",
    1240=>"111100000",
    1241=>"001011111",
    1242=>"110100000",
    1243=>"111111110",
    1244=>"010100001",
    1245=>"001011011",
    1246=>"010011011",
    1247=>"000100001",
    1248=>"110100100",
    1249=>"000011001",
    1250=>"001001000",
    1251=>"110100000",
    1252=>"001001001",
    1253=>"001100110",
    1254=>"011110100",
    1255=>"000001101",
    1256=>"000010111",
    1257=>"000011011",
    1258=>"000001001",
    1259=>"001010000",
    1260=>"100110110",
    1261=>"110110100",
    1262=>"110100100",
    1263=>"111111111",
    1264=>"111011001",
    1265=>"001010011",
    1266=>"101000100",
    1267=>"111100101",
    1268=>"001001101",
    1269=>"110110100",
    1270=>"100000000",
    1271=>"111100100",
    1272=>"011111000",
    1273=>"000111111",
    1274=>"111100100",
    1275=>"110100100",
    1276=>"111100000",
    1277=>"100000000",
    1278=>"000010101",
    1279=>"110100100",
    1280=>"100100011",
    1281=>"111011111",
    1282=>"010111001",
    1283=>"000000000",
    1284=>"001011000",
    1285=>"111111111",
    1286=>"011011011",
    1287=>"001000111",
    1288=>"000001000",
    1289=>"101001001",
    1290=>"110110010",
    1291=>"101000000",
    1292=>"000000011",
    1293=>"001011000",
    1294=>"111000100",
    1295=>"111011111",
    1296=>"000000111",
    1297=>"101000000",
    1298=>"011000100",
    1299=>"111011111",
    1300=>"001100100",
    1301=>"100000000",
    1302=>"000000000",
    1303=>"111100001",
    1304=>"000000000",
    1305=>"111011000",
    1306=>"011011001",
    1307=>"101100100",
    1308=>"011010000",
    1309=>"111111111",
    1310=>"111001111",
    1311=>"111110000",
    1312=>"100111011",
    1313=>"000010010",
    1314=>"111111000",
    1315=>"010001111",
    1316=>"101100010",
    1317=>"010011111",
    1318=>"011110101",
    1319=>"111111100",
    1320=>"101111111",
    1321=>"100000000",
    1322=>"111001111",
    1323=>"111111101",
    1324=>"101001111",
    1325=>"110000000",
    1326=>"000000001",
    1327=>"101111011",
    1328=>"100000000",
    1329=>"111011000",
    1330=>"000000001",
    1331=>"010110010",
    1332=>"000000000",
    1333=>"110100001",
    1334=>"110111111",
    1335=>"000111111",
    1336=>"110000000",
    1337=>"111001100",
    1338=>"100000000",
    1339=>"110100001",
    1340=>"001010010",
    1341=>"000101001",
    1342=>"111100101",
    1343=>"110100100",
    1344=>"000010010",
    1345=>"000000000",
    1346=>"001100100",
    1347=>"111101111",
    1348=>"100110100",
    1349=>"011010110",
    1350=>"000000000",
    1351=>"100100101",
    1352=>"000111110",
    1353=>"001101111",
    1354=>"100101011",
    1355=>"001111110",
    1356=>"000111111",
    1357=>"001111000",
    1358=>"000001101",
    1359=>"110101101",
    1360=>"111111000",
    1361=>"111000010",
    1362=>"000010010",
    1363=>"100000010",
    1364=>"010111000",
    1365=>"111111111",
    1366=>"111111111",
    1367=>"011111000",
    1368=>"111111110",
    1369=>"110101111",
    1370=>"110111011",
    1371=>"110100010",
    1372=>"010010010",
    1373=>"001101101",
    1374=>"010000010",
    1375=>"111111110",
    1376=>"011111011",
    1377=>"011011000",
    1378=>"000111010",
    1379=>"100010000",
    1380=>"000000000",
    1381=>"001111111",
    1382=>"110110000",
    1383=>"010110000",
    1384=>"011011101",
    1385=>"000000000",
    1386=>"000010001",
    1387=>"110001000",
    1388=>"100000000",
    1389=>"110000000",
    1390=>"111111111",
    1391=>"110110110",
    1392=>"011110110",
    1393=>"000101111",
    1394=>"011011011",
    1395=>"110111100",
    1396=>"110000000",
    1397=>"100111010",
    1398=>"011011001",
    1399=>"111111111",
    1400=>"100000010",
    1401=>"000110100",
    1402=>"010110100",
    1403=>"010110000",
    1404=>"110111010",
    1405=>"101000000",
    1406=>"100000010",
    1407=>"011111111",
    1408=>"000100001",
    1409=>"000000000",
    1410=>"000001100",
    1411=>"101101101",
    1412=>"000000000",
    1413=>"110111111",
    1414=>"101111111",
    1415=>"111111001",
    1416=>"000000101",
    1417=>"010111011",
    1418=>"000000000",
    1419=>"011111100",
    1420=>"000111011",
    1421=>"111111111",
    1422=>"000101100",
    1423=>"011010011",
    1424=>"111111110",
    1425=>"111110010",
    1426=>"111110101",
    1427=>"000010001",
    1428=>"111100100",
    1429=>"000100000",
    1430=>"000000010",
    1431=>"010000111",
    1432=>"000111000",
    1433=>"100111000",
    1434=>"111111111",
    1435=>"110001111",
    1436=>"111111110",
    1437=>"001111111",
    1438=>"000101010",
    1439=>"000000010",
    1440=>"011111111",
    1441=>"000000000",
    1442=>"111010000",
    1443=>"001000100",
    1444=>"010000111",
    1445=>"010111101",
    1446=>"000000000",
    1447=>"011101111",
    1448=>"101101000",
    1449=>"111111111",
    1450=>"011011001",
    1451=>"110000101",
    1452=>"000100110",
    1453=>"010101111",
    1454=>"110111111",
    1455=>"111111000",
    1456=>"000000000",
    1457=>"001000000",
    1458=>"111011000",
    1459=>"000010100",
    1460=>"111101101",
    1461=>"000001000",
    1462=>"111111011",
    1463=>"111111111",
    1464=>"110010010",
    1465=>"111101100",
    1466=>"111011111",
    1467=>"111111001",
    1468=>"000011011",
    1469=>"100000000",
    1470=>"001011001",
    1471=>"000000000",
    1472=>"111000000",
    1473=>"110000011",
    1474=>"111000000",
    1475=>"111000000",
    1476=>"111110000",
    1477=>"110111000",
    1478=>"111010000",
    1479=>"000000111",
    1480=>"111010101",
    1481=>"000001111",
    1482=>"111000001",
    1483=>"111100000",
    1484=>"111001111",
    1485=>"011111001",
    1486=>"111000000",
    1487=>"111000111",
    1488=>"111101001",
    1489=>"000111111",
    1490=>"110100000",
    1491=>"110001001",
    1492=>"001100100",
    1493=>"111000000",
    1494=>"001111111",
    1495=>"000010010",
    1496=>"001001111",
    1497=>"001111111",
    1498=>"001111110",
    1499=>"010001000",
    1500=>"011010100",
    1501=>"000111111",
    1502=>"111011000",
    1503=>"011010101",
    1504=>"110000001",
    1505=>"111000100",
    1506=>"111010010",
    1507=>"001100111",
    1508=>"011110100",
    1509=>"110000000",
    1510=>"001001010",
    1511=>"111010000",
    1512=>"111000000",
    1513=>"011000000",
    1514=>"111100100",
    1515=>"000011011",
    1516=>"011000000",
    1517=>"111011000",
    1518=>"100000111",
    1519=>"000000010",
    1520=>"100000111",
    1521=>"100000010",
    1522=>"100000001",
    1523=>"111010000",
    1524=>"111001000",
    1525=>"111011000",
    1526=>"111000000",
    1527=>"010000000",
    1528=>"000111011",
    1529=>"011000001",
    1530=>"011001000",
    1531=>"111001000",
    1532=>"001111110",
    1533=>"000000011",
    1534=>"111000000",
    1535=>"110111001",
    1536=>"101111110",
    1537=>"110111100",
    1538=>"000000000",
    1539=>"110110100",
    1540=>"000011111",
    1541=>"101101000",
    1542=>"100110010",
    1543=>"000011111",
    1544=>"011000000",
    1545=>"000110110",
    1546=>"111110110",
    1547=>"000000010",
    1548=>"101111111",
    1549=>"100100000",
    1550=>"000000001",
    1551=>"110100111",
    1552=>"100001110",
    1553=>"001101000",
    1554=>"010110110",
    1555=>"010011110",
    1556=>"000000000",
    1557=>"000010000",
    1558=>"011001001",
    1559=>"000001100",
    1560=>"000011011",
    1561=>"011110110",
    1562=>"001001000",
    1563=>"001011001",
    1564=>"000001001",
    1565=>"100100110",
    1566=>"001110111",
    1567=>"001011011",
    1568=>"000011001",
    1569=>"001001011",
    1570=>"111011011",
    1571=>"001001001",
    1572=>"111111011",
    1573=>"000111011",
    1574=>"011001000",
    1575=>"000101011",
    1576=>"111111110",
    1577=>"100100100",
    1578=>"110111110",
    1579=>"100101001",
    1580=>"110011111",
    1581=>"011011111",
    1582=>"000001001",
    1583=>"110110100",
    1584=>"001001011",
    1585=>"001100100",
    1586=>"000100111",
    1587=>"111111101",
    1588=>"001100100",
    1589=>"000000000",
    1590=>"111111011",
    1591=>"001001000",
    1592=>"100100001",
    1593=>"010000000",
    1594=>"001011011",
    1595=>"111111011",
    1596=>"001011011",
    1597=>"100001001",
    1598=>"001001010",
    1599=>"110110110",
    1600=>"001010110",
    1601=>"110010001",
    1602=>"111110000",
    1603=>"110101011",
    1604=>"101000000",
    1605=>"110100001",
    1606=>"101011100",
    1607=>"101001010",
    1608=>"111100000",
    1609=>"100100001",
    1610=>"000001111",
    1611=>"111100000",
    1612=>"101111101",
    1613=>"000110000",
    1614=>"100001000",
    1615=>"001011111",
    1616=>"100101001",
    1617=>"000011111",
    1618=>"001111001",
    1619=>"001011110",
    1620=>"110110000",
    1621=>"000001010",
    1622=>"010011110",
    1623=>"001011110",
    1624=>"110100000",
    1625=>"001011100",
    1626=>"001011110",
    1627=>"001110100",
    1628=>"001001011",
    1629=>"110100000",
    1630=>"110100110",
    1631=>"001011110",
    1632=>"011110101",
    1633=>"110010000",
    1634=>"100110100",
    1635=>"000000001",
    1636=>"000010111",
    1637=>"111110000",
    1638=>"000001011",
    1639=>"010111100",
    1640=>"111100000",
    1641=>"100001110",
    1642=>"001110100",
    1643=>"010101110",
    1644=>"101001000",
    1645=>"001011110",
    1646=>"111100001",
    1647=>"101101110",
    1648=>"111110000",
    1649=>"001010100",
    1650=>"011110001",
    1651=>"100010100",
    1652=>"100001101",
    1653=>"001010110",
    1654=>"001011110",
    1655=>"111110100",
    1656=>"001011110",
    1657=>"011111100",
    1658=>"011011010",
    1659=>"001011110",
    1660=>"001011111",
    1661=>"111100001",
    1662=>"001010110",
    1663=>"000001111",
    1664=>"011001001",
    1665=>"110111111",
    1666=>"001001001",
    1667=>"001001101",
    1668=>"001001001",
    1669=>"011000100",
    1670=>"101001011",
    1671=>"000000000",
    1672=>"011001101",
    1673=>"110110110",
    1674=>"101001001",
    1675=>"011001001",
    1676=>"101101100",
    1677=>"100110011",
    1678=>"011001001",
    1679=>"101000010",
    1680=>"100000000",
    1681=>"110110110",
    1682=>"011001001",
    1683=>"001011111",
    1684=>"001001000",
    1685=>"001001001",
    1686=>"110110110",
    1687=>"101100110",
    1688=>"110110010",
    1689=>"000100000",
    1690=>"110110110",
    1691=>"001111011",
    1692=>"001101001",
    1693=>"110110110",
    1694=>"001001001",
    1695=>"001001001",
    1696=>"001001001",
    1697=>"011001001",
    1698=>"111100010",
    1699=>"110110110",
    1700=>"011000100",
    1701=>"000001001",
    1702=>"100111011",
    1703=>"011001000",
    1704=>"001001001",
    1705=>"100100100",
    1706=>"111001001",
    1707=>"110110110",
    1708=>"001001001",
    1709=>"001001011",
    1710=>"011001001",
    1711=>"001001001",
    1712=>"111111110",
    1713=>"100101111",
    1714=>"010011011",
    1715=>"001001011",
    1716=>"001001001",
    1717=>"011001001",
    1718=>"001001001",
    1719=>"101101101",
    1720=>"100100110",
    1721=>"011011000",
    1722=>"001000000",
    1723=>"001001011",
    1724=>"001000000",
    1725=>"100100100",
    1726=>"001001011",
    1727=>"001001101",
    1728=>"000111011",
    1729=>"001001001",
    1730=>"111001000",
    1731=>"101000111",
    1732=>"111011011",
    1733=>"111001100",
    1734=>"101100100",
    1735=>"100111011",
    1736=>"110011001",
    1737=>"111010000",
    1738=>"000010111",
    1739=>"111001000",
    1740=>"111110010",
    1741=>"000110001",
    1742=>"010011001",
    1743=>"100100111",
    1744=>"000001000",
    1745=>"001100111",
    1746=>"011000000",
    1747=>"001100100",
    1748=>"010001000",
    1749=>"110000000",
    1750=>"001001111",
    1751=>"101100100",
    1752=>"111001000",
    1753=>"001100111",
    1754=>"100110111",
    1755=>"110100011",
    1756=>"111100100",
    1757=>"011001001",
    1758=>"010001101",
    1759=>"101100000",
    1760=>"110110010",
    1761=>"011100110",
    1762=>"010101000",
    1763=>"111001100",
    1764=>"110111110",
    1765=>"111001000",
    1766=>"000100000",
    1767=>"100100000",
    1768=>"111011001",
    1769=>"000100111",
    1770=>"011001000",
    1771=>"001000100",
    1772=>"011001000",
    1773=>"100110111",
    1774=>"111011011",
    1775=>"011000000",
    1776=>"001101101",
    1777=>"101100101",
    1778=>"011011000",
    1779=>"000000001",
    1780=>"100100110",
    1781=>"000111011",
    1782=>"100110011",
    1783=>"100100010",
    1784=>"001100110",
    1785=>"011111101",
    1786=>"000110011",
    1787=>"110111111",
    1788=>"001100111",
    1789=>"001000000",
    1790=>"100111111",
    1791=>"010010000",
    1792=>"100100101",
    1793=>"100111111",
    1794=>"001011011",
    1795=>"101101101",
    1796=>"000101110",
    1797=>"011100011",
    1798=>"000000010",
    1799=>"110000100",
    1800=>"001011011",
    1801=>"000001000",
    1802=>"010110111",
    1803=>"001000010",
    1804=>"111100111",
    1805=>"010011111",
    1806=>"110000100",
    1807=>"000000000",
    1808=>"111000000",
    1809=>"111100000",
    1810=>"100000000",
    1811=>"111011011",
    1812=>"111100110",
    1813=>"101011011",
    1814=>"011101111",
    1815=>"000010011",
    1816=>"000000000",
    1817=>"011010000",
    1818=>"111100011",
    1819=>"101000001",
    1820=>"011011010",
    1821=>"000001011",
    1822=>"100000000",
    1823=>"011001000",
    1824=>"111000111",
    1825=>"001000010",
    1826=>"111010010",
    1827=>"001100010",
    1828=>"111111110",
    1829=>"111001000",
    1830=>"011011011",
    1831=>"000101100",
    1832=>"000011000",
    1833=>"111100100",
    1834=>"111000100",
    1835=>"000100001",
    1836=>"101100100",
    1837=>"010011000",
    1838=>"111100101",
    1839=>"110110100",
    1840=>"010011010",
    1841=>"000011000",
    1842=>"111101100",
    1843=>"111110101",
    1844=>"000011001",
    1845=>"001001001",
    1846=>"101101100",
    1847=>"100100011",
    1848=>"111100111",
    1849=>"100001101",
    1850=>"110100000",
    1851=>"011100000",
    1852=>"111100100",
    1853=>"011100101",
    1854=>"100100101",
    1855=>"100000000",
    1856=>"000000010",
    1857=>"001001000",
    1858=>"110110110",
    1859=>"110100110",
    1860=>"100100100",
    1861=>"001001001",
    1862=>"000100000",
    1863=>"110000000",
    1864=>"110000100",
    1865=>"110100000",
    1866=>"110100100",
    1867=>"000000000",
    1868=>"101111001",
    1869=>"000100001",
    1870=>"110111111",
    1871=>"011101100",
    1872=>"001101000",
    1873=>"101101101",
    1874=>"000111011",
    1875=>"111010100",
    1876=>"101101110",
    1877=>"110110100",
    1878=>"011011111",
    1879=>"100000001",
    1880=>"001001011",
    1881=>"110100000",
    1882=>"001001000",
    1883=>"111110110",
    1884=>"110100100",
    1885=>"101001111",
    1886=>"111100010",
    1887=>"110100100",
    1888=>"001011011",
    1889=>"100110110",
    1890=>"111101001",
    1891=>"001001001",
    1892=>"000000000",
    1893=>"100100100",
    1894=>"110101001",
    1895=>"100110000",
    1896=>"000010010",
    1897=>"100100100",
    1898=>"101011011",
    1899=>"011111100",
    1900=>"100000100",
    1901=>"111100110",
    1902=>"001011111",
    1903=>"000001000",
    1904=>"111100100",
    1905=>"000001000",
    1906=>"001111111",
    1907=>"000000000",
    1908=>"000001011",
    1909=>"110110001",
    1910=>"111111110",
    1911=>"001001001",
    1912=>"011110100",
    1913=>"000000000",
    1914=>"101001101",
    1915=>"000000000",
    1916=>"001001111",
    1917=>"001011011",
    1918=>"110110110",
    1919=>"011011011",
    1920=>"001101010",
    1921=>"000100111",
    1922=>"111111110",
    1923=>"100111000",
    1924=>"000000101",
    1925=>"100001011",
    1926=>"000100110",
    1927=>"001001110",
    1928=>"111111001",
    1929=>"011010000",
    1930=>"100100110",
    1931=>"011110010",
    1932=>"101101100",
    1933=>"101100000",
    1934=>"000111001",
    1935=>"101001001",
    1936=>"101100100",
    1937=>"111011001",
    1938=>"000000001",
    1939=>"100110101",
    1940=>"111110101",
    1941=>"000000100",
    1942=>"100001100",
    1943=>"100100100",
    1944=>"001000100",
    1945=>"011001011",
    1946=>"100100100",
    1947=>"000100100",
    1948=>"000100110",
    1949=>"011011001",
    1950=>"100100110",
    1951=>"000100100",
    1952=>"100100100",
    1953=>"110111111",
    1954=>"001000000",
    1955=>"001000000",
    1956=>"000110001",
    1957=>"000011011",
    1958=>"100100110",
    1959=>"100110000",
    1960=>"101010111",
    1961=>"101111111",
    1962=>"100110000",
    1963=>"001100100",
    1964=>"011011010",
    1965=>"000100101",
    1966=>"100011110",
    1967=>"100100100",
    1968=>"001101001",
    1969=>"100001001",
    1970=>"100110011",
    1971=>"101111111",
    1972=>"100101101",
    1973=>"000111111",
    1974=>"000110011",
    1975=>"000100100",
    1976=>"100100100",
    1977=>"100101101",
    1978=>"100110111",
    1979=>"000000100",
    1980=>"010001100",
    1981=>"001100001",
    1982=>"100100110",
    1983=>"000000000",
    1984=>"110111111",
    1985=>"000111010",
    1986=>"000111000",
    1987=>"011010000",
    1988=>"000111111",
    1989=>"000000000",
    1990=>"000111000",
    1991=>"100100111",
    1992=>"000111111",
    1993=>"011101000",
    1994=>"000111111",
    1995=>"100000110",
    1996=>"000100111",
    1997=>"000011111",
    1998=>"011101101",
    1999=>"111000000",
    2000=>"000000000",
    2001=>"000000110",
    2002=>"001000000",
    2003=>"111000000",
    2004=>"000000100",
    2005=>"111100000",
    2006=>"111111111",
    2007=>"010000000",
    2008=>"000010000",
    2009=>"110000110",
    2010=>"100100000",
    2011=>"000011111",
    2012=>"111010000",
    2013=>"111001001",
    2014=>"000011000",
    2015=>"111010000",
    2016=>"000000000",
    2017=>"111000000",
    2018=>"011111100",
    2019=>"000000111",
    2020=>"111100111",
    2021=>"000000011",
    2022=>"111011000",
    2023=>"010101000",
    2024=>"100000000",
    2025=>"100000111",
    2026=>"100100001",
    2027=>"000010111",
    2028=>"101111111",
    2029=>"000100000",
    2030=>"111111000",
    2031=>"000000010",
    2032=>"000010111",
    2033=>"000111010",
    2034=>"011000000",
    2035=>"100010000",
    2036=>"000011011",
    2037=>"110001000",
    2038=>"001111111",
    2039=>"110111101",
    2040=>"000010010",
    2041=>"000101111",
    2042=>"010000010",
    2043=>"011010000",
    2044=>"000000000",
    2045=>"110000000",
    2046=>"110011000",
    2047=>"111000000",
    2048=>"100100100",
    2049=>"000010011",
    2050=>"001011111",
    2051=>"011000010",
    2052=>"011100000",
    2053=>"011100010",
    2054=>"001001011",
    2055=>"110110100",
    2056=>"011001000",
    2057=>"111101101",
    2058=>"110000110",
    2059=>"011001101",
    2060=>"111101000",
    2061=>"001001111",
    2062=>"011101101",
    2063=>"111000000",
    2064=>"111000100",
    2065=>"101000111",
    2066=>"011011001",
    2067=>"011001001",
    2068=>"001001000",
    2069=>"010000001",
    2070=>"001010111",
    2071=>"110100010",
    2072=>"000011011",
    2073=>"000111111",
    2074=>"110111010",
    2075=>"110000110",
    2076=>"001000001",
    2077=>"001011011",
    2078=>"100100110",
    2079=>"011000000",
    2080=>"111111000",
    2081=>"001001100",
    2082=>"000100010",
    2083=>"000100010",
    2084=>"110110100",
    2085=>"011011001",
    2086=>"100100101",
    2087=>"011011001",
    2088=>"100110101",
    2089=>"010100000",
    2090=>"011011001",
    2091=>"101000011",
    2092=>"001001001",
    2093=>"100100100",
    2094=>"111101000",
    2095=>"000001011",
    2096=>"111000001",
    2097=>"001101001",
    2098=>"011010101",
    2099=>"111101000",
    2100=>"111000100",
    2101=>"110100100",
    2102=>"010000101",
    2103=>"011001010",
    2104=>"110100111",
    2105=>"111000001",
    2106=>"110110100",
    2107=>"100100000",
    2108=>"101001010",
    2109=>"011001000",
    2110=>"110100100",
    2111=>"000000001",
    2112=>"110100100",
    2113=>"001011111",
    2114=>"011011111",
    2115=>"011011111",
    2116=>"011011111",
    2117=>"100001001",
    2118=>"011100101",
    2119=>"010100000",
    2120=>"001011111",
    2121=>"100100100",
    2122=>"001011111",
    2123=>"110100000",
    2124=>"101001111",
    2125=>"010000000",
    2126=>"110110000",
    2127=>"010010011",
    2128=>"101110001",
    2129=>"001011001",
    2130=>"100100100",
    2131=>"011100111",
    2132=>"110110000",
    2133=>"100100100",
    2134=>"110100000",
    2135=>"110001001",
    2136=>"011011011",
    2137=>"110100000",
    2138=>"110100000",
    2139=>"110100001",
    2140=>"100000000",
    2141=>"000000100",
    2142=>"111011011",
    2143=>"100100100",
    2144=>"100100000",
    2145=>"011111101",
    2146=>"111010100",
    2147=>"100000000",
    2148=>"110100100",
    2149=>"100100110",
    2150=>"011111111",
    2151=>"101100101",
    2152=>"011011111",
    2153=>"110100000",
    2154=>"110000000",
    2155=>"100100001",
    2156=>"100100101",
    2157=>"100100100",
    2158=>"100100100",
    2159=>"100000000",
    2160=>"101011111",
    2161=>"110000000",
    2162=>"100111010",
    2163=>"101101001",
    2164=>"001011111",
    2165=>"100100000",
    2166=>"110111001",
    2167=>"001001111",
    2168=>"100001011",
    2169=>"100100110",
    2170=>"010100000",
    2171=>"100100100",
    2172=>"011010001",
    2173=>"110100011",
    2174=>"011111011",
    2175=>"000100100",
    2176=>"011001000",
    2177=>"011011000",
    2178=>"100100110",
    2179=>"001111111",
    2180=>"100100110",
    2181=>"101100011",
    2182=>"111110111",
    2183=>"011001101",
    2184=>"100100110",
    2185=>"101111111",
    2186=>"101110001",
    2187=>"100110011",
    2188=>"101101111",
    2189=>"010010001",
    2190=>"100110010",
    2191=>"000100111",
    2192=>"011001001",
    2193=>"011001101",
    2194=>"100110010",
    2195=>"110010111",
    2196=>"110010011",
    2197=>"100100010",
    2198=>"011011101",
    2199=>"111011000",
    2200=>"111001001",
    2201=>"111001010",
    2202=>"011001101",
    2203=>"110000001",
    2204=>"100100110",
    2205=>"000100011",
    2206=>"001001001",
    2207=>"100010010",
    2208=>"100100110",
    2209=>"100100110",
    2210=>"100000011",
    2211=>"001001101",
    2212=>"000101101",
    2213=>"100100010",
    2214=>"011001001",
    2215=>"100110010",
    2216=>"000000010",
    2217=>"001000001",
    2218=>"110110011",
    2219=>"010011001",
    2220=>"100110010",
    2221=>"000000011",
    2222=>"100110110",
    2223=>"100110110",
    2224=>"011011001",
    2225=>"000010011",
    2226=>"001100010",
    2227=>"101110011",
    2228=>"111001001",
    2229=>"101000000",
    2230=>"100010110",
    2231=>"011001001",
    2232=>"101110010",
    2233=>"100110011",
    2234=>"011101101",
    2235=>"100000000",
    2236=>"110011101",
    2237=>"010000100",
    2238=>"001001001",
    2239=>"000100110",
    2240=>"000010100",
    2241=>"010101101",
    2242=>"111101111",
    2243=>"111010010",
    2244=>"100100001",
    2245=>"110100000",
    2246=>"101111110",
    2247=>"011101110",
    2248=>"000000000",
    2249=>"011000011",
    2250=>"001001000",
    2251=>"111111011",
    2252=>"111111111",
    2253=>"001001000",
    2254=>"011011110",
    2255=>"110111110",
    2256=>"000011110",
    2257=>"111101110",
    2258=>"111111111",
    2259=>"110111110",
    2260=>"000000000",
    2261=>"100111111",
    2262=>"000111000",
    2263=>"001011000",
    2264=>"000000101",
    2265=>"101011110",
    2266=>"001000000",
    2267=>"010110001",
    2268=>"000010001",
    2269=>"110000100",
    2270=>"111110111",
    2271=>"010010001",
    2272=>"111110100",
    2273=>"011110110",
    2274=>"111111111",
    2275=>"000000000",
    2276=>"011000000",
    2277=>"110100011",
    2278=>"110111011",
    2279=>"100111011",
    2280=>"110010101",
    2281=>"000000000",
    2282=>"100111010",
    2283=>"111111110",
    2284=>"111110111",
    2285=>"001000000",
    2286=>"111101000",
    2287=>"110110000",
    2288=>"010010001",
    2289=>"000000000",
    2290=>"101101011",
    2291=>"001001010",
    2292=>"011111111",
    2293=>"001111110",
    2294=>"111010101",
    2295=>"100000010",
    2296=>"111110110",
    2297=>"001011110",
    2298=>"100011110",
    2299=>"100000010",
    2300=>"000001001",
    2301=>"000000011",
    2302=>"111110110",
    2303=>"000000010",
    2304=>"110000001",
    2305=>"000111111",
    2306=>"000111111",
    2307=>"000111111",
    2308=>"001111111",
    2309=>"111101000",
    2310=>"001001011",
    2311=>"001100001",
    2312=>"010111111",
    2313=>"111000000",
    2314=>"100111111",
    2315=>"000001111",
    2316=>"111111110",
    2317=>"101000011",
    2318=>"111100000",
    2319=>"001101110",
    2320=>"111001000",
    2321=>"111110110",
    2322=>"111001010",
    2323=>"111111000",
    2324=>"001000110",
    2325=>"000101001",
    2326=>"000000101",
    2327=>"100100111",
    2328=>"000000000",
    2329=>"001000111",
    2330=>"111100001",
    2331=>"011001001",
    2332=>"010110110",
    2333=>"010011111",
    2334=>"010000110",
    2335=>"101101101",
    2336=>"100000000",
    2337=>"010111111",
    2338=>"111001101",
    2339=>"110000000",
    2340=>"001000000",
    2341=>"100000001",
    2342=>"110111111",
    2343=>"110111111",
    2344=>"000111111",
    2345=>"111000000",
    2346=>"111000000",
    2347=>"101100000",
    2348=>"011001101",
    2349=>"011100111",
    2350=>"000010111",
    2351=>"111011111",
    2352=>"000011111",
    2353=>"000000111",
    2354=>"100001110",
    2355=>"001000000",
    2356=>"000111111",
    2357=>"000001101",
    2358=>"111100001",
    2359=>"000010000",
    2360=>"111111000",
    2361=>"001000001",
    2362=>"111100100",
    2363=>"111101111",
    2364=>"001001001",
    2365=>"001001001",
    2366=>"110111111",
    2367=>"110001001",
    2368=>"010100100",
    2369=>"010010000",
    2370=>"011111100",
    2371=>"101101111",
    2372=>"010001011",
    2373=>"000010110",
    2374=>"111111111",
    2375=>"000001000",
    2376=>"011000010",
    2377=>"111011001",
    2378=>"010000001",
    2379=>"110010100",
    2380=>"111111011",
    2381=>"001011000",
    2382=>"001011000",
    2383=>"011111010",
    2384=>"010111011",
    2385=>"011001000",
    2386=>"001110000",
    2387=>"000001001",
    2388=>"111100100",
    2389=>"100000010",
    2390=>"010000010",
    2391=>"011001000",
    2392=>"110000000",
    2393=>"011111010",
    2394=>"100000001",
    2395=>"110110111",
    2396=>"111111111",
    2397=>"001100010",
    2398=>"111111111",
    2399=>"000000000",
    2400=>"000000000",
    2401=>"010010101",
    2402=>"001011101",
    2403=>"101100100",
    2404=>"001110100",
    2405=>"001111000",
    2406=>"000000001",
    2407=>"111110000",
    2408=>"111101000",
    2409=>"000000011",
    2410=>"000011001",
    2411=>"000001100",
    2412=>"000001000",
    2413=>"000011000",
    2414=>"111111101",
    2415=>"000101010",
    2416=>"100100101",
    2417=>"100101111",
    2418=>"010010000",
    2419=>"000000000",
    2420=>"000000000",
    2421=>"110100101",
    2422=>"001111111",
    2423=>"010010000",
    2424=>"010011110",
    2425=>"111001000",
    2426=>"110111000",
    2427=>"111111001",
    2428=>"010000000",
    2429=>"111000001",
    2430=>"111100011",
    2431=>"100000111",
    2432=>"111111011",
    2433=>"011000111",
    2434=>"000000000",
    2435=>"001100110",
    2436=>"000000110",
    2437=>"000111110",
    2438=>"110011001",
    2439=>"100010000",
    2440=>"010000000",
    2441=>"111001001",
    2442=>"000000000",
    2443=>"110110000",
    2444=>"111111100",
    2445=>"101011000",
    2446=>"011100100",
    2447=>"100111000",
    2448=>"111111111",
    2449=>"000000111",
    2450=>"010111010",
    2451=>"010010001",
    2452=>"001100111",
    2453=>"000000000",
    2454=>"000110110",
    2455=>"000000111",
    2456=>"000000101",
    2457=>"000000110",
    2458=>"000011011",
    2459=>"101100001",
    2460=>"111000100",
    2461=>"000000000",
    2462=>"011110111",
    2463=>"001000001",
    2464=>"011111000",
    2465=>"100110111",
    2466=>"111000111",
    2467=>"000000000",
    2468=>"110111110",
    2469=>"100111100",
    2470=>"001011111",
    2471=>"010000000",
    2472=>"000000000",
    2473=>"111001000",
    2474=>"111100111",
    2475=>"011011011",
    2476=>"111111101",
    2477=>"011000010",
    2478=>"100111000",
    2479=>"110111011",
    2480=>"000110111",
    2481=>"000000000",
    2482=>"001000000",
    2483=>"100000000",
    2484=>"000000111",
    2485=>"001111000",
    2486=>"001111000",
    2487=>"111111000",
    2488=>"001011011",
    2489=>"111011101",
    2490=>"001111010",
    2491=>"100000000",
    2492=>"000000111",
    2493=>"100111111",
    2494=>"000000000",
    2495=>"000000000",
    2496=>"001001000",
    2497=>"000000000",
    2498=>"111111011",
    2499=>"010010000",
    2500=>"111111111",
    2501=>"100000100",
    2502=>"000000000",
    2503=>"000111010",
    2504=>"111100111",
    2505=>"010111010",
    2506=>"111111101",
    2507=>"110111101",
    2508=>"110111010",
    2509=>"000100001",
    2510=>"111101101",
    2511=>"111001111",
    2512=>"000000000",
    2513=>"000000000",
    2514=>"011101100",
    2515=>"100000101",
    2516=>"000101000",
    2517=>"100100101",
    2518=>"100111000",
    2519=>"100000000",
    2520=>"000000000",
    2521=>"011001101",
    2522=>"001001000",
    2523=>"100001111",
    2524=>"111111000",
    2525=>"011111011",
    2526=>"000000000",
    2527=>"111111101",
    2528=>"000101101",
    2529=>"011011100",
    2530=>"000000000",
    2531=>"101000100",
    2532=>"111111111",
    2533=>"011111010",
    2534=>"000111011",
    2535=>"011110110",
    2536=>"101111110",
    2537=>"000000000",
    2538=>"110000100",
    2539=>"100000000",
    2540=>"000000001",
    2541=>"001101001",
    2542=>"111111111",
    2543=>"010101111",
    2544=>"100100111",
    2545=>"100101001",
    2546=>"000000010",
    2547=>"000101001",
    2548=>"101111111",
    2549=>"111111011",
    2550=>"111001111",
    2551=>"001100100",
    2552=>"000001001",
    2553=>"001100001",
    2554=>"110100000",
    2555=>"100011101",
    2556=>"000000000",
    2557=>"100000001",
    2558=>"111111111",
    2559=>"101101000",
    2560=>"111111100",
    2561=>"000010000",
    2562=>"000000111",
    2563=>"000000111",
    2564=>"000000000",
    2565=>"110111001",
    2566=>"000111100",
    2567=>"001001111",
    2568=>"110111111",
    2569=>"110001100",
    2570=>"001011000",
    2571=>"110010000",
    2572=>"111000111",
    2573=>"000000000",
    2574=>"000010101",
    2575=>"000000111",
    2576=>"111110000",
    2577=>"010111111",
    2578=>"010101000",
    2579=>"101011010",
    2580=>"111011000",
    2581=>"011000000",
    2582=>"011011101",
    2583=>"000011000",
    2584=>"111010000",
    2585=>"010011000",
    2586=>"001111100",
    2587=>"111001000",
    2588=>"000110010",
    2589=>"111100011",
    2590=>"010011001",
    2591=>"000111111",
    2592=>"011101010",
    2593=>"000110111",
    2594=>"000000000",
    2595=>"011000110",
    2596=>"111111111",
    2597=>"111000011",
    2598=>"000001111",
    2599=>"111110000",
    2600=>"111000110",
    2601=>"111000001",
    2602=>"111111000",
    2603=>"000000000",
    2604=>"110110001",
    2605=>"111111000",
    2606=>"111000000",
    2607=>"010110010",
    2608=>"000111110",
    2609=>"111111000",
    2610=>"100110011",
    2611=>"101110000",
    2612=>"101110111",
    2613=>"100000000",
    2614=>"001000110",
    2615=>"011111000",
    2616=>"000010001",
    2617=>"010000111",
    2618=>"011111000",
    2619=>"001111100",
    2620=>"000010000",
    2621=>"110000011",
    2622=>"111010111",
    2623=>"111111000",
    2624=>"101000010",
    2625=>"001110000",
    2626=>"110111011",
    2627=>"111110000",
    2628=>"000000011",
    2629=>"100100001",
    2630=>"110011010",
    2631=>"011010010",
    2632=>"000001011",
    2633=>"110100101",
    2634=>"000011111",
    2635=>"001000010",
    2636=>"111111010",
    2637=>"100111101",
    2638=>"000001010",
    2639=>"110110000",
    2640=>"101001010",
    2641=>"010111100",
    2642=>"011001000",
    2643=>"000000011",
    2644=>"111100000",
    2645=>"000001111",
    2646=>"100000110",
    2647=>"001011111",
    2648=>"100100011",
    2649=>"101001110",
    2650=>"101000000",
    2651=>"010001001",
    2652=>"000001111",
    2653=>"111100000",
    2654=>"101000101",
    2655=>"000000000",
    2656=>"001000111",
    2657=>"000101111",
    2658=>"101111111",
    2659=>"111000000",
    2660=>"111110000",
    2661=>"111110100",
    2662=>"111001001",
    2663=>"000011111",
    2664=>"001001001",
    2665=>"000000011",
    2666=>"000000011",
    2667=>"110111001",
    2668=>"000000011",
    2669=>"000000001",
    2670=>"011111000",
    2671=>"111000111",
    2672=>"011111110",
    2673=>"000001111",
    2674=>"010110100",
    2675=>"001011111",
    2676=>"011011010",
    2677=>"100001111",
    2678=>"010000001",
    2679=>"000100111",
    2680=>"101001001",
    2681=>"001000110",
    2682=>"000100000",
    2683=>"011000000",
    2684=>"110100101",
    2685=>"110100000",
    2686=>"000001011",
    2687=>"000000011",
    2688=>"001001010",
    2689=>"100100000",
    2690=>"010011111",
    2691=>"001010010",
    2692=>"011111111",
    2693=>"101001101",
    2694=>"110110100",
    2695=>"011011110",
    2696=>"000011000",
    2697=>"011010010",
    2698=>"111110111",
    2699=>"001001011",
    2700=>"101111111",
    2701=>"111010000",
    2702=>"001011011",
    2703=>"011110100",
    2704=>"010110001",
    2705=>"110100100",
    2706=>"000000001",
    2707=>"010110101",
    2708=>"101111010",
    2709=>"001000000",
    2710=>"111101001",
    2711=>"110100100",
    2712=>"100001011",
    2713=>"100101111",
    2714=>"110100100",
    2715=>"010100000",
    2716=>"100100101",
    2717=>"011011001",
    2718=>"000001001",
    2719=>"101001001",
    2720=>"001011110",
    2721=>"000001001",
    2722=>"100001101",
    2723=>"100110000",
    2724=>"010101111",
    2725=>"001001011",
    2726=>"110100100",
    2727=>"000000000",
    2728=>"001011011",
    2729=>"100100100",
    2730=>"100001111",
    2731=>"100100000",
    2732=>"001001111",
    2733=>"010101111",
    2734=>"011011010",
    2735=>"011111011",
    2736=>"110100100",
    2737=>"110100000",
    2738=>"001001101",
    2739=>"000000000",
    2740=>"110110000",
    2741=>"000010110",
    2742=>"011010110",
    2743=>"000001001",
    2744=>"110100100",
    2745=>"001111011",
    2746=>"001011110",
    2747=>"001011110",
    2748=>"100100101",
    2749=>"100001100",
    2750=>"000011110",
    2751=>"010001001",
    2752=>"101101100",
    2753=>"101100100",
    2754=>"110001000",
    2755=>"001011011",
    2756=>"101101111",
    2757=>"100000100",
    2758=>"110010110",
    2759=>"011101101",
    2760=>"111110110",
    2761=>"010000000",
    2762=>"101101111",
    2763=>"111111110",
    2764=>"101101101",
    2765=>"101011010",
    2766=>"000000000",
    2767=>"101110100",
    2768=>"001000000",
    2769=>"111111111",
    2770=>"010001001",
    2771=>"111000110",
    2772=>"100010100",
    2773=>"100100000",
    2774=>"011011101",
    2775=>"111110110",
    2776=>"100001000",
    2777=>"001001011",
    2778=>"101010100",
    2779=>"111111111",
    2780=>"001011011",
    2781=>"011111111",
    2782=>"100000011",
    2783=>"100100100",
    2784=>"011001100",
    2785=>"101101101",
    2786=>"000011000",
    2787=>"000001011",
    2788=>"001010000",
    2789=>"100000001",
    2790=>"100101000",
    2791=>"110110110",
    2792=>"010110000",
    2793=>"011011111",
    2794=>"111011110",
    2795=>"001011001",
    2796=>"111111101",
    2797=>"000000000",
    2798=>"001000101",
    2799=>"001011010",
    2800=>"001001001",
    2801=>"001011000",
    2802=>"101110011",
    2803=>"000111000",
    2804=>"100100100",
    2805=>"111111111",
    2806=>"111001101",
    2807=>"001001001",
    2808=>"100000000",
    2809=>"000000000",
    2810=>"110010000",
    2811=>"111111111",
    2812=>"100101110",
    2813=>"000001011",
    2814=>"011110101",
    2815=>"000000010",
    2816=>"010001000",
    2817=>"111011000",
    2818=>"110010001",
    2819=>"100111111",
    2820=>"011000100",
    2821=>"000011101",
    2822=>"000110001",
    2823=>"011100000",
    2824=>"101110101",
    2825=>"111000000",
    2826=>"111101000",
    2827=>"111000100",
    2828=>"101101111",
    2829=>"011110011",
    2830=>"111000000",
    2831=>"011010000",
    2832=>"001110010",
    2833=>"010100111",
    2834=>"000100111",
    2835=>"001011101",
    2836=>"100001101",
    2837=>"111001000",
    2838=>"100111111",
    2839=>"011000000",
    2840=>"000001100",
    2841=>"000000101",
    2842=>"001001000",
    2843=>"111111111",
    2844=>"100000000",
    2845=>"111011011",
    2846=>"100010011",
    2847=>"111101011",
    2848=>"111001000",
    2849=>"011001100",
    2850=>"111011111",
    2851=>"001100101",
    2852=>"101110011",
    2853=>"001100000",
    2854=>"011001000",
    2855=>"101110010",
    2856=>"010000010",
    2857=>"000010110",
    2858=>"000000000",
    2859=>"000100100",
    2860=>"010111011",
    2861=>"111000000",
    2862=>"111111001",
    2863=>"111110110",
    2864=>"000100111",
    2865=>"111001000",
    2866=>"111110011",
    2867=>"111011000",
    2868=>"111011000",
    2869=>"000000000",
    2870=>"111010001",
    2871=>"001000100",
    2872=>"011000100",
    2873=>"110011001",
    2874=>"010110000",
    2875=>"011001010",
    2876=>"011001001",
    2877=>"000000000",
    2878=>"110110001",
    2879=>"000100110",
    2880=>"000101001",
    2881=>"010111000",
    2882=>"010010000",
    2883=>"111111010",
    2884=>"000000000",
    2885=>"011000101",
    2886=>"000000000",
    2887=>"100111000",
    2888=>"000000000",
    2889=>"101010110",
    2890=>"000000000",
    2891=>"001101100",
    2892=>"110111011",
    2893=>"111011000",
    2894=>"011111100",
    2895=>"010010000",
    2896=>"111000100",
    2897=>"111000000",
    2898=>"000000111",
    2899=>"111110001",
    2900=>"000000111",
    2901=>"111000000",
    2902=>"000100000",
    2903=>"110000000",
    2904=>"011011111",
    2905=>"111011110",
    2906=>"100000011",
    2907=>"111000111",
    2908=>"000111110",
    2909=>"101111111",
    2910=>"010000000",
    2911=>"000000111",
    2912=>"100111101",
    2913=>"111111110",
    2914=>"111001111",
    2915=>"100000110",
    2916=>"001000100",
    2917=>"000001000",
    2918=>"111111110",
    2919=>"111011100",
    2920=>"000010110",
    2921=>"111101111",
    2922=>"111000000",
    2923=>"000000001",
    2924=>"001111110",
    2925=>"110000111",
    2926=>"000101111",
    2927=>"110111111",
    2928=>"000000111",
    2929=>"100000000",
    2930=>"011011000",
    2931=>"000100111",
    2932=>"000010110",
    2933=>"100101011",
    2934=>"001111111",
    2935=>"111111000",
    2936=>"110101010",
    2937=>"110100000",
    2938=>"110100000",
    2939=>"111111101",
    2940=>"001001111",
    2941=>"011001101",
    2942=>"110110111",
    2943=>"111111000",
    2944=>"001100100",
    2945=>"011111011",
    2946=>"111111010",
    2947=>"111010000",
    2948=>"111101000",
    2949=>"111001101",
    2950=>"110111110",
    2951=>"011111110",
    2952=>"111011100",
    2953=>"000000111",
    2954=>"111110000",
    2955=>"110011001",
    2956=>"010010110",
    2957=>"000100111",
    2958=>"000001100",
    2959=>"111000000",
    2960=>"101111110",
    2961=>"111111000",
    2962=>"001100101",
    2963=>"111010100",
    2964=>"100100000",
    2965=>"000100111",
    2966=>"111000000",
    2967=>"010101011",
    2968=>"000000000",
    2969=>"000001111",
    2970=>"111100100",
    2971=>"010000011",
    2972=>"000010110",
    2973=>"111000000",
    2974=>"010111011",
    2975=>"000100111",
    2976=>"111010000",
    2977=>"111111000",
    2978=>"011001000",
    2979=>"111100100",
    2980=>"110001101",
    2981=>"100111011",
    2982=>"111000000",
    2983=>"001100110",
    2984=>"111111001",
    2985=>"000000111",
    2986=>"111100011",
    2987=>"001000000",
    2988=>"000001001",
    2989=>"100001000",
    2990=>"111111010",
    2991=>"011111101",
    2992=>"110111110",
    2993=>"100110010",
    2994=>"111111001",
    2995=>"010010110",
    2996=>"010011010",
    2997=>"100001011",
    2998=>"110110101",
    2999=>"101000000",
    3000=>"111110101",
    3001=>"000000100",
    3002=>"110001011",
    3003=>"101101001",
    3004=>"111101000",
    3005=>"101100100",
    3006=>"110111111",
    3007=>"011011000",
    3008=>"011111111",
    3009=>"111000000",
    3010=>"000000100",
    3011=>"010011000",
    3012=>"111111010",
    3013=>"001011100",
    3014=>"100000001",
    3015=>"000111010",
    3016=>"011001001",
    3017=>"100000001",
    3018=>"111111000",
    3019=>"001011000",
    3020=>"111010010",
    3021=>"001010000",
    3022=>"100000000",
    3023=>"000101111",
    3024=>"111011101",
    3025=>"011111110",
    3026=>"000001100",
    3027=>"111111111",
    3028=>"110110010",
    3029=>"000000100",
    3030=>"010010000",
    3031=>"000000000",
    3032=>"000000000",
    3033=>"001000111",
    3034=>"100110001",
    3035=>"100011001",
    3036=>"100000100",
    3037=>"000111000",
    3038=>"001000100",
    3039=>"000000000",
    3040=>"000000001",
    3041=>"110011110",
    3042=>"011111111",
    3043=>"000101000",
    3044=>"110111010",
    3045=>"100111100",
    3046=>"110111001",
    3047=>"100001101",
    3048=>"000000101",
    3049=>"000000001",
    3050=>"000110001",
    3051=>"100110000",
    3052=>"110111111",
    3053=>"100000000",
    3054=>"000111000",
    3055=>"000000000",
    3056=>"111111111",
    3057=>"000000111",
    3058=>"011011110",
    3059=>"010100111",
    3060=>"100111111",
    3061=>"001000011",
    3062=>"000100000",
    3063=>"111000000",
    3064=>"010011000",
    3065=>"001010110",
    3066=>"100100000",
    3067=>"100010000",
    3068=>"110010000",
    3069=>"100101011",
    3070=>"001000001",
    3071=>"011010000",
    3072=>"011000000",
    3073=>"000000110",
    3074=>"111101101",
    3075=>"000011111",
    3076=>"111100000",
    3077=>"001011001",
    3078=>"000010011",
    3079=>"100100110",
    3080=>"000110111",
    3081=>"000010111",
    3082=>"011011011",
    3083=>"101100100",
    3084=>"000111111",
    3085=>"000100100",
    3086=>"111101100",
    3087=>"000110101",
    3088=>"110010110",
    3089=>"111111000",
    3090=>"001100100",
    3091=>"000001111",
    3092=>"001000100",
    3093=>"111000000",
    3094=>"111101000",
    3095=>"000100111",
    3096=>"000000000",
    3097=>"111000000",
    3098=>"100100100",
    3099=>"111100000",
    3100=>"111100110",
    3101=>"111011000",
    3102=>"000000000",
    3103=>"111111000",
    3104=>"000000111",
    3105=>"111100100",
    3106=>"000000000",
    3107=>"000100100",
    3108=>"001000011",
    3109=>"000011011",
    3110=>"001011011",
    3111=>"100100111",
    3112=>"111101100",
    3113=>"110010010",
    3114=>"100000001",
    3115=>"110010011",
    3116=>"111001000",
    3117=>"111011011",
    3118=>"000110111",
    3119=>"101101011",
    3120=>"111001000",
    3121=>"000000011",
    3122=>"011011011",
    3123=>"001001001",
    3124=>"000000110",
    3125=>"101001001",
    3126=>"101101101",
    3127=>"000000110",
    3128=>"101011011",
    3129=>"011001111",
    3130=>"111011011",
    3131=>"011001001",
    3132=>"111111000",
    3133=>"001001001",
    3134=>"001011011",
    3135=>"111111011",
    3136=>"000100000",
    3137=>"010101111",
    3138=>"111111111",
    3139=>"111111010",
    3140=>"001001100",
    3141=>"001001110",
    3142=>"111010101",
    3143=>"111011011",
    3144=>"001000010",
    3145=>"110110010",
    3146=>"101000111",
    3147=>"001000100",
    3148=>"111101111",
    3149=>"110100000",
    3150=>"101111111",
    3151=>"110100000",
    3152=>"110010001",
    3153=>"101011001",
    3154=>"111111100",
    3155=>"001111011",
    3156=>"101110100",
    3157=>"000000000",
    3158=>"000000000",
    3159=>"000000000",
    3160=>"101000100",
    3161=>"110111010",
    3162=>"011010010",
    3163=>"111100101",
    3164=>"001100111",
    3165=>"001001001",
    3166=>"011110111",
    3167=>"100010000",
    3168=>"000000100",
    3169=>"001100101",
    3170=>"010000110",
    3171=>"001000100",
    3172=>"001011100",
    3173=>"000001000",
    3174=>"010101111",
    3175=>"101110010",
    3176=>"011010011",
    3177=>"110110110",
    3178=>"101000001",
    3179=>"100000110",
    3180=>"001101100",
    3181=>"000000000",
    3182=>"000000000",
    3183=>"100000000",
    3184=>"101001000",
    3185=>"111001000",
    3186=>"111001101",
    3187=>"000000000",
    3188=>"000100000",
    3189=>"000000001",
    3190=>"000001100",
    3191=>"111111000",
    3192=>"111111111",
    3193=>"101100101",
    3194=>"101011110",
    3195=>"111111111",
    3196=>"000100110",
    3197=>"110010101",
    3198=>"001101011",
    3199=>"111000000",
    3200=>"010110011",
    3201=>"001001000",
    3202=>"000000100",
    3203=>"011010110",
    3204=>"110011001",
    3205=>"110001000",
    3206=>"000000100",
    3207=>"001100111",
    3208=>"111011001",
    3209=>"000100101",
    3210=>"100100110",
    3211=>"110111001",
    3212=>"011100111",
    3213=>"011000000",
    3214=>"110011001",
    3215=>"111011001",
    3216=>"100011001",
    3217=>"110011001",
    3218=>"110010001",
    3219=>"001000110",
    3220=>"110011000",
    3221=>"100010001",
    3222=>"111011010",
    3223=>"110011001",
    3224=>"001100110",
    3225=>"010001100",
    3226=>"001100111",
    3227=>"100110110",
    3228=>"010001000",
    3229=>"000101111",
    3230=>"111011001",
    3231=>"111011001",
    3232=>"001100110",
    3233=>"011001000",
    3234=>"111011000",
    3235=>"100000111",
    3236=>"110111001",
    3237=>"010011000",
    3238=>"000100010",
    3239=>"110010001",
    3240=>"000100000",
    3241=>"110001100",
    3242=>"110111001",
    3243=>"000000001",
    3244=>"000000110",
    3245=>"000100010",
    3246=>"001100110",
    3247=>"100001000",
    3248=>"110011010",
    3249=>"010001100",
    3250=>"111000000",
    3251=>"010011010",
    3252=>"111001000",
    3253=>"001100000",
    3254=>"100011000",
    3255=>"100100111",
    3256=>"101010001",
    3257=>"110011001",
    3258=>"110110011",
    3259=>"000000110",
    3260=>"111111011",
    3261=>"111010000",
    3262=>"111111111",
    3263=>"100011001",
    3264=>"000000001",
    3265=>"000011111",
    3266=>"011000000",
    3267=>"011011110",
    3268=>"111101011",
    3269=>"000000000",
    3270=>"110100111",
    3271=>"000100000",
    3272=>"100100100",
    3273=>"000001111",
    3274=>"111111111",
    3275=>"111100100",
    3276=>"111100100",
    3277=>"010001000",
    3278=>"000000000",
    3279=>"000111110",
    3280=>"000000000",
    3281=>"100111110",
    3282=>"001000000",
    3283=>"000000000",
    3284=>"000100101",
    3285=>"000000001",
    3286=>"111110000",
    3287=>"100010111",
    3288=>"101000000",
    3289=>"001001011",
    3290=>"100000000",
    3291=>"001001011",
    3292=>"100101011",
    3293=>"111110000",
    3294=>"100100111",
    3295=>"110001111",
    3296=>"010100110",
    3297=>"000000111",
    3298=>"000000000",
    3299=>"111000101",
    3300=>"101000001",
    3301=>"111111001",
    3302=>"001011111",
    3303=>"000000001",
    3304=>"011011011",
    3305=>"000000000",
    3306=>"000000101",
    3307=>"110110000",
    3308=>"000000011",
    3309=>"111111111",
    3310=>"111110110",
    3311=>"011011111",
    3312=>"000000001",
    3313=>"000000111",
    3314=>"011111111",
    3315=>"001001001",
    3316=>"010100101",
    3317=>"001001001",
    3318=>"000000101",
    3319=>"100000000",
    3320=>"000001001",
    3321=>"000001111",
    3322=>"000000100",
    3323=>"000001111",
    3324=>"111101001",
    3325=>"111110100",
    3326=>"001111111",
    3327=>"001111111",
    3328=>"001111101",
    3329=>"111110111",
    3330=>"010000000",
    3331=>"110110100",
    3332=>"111101111",
    3333=>"110110101",
    3334=>"110011001",
    3335=>"100010011",
    3336=>"111011001",
    3337=>"011001001",
    3338=>"101100110",
    3339=>"111001001",
    3340=>"100101101",
    3341=>"000001010",
    3342=>"011001001",
    3343=>"001001011",
    3344=>"100100011",
    3345=>"101100100",
    3346=>"101101111",
    3347=>"010000000",
    3348=>"000000000",
    3349=>"001001001",
    3350=>"110110110",
    3351=>"111110100",
    3352=>"100110100",
    3353=>"001001001",
    3354=>"100110111",
    3355=>"001011001",
    3356=>"001001001",
    3357=>"100001111",
    3358=>"011010001",
    3359=>"011001001",
    3360=>"100110110",
    3361=>"101101101",
    3362=>"100100110",
    3363=>"100100100",
    3364=>"100001000",
    3365=>"100000001",
    3366=>"000110101",
    3367=>"110010111",
    3368=>"111010101",
    3369=>"001001001",
    3370=>"101011100",
    3371=>"110100101",
    3372=>"001000100",
    3373=>"000000000",
    3374=>"100110010",
    3375=>"011011011",
    3376=>"001001001",
    3377=>"001001000",
    3378=>"111110100",
    3379=>"111001111",
    3380=>"001010000",
    3381=>"001000110",
    3382=>"000000000",
    3383=>"110110110",
    3384=>"110110100",
    3385=>"110001100",
    3386=>"001000001",
    3387=>"111110100",
    3388=>"100100110",
    3389=>"100100110",
    3390=>"001011010",
    3391=>"011010001",
    3392=>"010110100",
    3393=>"000111111",
    3394=>"110111011",
    3395=>"010111011",
    3396=>"011001001",
    3397=>"110110111",
    3398=>"100001111",
    3399=>"011001000",
    3400=>"010111101",
    3401=>"010000000",
    3402=>"000100000",
    3403=>"101100111",
    3404=>"010011111",
    3405=>"001111110",
    3406=>"110011001",
    3407=>"111111111",
    3408=>"111100101",
    3409=>"000011111",
    3410=>"111110110",
    3411=>"101011000",
    3412=>"111001000",
    3413=>"010111111",
    3414=>"000000000",
    3415=>"000111001",
    3416=>"000101100",
    3417=>"111111100",
    3418=>"011111101",
    3419=>"000001010",
    3420=>"000111111",
    3421=>"111000000",
    3422=>"000111111",
    3423=>"000010110",
    3424=>"110110011",
    3425=>"000110111",
    3426=>"110010100",
    3427=>"111000000",
    3428=>"100000000",
    3429=>"110000000",
    3430=>"000001111",
    3431=>"011111011",
    3432=>"010111111",
    3433=>"111111111",
    3434=>"110110000",
    3435=>"000100101",
    3436=>"111101001",
    3437=>"000111111",
    3438=>"111001111",
    3439=>"111110111",
    3440=>"000000000",
    3441=>"111111000",
    3442=>"101111011",
    3443=>"000110111",
    3444=>"000000010",
    3445=>"001000001",
    3446=>"100011111",
    3447=>"000001011",
    3448=>"101101111",
    3449=>"000000110",
    3450=>"110001001",
    3451=>"111110100",
    3452=>"000111111",
    3453=>"111010000",
    3454=>"001011111",
    3455=>"000111000",
    3456=>"011100111",
    3457=>"111001111",
    3458=>"111111111",
    3459=>"010111000",
    3460=>"100100110",
    3461=>"111001111",
    3462=>"001101101",
    3463=>"000000100",
    3464=>"000100000",
    3465=>"111111101",
    3466=>"001011110",
    3467=>"000001000",
    3468=>"100111100",
    3469=>"111111111",
    3470=>"110001001",
    3471=>"000110111",
    3472=>"101111101",
    3473=>"110111000",
    3474=>"111101111",
    3475=>"100011111",
    3476=>"011001000",
    3477=>"110110110",
    3478=>"000000000",
    3479=>"111000000",
    3480=>"000000000",
    3481=>"111111000",
    3482=>"111100011",
    3483=>"110110000",
    3484=>"000111110",
    3485=>"000000000",
    3486=>"111111111",
    3487=>"110000000",
    3488=>"111000000",
    3489=>"011111100",
    3490=>"111000110",
    3491=>"000000000",
    3492=>"001000010",
    3493=>"100000001",
    3494=>"110011110",
    3495=>"111110111",
    3496=>"111110111",
    3497=>"111111100",
    3498=>"011111100",
    3499=>"011000100",
    3500=>"110101111",
    3501=>"000010100",
    3502=>"011000011",
    3503=>"000111101",
    3504=>"110111000",
    3505=>"111111110",
    3506=>"100011101",
    3507=>"110111110",
    3508=>"000100000",
    3509=>"100000001",
    3510=>"000000000",
    3511=>"101000111",
    3512=>"111111111",
    3513=>"110110000",
    3514=>"111100110",
    3515=>"000000000",
    3516=>"000000000",
    3517=>"000000001",
    3518=>"001101111",
    3519=>"000000000",
    3520=>"100100111",
    3521=>"010111010",
    3522=>"010011011",
    3523=>"010111010",
    3524=>"000011110",
    3525=>"000000100",
    3526=>"000000001",
    3527=>"101000001",
    3528=>"000001000",
    3529=>"111111101",
    3530=>"000010011",
    3531=>"000100110",
    3532=>"011111010",
    3533=>"111111111",
    3534=>"001101001",
    3535=>"000001000",
    3536=>"000000000",
    3537=>"010000000",
    3538=>"000000100",
    3539=>"110100100",
    3540=>"000000111",
    3541=>"010111100",
    3542=>"111101101",
    3543=>"110000000",
    3544=>"000000000",
    3545=>"101100111",
    3546=>"100000001",
    3547=>"000001011",
    3548=>"000000010",
    3549=>"000000100",
    3550=>"110010110",
    3551=>"111111111",
    3552=>"110100000",
    3553=>"000000110",
    3554=>"011001000",
    3555=>"000000100",
    3556=>"011101111",
    3557=>"100000100",
    3558=>"000010111",
    3559=>"111011111",
    3560=>"000001110",
    3561=>"010110000",
    3562=>"010001110",
    3563=>"001101011",
    3564=>"111011110",
    3565=>"000000001",
    3566=>"101000100",
    3567=>"111111111",
    3568=>"100000000",
    3569=>"000000010",
    3570=>"101000100",
    3571=>"000000000",
    3572=>"010010010",
    3573=>"100100000",
    3574=>"101101001",
    3575=>"111011010",
    3576=>"010001010",
    3577=>"000100111",
    3578=>"100000000",
    3579=>"000000111",
    3580=>"001000100",
    3581=>"001000001",
    3582=>"111111111",
    3583=>"010000100",
    3584=>"111111000",
    3585=>"000110111",
    3586=>"111111101",
    3587=>"001011011",
    3588=>"111111001",
    3589=>"000100111",
    3590=>"000000000",
    3591=>"101101001",
    3592=>"111100000",
    3593=>"011111000",
    3594=>"111011011",
    3595=>"111100001",
    3596=>"111110111",
    3597=>"000111111",
    3598=>"111011000",
    3599=>"111101010",
    3600=>"010000111",
    3601=>"010000111",
    3602=>"000000000",
    3603=>"110001111",
    3604=>"001000000",
    3605=>"010110110",
    3606=>"000000111",
    3607=>"000111111",
    3608=>"000010111",
    3609=>"110110110",
    3610=>"000011110",
    3611=>"000011011",
    3612=>"110110000",
    3613=>"111000001",
    3614=>"000000000",
    3615=>"110110100",
    3616=>"101000000",
    3617=>"011011000",
    3618=>"010111111",
    3619=>"000000100",
    3620=>"001000000",
    3621=>"111111000",
    3622=>"100000011",
    3623=>"111011100",
    3624=>"111110000",
    3625=>"011000000",
    3626=>"011111100",
    3627=>"000110110",
    3628=>"001101000",
    3629=>"111011000",
    3630=>"111101000",
    3631=>"101001111",
    3632=>"110110000",
    3633=>"000000000",
    3634=>"011000100",
    3635=>"100000000",
    3636=>"000001111",
    3637=>"011011000",
    3638=>"011001000",
    3639=>"000001111",
    3640=>"000011111",
    3641=>"111100001",
    3642=>"000000000",
    3643=>"101101000",
    3644=>"000000111",
    3645=>"100000010",
    3646=>"101111011",
    3647=>"000000111",
    3648=>"111000010",
    3649=>"111011100",
    3650=>"011111110",
    3651=>"100111111",
    3652=>"110110110",
    3653=>"100010101",
    3654=>"010000100",
    3655=>"001101010",
    3656=>"011001110",
    3657=>"111000000",
    3658=>"111010000",
    3659=>"100111000",
    3660=>"111111111",
    3661=>"110000000",
    3662=>"011110001",
    3663=>"000011010",
    3664=>"000000000",
    3665=>"001111010",
    3666=>"110000100",
    3667=>"000101111",
    3668=>"011000000",
    3669=>"111000000",
    3670=>"011000000",
    3671=>"000011111",
    3672=>"011000000",
    3673=>"110000101",
    3674=>"001100110",
    3675=>"010111010",
    3676=>"111000000",
    3677=>"000101111",
    3678=>"011001001",
    3679=>"111000000",
    3680=>"111001001",
    3681=>"101001001",
    3682=>"110011111",
    3683=>"011100110",
    3684=>"000000111",
    3685=>"111111100",
    3686=>"001101100",
    3687=>"110100001",
    3688=>"000110011",
    3689=>"001000000",
    3690=>"000110110",
    3691=>"011010000",
    3692=>"111101011",
    3693=>"001000111",
    3694=>"101001000",
    3695=>"110000000",
    3696=>"110001010",
    3697=>"000000000",
    3698=>"011100001",
    3699=>"100111111",
    3700=>"101111010",
    3701=>"011000000",
    3702=>"001000110",
    3703=>"010010000",
    3704=>"110010011",
    3705=>"100111011",
    3706=>"111000011",
    3707=>"110000000",
    3708=>"100110001",
    3709=>"010001010",
    3710=>"011111001",
    3711=>"100000000",
    3712=>"000001110",
    3713=>"100000001",
    3714=>"000011111",
    3715=>"111000101",
    3716=>"111110100",
    3717=>"100000000",
    3718=>"001001010",
    3719=>"100000111",
    3720=>"110110100",
    3721=>"001010111",
    3722=>"011100100",
    3723=>"011111110",
    3724=>"101011111",
    3725=>"011110111",
    3726=>"001011111",
    3727=>"111110000",
    3728=>"000000101",
    3729=>"110100000",
    3730=>"011111100",
    3731=>"001111000",
    3732=>"011111000",
    3733=>"110110000",
    3734=>"111101001",
    3735=>"110100001",
    3736=>"000001111",
    3737=>"100001001",
    3738=>"101001111",
    3739=>"001001011",
    3740=>"110110000",
    3741=>"011111110",
    3742=>"100100101",
    3743=>"001000101",
    3744=>"000011110",
    3745=>"110110000",
    3746=>"110100001",
    3747=>"000100000",
    3748=>"110100000",
    3749=>"000011110",
    3750=>"101001101",
    3751=>"011111100",
    3752=>"000011111",
    3753=>"000000000",
    3754=>"111110000",
    3755=>"101000001",
    3756=>"000011111",
    3757=>"000000011",
    3758=>"001011110",
    3759=>"010000111",
    3760=>"110110001",
    3761=>"100100100",
    3762=>"111110100",
    3763=>"110011001",
    3764=>"111000001",
    3765=>"001010111",
    3766=>"011000110",
    3767=>"000100000",
    3768=>"110100001",
    3769=>"000111101",
    3770=>"110100000",
    3771=>"000000011",
    3772=>"111100000",
    3773=>"111111110",
    3774=>"100000000",
    3775=>"100110000",
    3776=>"111101101",
    3777=>"000010000",
    3778=>"110011011",
    3779=>"000000000",
    3780=>"000000110",
    3781=>"100001101",
    3782=>"000000000",
    3783=>"011110110",
    3784=>"001100110",
    3785=>"010010110",
    3786=>"001001111",
    3787=>"111110110",
    3788=>"111111111",
    3789=>"111111010",
    3790=>"011001100",
    3791=>"011010000",
    3792=>"000111111",
    3793=>"111111101",
    3794=>"000000000",
    3795=>"111111111",
    3796=>"001000000",
    3797=>"000000000",
    3798=>"001001001",
    3799=>"101100101",
    3800=>"110111010",
    3801=>"000101000",
    3802=>"001110101",
    3803=>"101110101",
    3804=>"111101000",
    3805=>"111011110",
    3806=>"000000000",
    3807=>"111101000",
    3808=>"110001111",
    3809=>"001000000",
    3810=>"111111111",
    3811=>"000000000",
    3812=>"011101011",
    3813=>"110000110",
    3814=>"100100000",
    3815=>"111111111",
    3816=>"000000000",
    3817=>"110111111",
    3818=>"001100111",
    3819=>"000000001",
    3820=>"011011111",
    3821=>"001001011",
    3822=>"111000010",
    3823=>"110100010",
    3824=>"111101011",
    3825=>"010111000",
    3826=>"111111011",
    3827=>"000001001",
    3828=>"111101000",
    3829=>"000000000",
    3830=>"000000000",
    3831=>"011100011",
    3832=>"000000000",
    3833=>"100001111",
    3834=>"101101010",
    3835=>"000000000",
    3836=>"001101001",
    3837=>"000000000",
    3838=>"111111111",
    3839=>"000010000",
    3840=>"101101001",
    3841=>"000010011",
    3842=>"000100000",
    3843=>"011000110",
    3844=>"111111111",
    3845=>"111111111",
    3846=>"000001011",
    3847=>"111111000",
    3848=>"111001000",
    3849=>"111111000",
    3850=>"111111111",
    3851=>"101110011",
    3852=>"011111000",
    3853=>"001000000",
    3854=>"011101000",
    3855=>"110000000",
    3856=>"001111111",
    3857=>"000000111",
    3858=>"001101110",
    3859=>"000000000",
    3860=>"011000101",
    3861=>"001111001",
    3862=>"001001111",
    3863=>"000000111",
    3864=>"011011010",
    3865=>"111111011",
    3866=>"111111111",
    3867=>"000001111",
    3868=>"000001001",
    3869=>"111000000",
    3870=>"000000111",
    3871=>"001000000",
    3872=>"111111111",
    3873=>"110111111",
    3874=>"011000110",
    3875=>"001011001",
    3876=>"011101101",
    3877=>"111111010",
    3878=>"011111111",
    3879=>"000000000",
    3880=>"111110010",
    3881=>"111111111",
    3882=>"001011000",
    3883=>"001111111",
    3884=>"111101101",
    3885=>"111101111",
    3886=>"111111100",
    3887=>"000000001",
    3888=>"001000100",
    3889=>"010001111",
    3890=>"011111111",
    3891=>"000000000",
    3892=>"010111111",
    3893=>"100100011",
    3894=>"000000000",
    3895=>"110111111",
    3896=>"000110111",
    3897=>"101000000",
    3898=>"011111111",
    3899=>"001000000",
    3900=>"111111111",
    3901=>"100111001",
    3902=>"000000000",
    3903=>"001001001",
    3904=>"100101011",
    3905=>"111111010",
    3906=>"111011111",
    3907=>"110110000",
    3908=>"111011111",
    3909=>"000100100",
    3910=>"111111111",
    3911=>"111001001",
    3912=>"111001111",
    3913=>"101001100",
    3914=>"111110110",
    3915=>"001001001",
    3916=>"111111110",
    3917=>"111010010",
    3918=>"001110100",
    3919=>"000000110",
    3920=>"000000101",
    3921=>"010000111",
    3922=>"011100100",
    3923=>"000000101",
    3924=>"000100111",
    3925=>"010001101",
    3926=>"000000101",
    3927=>"000101111",
    3928=>"000000000",
    3929=>"001001111",
    3930=>"000001001",
    3931=>"001011011",
    3932=>"111000100",
    3933=>"000000101",
    3934=>"111111111",
    3935=>"111000000",
    3936=>"111111101",
    3937=>"100110011",
    3938=>"000000000",
    3939=>"000000001",
    3940=>"000001111",
    3941=>"101110110",
    3942=>"000111100",
    3943=>"000000001",
    3944=>"111111100",
    3945=>"000111011",
    3946=>"011110100",
    3947=>"000000000",
    3948=>"111011100",
    3949=>"000000101",
    3950=>"100101111",
    3951=>"110001101",
    3952=>"110111000",
    3953=>"000000000",
    3954=>"011000000",
    3955=>"000001011",
    3956=>"010111010",
    3957=>"001001100",
    3958=>"111111111",
    3959=>"000000000",
    3960=>"110010000",
    3961=>"000110011",
    3962=>"110001101",
    3963=>"000011011",
    3964=>"110110111",
    3965=>"010000100",
    3966=>"011110000",
    3967=>"111000001",
    3968=>"110101001",
    3969=>"101100101",
    3970=>"101111110",
    3971=>"001011111",
    3972=>"000010111",
    3973=>"001001111",
    3974=>"000100001",
    3975=>"111100000",
    3976=>"001011111",
    3977=>"110000000",
    3978=>"111011101",
    3979=>"000011111",
    3980=>"101001110",
    3981=>"100001100",
    3982=>"001110110",
    3983=>"001011111",
    3984=>"110100001",
    3985=>"101001111",
    3986=>"000111110",
    3987=>"000111110",
    3988=>"000011111",
    3989=>"000000000",
    3990=>"100100111",
    3991=>"110001001",
    3992=>"110100001",
    3993=>"100101111",
    3994=>"111100000",
    3995=>"111000001",
    3996=>"011111001",
    3997=>"100110110",
    3998=>"001001001",
    3999=>"000001011",
    4000=>"011010100",
    4001=>"100001010",
    4002=>"000001001",
    4003=>"100000000",
    4004=>"011001011",
    4005=>"001011110",
    4006=>"111101011",
    4007=>"000111111",
    4008=>"011100000",
    4009=>"000000101",
    4010=>"100011011",
    4011=>"100100000",
    4012=>"000111110",
    4013=>"110100000",
    4014=>"011111000",
    4015=>"000010000",
    4016=>"100101111",
    4017=>"000001111",
    4018=>"000000000",
    4019=>"001101101",
    4020=>"011001001",
    4021=>"010100000",
    4022=>"110100000",
    4023=>"001011110",
    4024=>"101000001",
    4025=>"010010111",
    4026=>"100000000",
    4027=>"111110000",
    4028=>"000001111",
    4029=>"000111001",
    4030=>"111000000",
    4031=>"010110001",
    4032=>"001101001",
    4033=>"010111110",
    4034=>"000111010",
    4035=>"111001001",
    4036=>"111000010",
    4037=>"000000100",
    4038=>"110110010",
    4039=>"101001001",
    4040=>"001011001",
    4041=>"000010001",
    4042=>"111011100",
    4043=>"001010000",
    4044=>"111111111",
    4045=>"111110010",
    4046=>"000001110",
    4047=>"010110111",
    4048=>"000000111",
    4049=>"111111001",
    4050=>"010101111",
    4051=>"000000111",
    4052=>"111011101",
    4053=>"110100110",
    4054=>"111001001",
    4055=>"010101110",
    4056=>"011001001",
    4057=>"010110110",
    4058=>"001001000",
    4059=>"000001110",
    4060=>"111000001",
    4061=>"000100110",
    4062=>"110110100",
    4063=>"011011001",
    4064=>"000000011",
    4065=>"000000101",
    4066=>"010000011",
    4067=>"101000101",
    4068=>"000010111",
    4069=>"001000111",
    4070=>"000001101",
    4071=>"010000111",
    4072=>"101111001",
    4073=>"000000000",
    4074=>"101010011",
    4075=>"101001001",
    4076=>"000000001",
    4077=>"111110011",
    4078=>"101001100",
    4079=>"100000000",
    4080=>"111000001",
    4081=>"000000000",
    4082=>"011000001",
    4083=>"110010110",
    4084=>"111110011",
    4085=>"100000100",
    4086=>"011010011",
    4087=>"000000000",
    4088=>"100100000",
    4089=>"010110000",
    4090=>"110101101",
    4091=>"100100100",
    4092=>"011001000",
    4093=>"001001001",
    4094=>"110110101",
    4095=>"110000000",
    4096=>"100100000",
    4097=>"110111001",
    4098=>"110110111",
    4099=>"111001001",
    4100=>"000000000",
    4101=>"000100110",
    4102=>"100110110",
    4103=>"001101101",
    4104=>"111011101",
    4105=>"000110000",
    4106=>"000100000",
    4107=>"101011001",
    4108=>"110111111",
    4109=>"111111111",
    4110=>"000100110",
    4111=>"100110001",
    4112=>"010110100",
    4113=>"111110010",
    4114=>"000001101",
    4115=>"000000101",
    4116=>"111001101",
    4117=>"000000000",
    4118=>"100100100",
    4119=>"000001010",
    4120=>"111000101",
    4121=>"000110000",
    4122=>"001101011",
    4123=>"110110100",
    4124=>"000001000",
    4125=>"001001111",
    4126=>"100000110",
    4127=>"000010000",
    4128=>"000000010",
    4129=>"001100100",
    4130=>"111010000",
    4131=>"110100000",
    4132=>"000000000",
    4133=>"000110101",
    4134=>"000010110",
    4135=>"110111111",
    4136=>"110111111",
    4137=>"000110111",
    4138=>"000100110",
    4139=>"010000001",
    4140=>"101001101",
    4141=>"001101101",
    4142=>"010000000",
    4143=>"110110100",
    4144=>"111111111",
    4145=>"000010000",
    4146=>"110111001",
    4147=>"111101111",
    4148=>"111011001",
    4149=>"110000001",
    4150=>"000010000",
    4151=>"000110010",
    4152=>"101110001",
    4153=>"110011011",
    4154=>"000101111",
    4155=>"001011011",
    4156=>"100000000",
    4157=>"000010111",
    4158=>"000111101",
    4159=>"110111111",
    4160=>"010010100",
    4161=>"000100011",
    4162=>"110111001",
    4163=>"111111100",
    4164=>"100100110",
    4165=>"100101001",
    4166=>"111111110",
    4167=>"011001110",
    4168=>"111100010",
    4169=>"101101000",
    4170=>"001001111",
    4171=>"000010011",
    4172=>"101001111",
    4173=>"000000000",
    4174=>"000010010",
    4175=>"111000101",
    4176=>"000111111",
    4177=>"101100101",
    4178=>"111111011",
    4179=>"000000000",
    4180=>"100011001",
    4181=>"000000100",
    4182=>"000111111",
    4183=>"000111100",
    4184=>"000100010",
    4185=>"000000111",
    4186=>"001101100",
    4187=>"011010000",
    4188=>"000101111",
    4189=>"111101001",
    4190=>"100111011",
    4191=>"000011010",
    4192=>"010010010",
    4193=>"011011001",
    4194=>"000011000",
    4195=>"001010110",
    4196=>"001111011",
    4197=>"110000011",
    4198=>"110110100",
    4199=>"000000000",
    4200=>"111011010",
    4201=>"000000000",
    4202=>"100010010",
    4203=>"001111111",
    4204=>"010010011",
    4205=>"001010110",
    4206=>"111001101",
    4207=>"000010000",
    4208=>"001000000",
    4209=>"000000111",
    4210=>"101100011",
    4211=>"011000000",
    4212=>"111110000",
    4213=>"111110110",
    4214=>"000010000",
    4215=>"000010011",
    4216=>"000010110",
    4217=>"100010110",
    4218=>"111111110",
    4219=>"001011110",
    4220=>"000101101",
    4221=>"100000001",
    4222=>"000000000",
    4223=>"000010111",
    4224=>"000101111",
    4225=>"111111000",
    4226=>"100111111",
    4227=>"011010111",
    4228=>"000110111",
    4229=>"101111111",
    4230=>"110100001",
    4231=>"000100111",
    4232=>"101100000",
    4233=>"111110000",
    4234=>"011110111",
    4235=>"000000011",
    4236=>"011000111",
    4237=>"101000000",
    4238=>"111001001",
    4239=>"111000000",
    4240=>"100000011",
    4241=>"111000000",
    4242=>"001011100",
    4243=>"111011001",
    4244=>"001000010",
    4245=>"111000000",
    4246=>"000111111",
    4247=>"111110000",
    4248=>"000010111",
    4249=>"111000000",
    4250=>"101011111",
    4251=>"110000001",
    4252=>"111100010",
    4253=>"111000111",
    4254=>"111111000",
    4255=>"111010000",
    4256=>"000001111",
    4257=>"111001000",
    4258=>"100000000",
    4259=>"000000111",
    4260=>"111010010",
    4261=>"000000111",
    4262=>"111001000",
    4263=>"111111101",
    4264=>"000001111",
    4265=>"111110000",
    4266=>"111011000",
    4267=>"111000011",
    4268=>"001101111",
    4269=>"110000111",
    4270=>"000001111",
    4271=>"001101000",
    4272=>"111000000",
    4273=>"111000000",
    4274=>"000000111",
    4275=>"001001000",
    4276=>"111110000",
    4277=>"000000001",
    4278=>"000110110",
    4279=>"000100111",
    4280=>"111011000",
    4281=>"001011111",
    4282=>"100010001",
    4283=>"110011111",
    4284=>"000001111",
    4285=>"000001111",
    4286=>"111111001",
    4287=>"111000010",
    4288=>"000111001",
    4289=>"111010010",
    4290=>"011111001",
    4291=>"100001111",
    4292=>"011011100",
    4293=>"000110110",
    4294=>"111011110",
    4295=>"110101001",
    4296=>"111011000",
    4297=>"101101001",
    4298=>"110100000",
    4299=>"101110100",
    4300=>"111111010",
    4301=>"010010000",
    4302=>"001101100",
    4303=>"001001101",
    4304=>"110010110",
    4305=>"110000010",
    4306=>"011110100",
    4307=>"010000001",
    4308=>"111000000",
    4309=>"010010000",
    4310=>"110000111",
    4311=>"010010011",
    4312=>"010010010",
    4313=>"010010010",
    4314=>"100011011",
    4315=>"110111010",
    4316=>"000010010",
    4317=>"001101111",
    4318=>"011111010",
    4319=>"000000000",
    4320=>"111111000",
    4321=>"001110110",
    4322=>"000000110",
    4323=>"000000111",
    4324=>"000000000",
    4325=>"001100100",
    4326=>"010011011",
    4327=>"000000000",
    4328=>"111111100",
    4329=>"101111000",
    4330=>"001101110",
    4331=>"010000011",
    4332=>"001111100",
    4333=>"111111001",
    4334=>"111101101",
    4335=>"000000000",
    4336=>"111111110",
    4337=>"111011000",
    4338=>"011001000",
    4339=>"111111110",
    4340=>"000000000",
    4341=>"100111001",
    4342=>"000001001",
    4343=>"000111010",
    4344=>"110010011",
    4345=>"111101001",
    4346=>"110111001",
    4347=>"100111000",
    4348=>"111110111",
    4349=>"011001000",
    4350=>"000000000",
    4351=>"000000000",
    4352=>"000001000",
    4353=>"110110011",
    4354=>"100010001",
    4355=>"001110011",
    4356=>"111011000",
    4357=>"100110111",
    4358=>"001010000",
    4359=>"011111001",
    4360=>"011001001",
    4361=>"011010100",
    4362=>"001001011",
    4363=>"000110011",
    4364=>"111011111",
    4365=>"110011000",
    4366=>"010001100",
    4367=>"110100011",
    4368=>"000000000",
    4369=>"111110001",
    4370=>"111001101",
    4371=>"111100000",
    4372=>"011001100",
    4373=>"001100100",
    4374=>"011111100",
    4375=>"101001001",
    4376=>"111000100",
    4377=>"101001110",
    4378=>"111000011",
    4379=>"011001101",
    4380=>"100100001",
    4381=>"100011100",
    4382=>"000000110",
    4383=>"001011100",
    4384=>"011100110",
    4385=>"000100110",
    4386=>"000110110",
    4387=>"111100000",
    4388=>"100011111",
    4389=>"001100110",
    4390=>"111110100",
    4391=>"001000110",
    4392=>"001010100",
    4393=>"101001101",
    4394=>"101001000",
    4395=>"000001100",
    4396=>"101100101",
    4397=>"000110000",
    4398=>"011110110",
    4399=>"101001101",
    4400=>"001011010",
    4401=>"001011011",
    4402=>"111110111",
    4403=>"000100110",
    4404=>"001110001",
    4405=>"110100000",
    4406=>"101100010",
    4407=>"001100101",
    4408=>"110001011",
    4409=>"011001110",
    4410=>"101111011",
    4411=>"000110100",
    4412=>"100100010",
    4413=>"000000001",
    4414=>"110100101",
    4415=>"001100100",
    4416=>"001111011",
    4417=>"101100011",
    4418=>"011111010",
    4419=>"011011001",
    4420=>"111111110",
    4421=>"010011110",
    4422=>"111111011",
    4423=>"100000000",
    4424=>"111111110",
    4425=>"111111110",
    4426=>"000000000",
    4427=>"001101101",
    4428=>"111111110",
    4429=>"110010010",
    4430=>"110101100",
    4431=>"010011111",
    4432=>"111111011",
    4433=>"011111111",
    4434=>"001101111",
    4435=>"110110110",
    4436=>"011011111",
    4437=>"100100100",
    4438=>"000010111",
    4439=>"110100011",
    4440=>"101101101",
    4441=>"100100100",
    4442=>"110011010",
    4443=>"101000100",
    4444=>"010000011",
    4445=>"000010110",
    4446=>"011011111",
    4447=>"001000001",
    4448=>"001001011",
    4449=>"000000000",
    4450=>"000100100",
    4451=>"000000000",
    4452=>"111111110",
    4453=>"000000100",
    4454=>"110111111",
    4455=>"100101111",
    4456=>"000001000",
    4457=>"110111111",
    4458=>"101001101",
    4459=>"000000000",
    4460=>"101101101",
    4461=>"000000001",
    4462=>"000110010",
    4463=>"000001001",
    4464=>"000101101",
    4465=>"000100100",
    4466=>"011010011",
    4467=>"000101011",
    4468=>"000011011",
    4469=>"111111111",
    4470=>"101100100",
    4471=>"100000100",
    4472=>"101001111",
    4473=>"100101101",
    4474=>"100111001",
    4475=>"100000000",
    4476=>"000000010",
    4477=>"000000000",
    4478=>"111100101",
    4479=>"100000000",
    4480=>"000000000",
    4481=>"111000000",
    4482=>"000100000",
    4483=>"000011000",
    4484=>"011011000",
    4485=>"010111000",
    4486=>"110111011",
    4487=>"110111000",
    4488=>"000100100",
    4489=>"111111111",
    4490=>"111111110",
    4491=>"111111001",
    4492=>"010110010",
    4493=>"111111111",
    4494=>"000111110",
    4495=>"111101000",
    4496=>"000010101",
    4497=>"110010110",
    4498=>"010100100",
    4499=>"000111000",
    4500=>"110111111",
    4501=>"010111010",
    4502=>"011011011",
    4503=>"110000111",
    4504=>"000110101",
    4505=>"000000110",
    4506=>"000011001",
    4507=>"010110001",
    4508=>"111101111",
    4509=>"000111000",
    4510=>"101111010",
    4511=>"000101111",
    4512=>"110011000",
    4513=>"100110110",
    4514=>"001000000",
    4515=>"000010000",
    4516=>"111011100",
    4517=>"111111100",
    4518=>"000111010",
    4519=>"000001100",
    4520=>"000010110",
    4521=>"100100000",
    4522=>"101011010",
    4523=>"111100111",
    4524=>"000010000",
    4525=>"000000000",
    4526=>"010010010",
    4527=>"011100000",
    4528=>"000000000",
    4529=>"010011001",
    4530=>"000111000",
    4531=>"000000100",
    4532=>"100111111",
    4533=>"100110100",
    4534=>"110111011",
    4535=>"110110000",
    4536=>"000100000",
    4537=>"011111100",
    4538=>"010010110",
    4539=>"000111000",
    4540=>"000010000",
    4541=>"011001110",
    4542=>"110110010",
    4543=>"111111111",
    4544=>"101001000",
    4545=>"000100110",
    4546=>"111111001",
    4547=>"111010000",
    4548=>"111111000",
    4549=>"001000101",
    4550=>"000000111",
    4551=>"111111000",
    4552=>"111000000",
    4553=>"010000111",
    4554=>"111010000",
    4555=>"001000110",
    4556=>"111000000",
    4557=>"010100010",
    4558=>"010100011",
    4559=>"111101000",
    4560=>"000000111",
    4561=>"000000111",
    4562=>"000101000",
    4563=>"011000001",
    4564=>"011110111",
    4565=>"000000111",
    4566=>"000000111",
    4567=>"000111111",
    4568=>"111110110",
    4569=>"000001111",
    4570=>"100000111",
    4571=>"000000111",
    4572=>"000101111",
    4573=>"111111000",
    4574=>"000000111",
    4575=>"000000111",
    4576=>"111111000",
    4577=>"000110110",
    4578=>"011110101",
    4579=>"111111000",
    4580=>"000101111",
    4581=>"111111000",
    4582=>"000001011",
    4583=>"111011101",
    4584=>"111111001",
    4585=>"000100111",
    4586=>"000011111",
    4587=>"000000100",
    4588=>"100101000",
    4589=>"000000111",
    4590=>"111111000",
    4591=>"000100111",
    4592=>"000010110",
    4593=>"000111111",
    4594=>"001101000",
    4595=>"001001111",
    4596=>"000000111",
    4597=>"111101000",
    4598=>"000100001",
    4599=>"111111000",
    4600=>"000000111",
    4601=>"111011110",
    4602=>"000100000",
    4603=>"111111000",
    4604=>"110000010",
    4605=>"111101000",
    4606=>"110110000",
    4607=>"000011000",
    4608=>"100111011",
    4609=>"110111011",
    4610=>"000000000",
    4611=>"010111011",
    4612=>"000000011",
    4613=>"000000000",
    4614=>"111111111",
    4615=>"111111111",
    4616=>"000000000",
    4617=>"010110101",
    4618=>"111110101",
    4619=>"100000000",
    4620=>"010111000",
    4621=>"101011010",
    4622=>"100000000",
    4623=>"000110000",
    4624=>"111011100",
    4625=>"011110000",
    4626=>"000000000",
    4627=>"101101000",
    4628=>"000000101",
    4629=>"000000000",
    4630=>"001001011",
    4631=>"110100110",
    4632=>"001011011",
    4633=>"011100000",
    4634=>"111111111",
    4635=>"110110110",
    4636=>"100101110",
    4637=>"000000000",
    4638=>"000000000",
    4639=>"100100001",
    4640=>"110100011",
    4641=>"010110000",
    4642=>"100100101",
    4643=>"101011101",
    4644=>"010111001",
    4645=>"000000000",
    4646=>"111111000",
    4647=>"000000000",
    4648=>"111111111",
    4649=>"010010000",
    4650=>"000100010",
    4651=>"001000101",
    4652=>"100000010",
    4653=>"110111011",
    4654=>"100100100",
    4655=>"111111100",
    4656=>"100100100",
    4657=>"110110000",
    4658=>"000000001",
    4659=>"001011100",
    4660=>"000111001",
    4661=>"010101001",
    4662=>"000110110",
    4663=>"100000001",
    4664=>"011110000",
    4665=>"110100000",
    4666=>"100100100",
    4667=>"110110111",
    4668=>"001000010",
    4669=>"000000000",
    4670=>"110111111",
    4671=>"011000001",
    4672=>"100000100",
    4673=>"000000010",
    4674=>"011101111",
    4675=>"000111111",
    4676=>"000110110",
    4677=>"000000100",
    4678=>"111111111",
    4679=>"100000110",
    4680=>"111110110",
    4681=>"010010010",
    4682=>"110011011",
    4683=>"101111101",
    4684=>"110111111",
    4685=>"010000100",
    4686=>"011011101",
    4687=>"000111101",
    4688=>"001110111",
    4689=>"000101101",
    4690=>"000100011",
    4691=>"110101110",
    4692=>"001000000",
    4693=>"011111011",
    4694=>"101101000",
    4695=>"010010100",
    4696=>"001000000",
    4697=>"111110100",
    4698=>"001000100",
    4699=>"111010010",
    4700=>"111110010",
    4701=>"100000000",
    4702=>"011111100",
    4703=>"011011000",
    4704=>"101001111",
    4705=>"010001000",
    4706=>"001001100",
    4707=>"100000100",
    4708=>"000000000",
    4709=>"100100011",
    4710=>"100100000",
    4711=>"000101011",
    4712=>"111110111",
    4713=>"011010010",
    4714=>"011001001",
    4715=>"001000000",
    4716=>"100000001",
    4717=>"011110011",
    4718=>"100000011",
    4719=>"110100100",
    4720=>"001111000",
    4721=>"000000010",
    4722=>"001000101",
    4723=>"111110110",
    4724=>"010011000",
    4725=>"111001001",
    4726=>"111111111",
    4727=>"100000100",
    4728=>"000110100",
    4729=>"110111001",
    4730=>"001101111",
    4731=>"110110100",
    4732=>"101101101",
    4733=>"000000001",
    4734=>"001101101",
    4735=>"100100000",
    4736=>"111010000",
    4737=>"110111111",
    4738=>"110110111",
    4739=>"110111111",
    4740=>"111101110",
    4741=>"101100110",
    4742=>"111111011",
    4743=>"001000101",
    4744=>"110110001",
    4745=>"011000100",
    4746=>"011001111",
    4747=>"000000000",
    4748=>"101101101",
    4749=>"111100010",
    4750=>"111111011",
    4751=>"011001001",
    4752=>"000100110",
    4753=>"000000000",
    4754=>"000110010",
    4755=>"100001110",
    4756=>"111100010",
    4757=>"000000110",
    4758=>"000100101",
    4759=>"111111111",
    4760=>"001100110",
    4761=>"001101101",
    4762=>"010101111",
    4763=>"111000101",
    4764=>"000110111",
    4765=>"110100000",
    4766=>"110010001",
    4767=>"100100001",
    4768=>"000100111",
    4769=>"111000111",
    4770=>"011100110",
    4771=>"001100100",
    4772=>"111111110",
    4773=>"111110010",
    4774=>"101000110",
    4775=>"110111111",
    4776=>"111111110",
    4777=>"111011000",
    4778=>"100100111",
    4779=>"011101101",
    4780=>"111000001",
    4781=>"000000111",
    4782=>"000100111",
    4783=>"110110010",
    4784=>"111111001",
    4785=>"100101001",
    4786=>"000111101",
    4787=>"100010110",
    4788=>"111001000",
    4789=>"110110110",
    4790=>"111001000",
    4791=>"000000100",
    4792=>"000000000",
    4793=>"100100111",
    4794=>"010010100",
    4795=>"111101000",
    4796=>"100101111",
    4797=>"000000011",
    4798=>"110011101",
    4799=>"111101000",
    4800=>"110110111",
    4801=>"011000011",
    4802=>"010000001",
    4803=>"100000000",
    4804=>"001011010",
    4805=>"111111111",
    4806=>"111011001",
    4807=>"111011111",
    4808=>"000011000",
    4809=>"000000000",
    4810=>"000110000",
    4811=>"111111100",
    4812=>"000111010",
    4813=>"110010010",
    4814=>"110111011",
    4815=>"000000000",
    4816=>"111111111",
    4817=>"000000100",
    4818=>"111111111",
    4819=>"111111101",
    4820=>"110110111",
    4821=>"111011010",
    4822=>"111111111",
    4823=>"011011110",
    4824=>"111111111",
    4825=>"001000111",
    4826=>"111111111",
    4827=>"111110100",
    4828=>"111111111",
    4829=>"101101001",
    4830=>"111111110",
    4831=>"111000000",
    4832=>"111111111",
    4833=>"000010011",
    4834=>"111111111",
    4835=>"000000011",
    4836=>"111111111",
    4837=>"111111111",
    4838=>"000011110",
    4839=>"111111011",
    4840=>"111111111",
    4841=>"000000000",
    4842=>"011001011",
    4843=>"111111000",
    4844=>"111111111",
    4845=>"111110101",
    4846=>"110100111",
    4847=>"111011111",
    4848=>"000000110",
    4849=>"010011100",
    4850=>"111111111",
    4851=>"111111101",
    4852=>"000110111",
    4853=>"111111011",
    4854=>"111110110",
    4855=>"100111110",
    4856=>"110110101",
    4857=>"110111100",
    4858=>"111111110",
    4859=>"111110111",
    4860=>"111111111",
    4861=>"000000001",
    4862=>"111110111",
    4863=>"111110010",
    4864=>"111101111",
    4865=>"000010010",
    4866=>"000110010",
    4867=>"010010010",
    4868=>"111111111",
    4869=>"010000100",
    4870=>"011100011",
    4871=>"110111101",
    4872=>"111111111",
    4873=>"100100111",
    4874=>"111111111",
    4875=>"011001100",
    4876=>"111111110",
    4877=>"000000011",
    4878=>"000000011",
    4879=>"101001001",
    4880=>"111100110",
    4881=>"111101000",
    4882=>"011001100",
    4883=>"110001011",
    4884=>"111111111",
    4885=>"000000111",
    4886=>"000000000",
    4887=>"110110010",
    4888=>"101111111",
    4889=>"111001011",
    4890=>"110000001",
    4891=>"100000001",
    4892=>"100000000",
    4893=>"111000101",
    4894=>"001000110",
    4895=>"011001000",
    4896=>"000111101",
    4897=>"000000000",
    4898=>"000000000",
    4899=>"010111101",
    4900=>"111111111",
    4901=>"001000110",
    4902=>"000000000",
    4903=>"000000010",
    4904=>"000010011",
    4905=>"000001111",
    4906=>"011000111",
    4907=>"111010010",
    4908=>"001101111",
    4909=>"111100001",
    4910=>"000000000",
    4911=>"111111111",
    4912=>"111111000",
    4913=>"111111111",
    4914=>"111001000",
    4915=>"010001110",
    4916=>"110110010",
    4917=>"100001100",
    4918=>"000100111",
    4919=>"000111000",
    4920=>"110000000",
    4921=>"000100011",
    4922=>"110110101",
    4923=>"100101010",
    4924=>"101000000",
    4925=>"001110001",
    4926=>"000001000",
    4927=>"000000111",
    4928=>"100100000",
    4929=>"110110110",
    4930=>"011011010",
    4931=>"000110110",
    4932=>"001110110",
    4933=>"000101101",
    4934=>"110110111",
    4935=>"100000000",
    4936=>"011011111",
    4937=>"001011010",
    4938=>"100110110",
    4939=>"011011011",
    4940=>"110111111",
    4941=>"000010000",
    4942=>"100100000",
    4943=>"000000010",
    4944=>"100111111",
    4945=>"000000000",
    4946=>"010100110",
    4947=>"010111110",
    4948=>"111001001",
    4949=>"000000110",
    4950=>"101001001",
    4951=>"000000110",
    4952=>"111001000",
    4953=>"110110000",
    4954=>"001001001",
    4955=>"000011011",
    4956=>"101000000",
    4957=>"001011000",
    4958=>"000111010",
    4959=>"110111111",
    4960=>"111001001",
    4961=>"100111110",
    4962=>"111101101",
    4963=>"110000011",
    4964=>"000000000",
    4965=>"111000111",
    4966=>"110111111",
    4967=>"010110111",
    4968=>"100111111",
    4969=>"010111110",
    4970=>"011111001",
    4971=>"001000101",
    4972=>"001011000",
    4973=>"010110000",
    4974=>"101001001",
    4975=>"110110001",
    4976=>"011111111",
    4977=>"110101101",
    4978=>"011000000",
    4979=>"100010000",
    4980=>"000111110",
    4981=>"011110010",
    4982=>"001011111",
    4983=>"000000000",
    4984=>"010000001",
    4985=>"000000110",
    4986=>"010001111",
    4987=>"001000000",
    4988=>"110000101",
    4989=>"110000000",
    4990=>"100111111",
    4991=>"110111001",
    4992=>"100101011",
    4993=>"010111111",
    4994=>"110011010",
    4995=>"000111111",
    4996=>"111110000",
    4997=>"000001101",
    4998=>"000000001",
    4999=>"110100111",
    5000=>"111000000",
    5001=>"111111000",
    5002=>"111110000",
    5003=>"001111111",
    5004=>"111110000",
    5005=>"010000000",
    5006=>"111011001",
    5007=>"101111111",
    5008=>"000000000",
    5009=>"101001111",
    5010=>"001100111",
    5011=>"100000000",
    5012=>"001000100",
    5013=>"101111011",
    5014=>"111101111",
    5015=>"110010000",
    5016=>"000100000",
    5017=>"111001111",
    5018=>"111001101",
    5019=>"000000110",
    5020=>"111000000",
    5021=>"101000111",
    5022=>"000000000",
    5023=>"111101101",
    5024=>"111011011",
    5025=>"000011111",
    5026=>"000000011",
    5027=>"101100100",
    5028=>"111111111",
    5029=>"101100100",
    5030=>"000011111",
    5031=>"101111100",
    5032=>"010001000",
    5033=>"000000000",
    5034=>"110110110",
    5035=>"111000001",
    5036=>"000001101",
    5037=>"110000001",
    5038=>"111100111",
    5039=>"111000001",
    5040=>"111100000",
    5041=>"111000100",
    5042=>"101000100",
    5043=>"000111111",
    5044=>"000010111",
    5045=>"001001101",
    5046=>"100110111",
    5047=>"000111000",
    5048=>"011011111",
    5049=>"000001011",
    5050=>"111000000",
    5051=>"100000001",
    5052=>"000000011",
    5053=>"101001001",
    5054=>"101010000",
    5055=>"101001111",
    5056=>"110100100",
    5057=>"011101110",
    5058=>"100101001",
    5059=>"111111111",
    5060=>"001101100",
    5061=>"110011011",
    5062=>"101011011",
    5063=>"111001000",
    5064=>"011111111",
    5065=>"110000000",
    5066=>"100101011",
    5067=>"000000000",
    5068=>"111110111",
    5069=>"010011000",
    5070=>"000000000",
    5071=>"010010111",
    5072=>"000110010",
    5073=>"000000111",
    5074=>"110110110",
    5075=>"000100111",
    5076=>"001000100",
    5077=>"101101111",
    5078=>"000000101",
    5079=>"000000000",
    5080=>"000001101",
    5081=>"110100000",
    5082=>"001111110",
    5083=>"101000001",
    5084=>"000000111",
    5085=>"100000000",
    5086=>"111111111",
    5087=>"101000101",
    5088=>"001001110",
    5089=>"001000101",
    5090=>"000011101",
    5091=>"001100100",
    5092=>"000010100",
    5093=>"111010011",
    5094=>"001100001",
    5095=>"001110111",
    5096=>"111111011",
    5097=>"111111010",
    5098=>"100000100",
    5099=>"000000000",
    5100=>"001011100",
    5101=>"000000001",
    5102=>"000000101",
    5103=>"011111101",
    5104=>"111111111",
    5105=>"010001110",
    5106=>"000010100",
    5107=>"111111010",
    5108=>"111111111",
    5109=>"000000101",
    5110=>"111111111",
    5111=>"000000100",
    5112=>"000000000",
    5113=>"101000101",
    5114=>"111011011",
    5115=>"000000000",
    5116=>"000101111",
    5117=>"000000001",
    5118=>"110111111",
    5119=>"100000101",
    5120=>"001000000",
    5121=>"111111111",
    5122=>"000000000",
    5123=>"010111010",
    5124=>"110000001",
    5125=>"111101111",
    5126=>"011111111",
    5127=>"000000000",
    5128=>"111111111",
    5129=>"000111110",
    5130=>"101111111",
    5131=>"100000111",
    5132=>"010111110",
    5133=>"000111101",
    5134=>"001000001",
    5135=>"001001000",
    5136=>"110110111",
    5137=>"111001101",
    5138=>"000000001",
    5139=>"110101111",
    5140=>"100111000",
    5141=>"000101001",
    5142=>"011000000",
    5143=>"110111111",
    5144=>"101000100",
    5145=>"001000101",
    5146=>"001101111",
    5147=>"000101101",
    5148=>"111000111",
    5149=>"111000111",
    5150=>"110111111",
    5151=>"101000000",
    5152=>"111111111",
    5153=>"110111111",
    5154=>"111111111",
    5155=>"101000100",
    5156=>"111101101",
    5157=>"001000000",
    5158=>"111111110",
    5159=>"000000000",
    5160=>"000000000",
    5161=>"000000000",
    5162=>"100111111",
    5163=>"010110111",
    5164=>"000001001",
    5165=>"001001110",
    5166=>"111111111",
    5167=>"100110101",
    5168=>"110100100",
    5169=>"000111101",
    5170=>"001001111",
    5171=>"000000011",
    5172=>"011111110",
    5173=>"001000000",
    5174=>"000000000",
    5175=>"101100000",
    5176=>"111111111",
    5177=>"000000000",
    5178=>"100001001",
    5179=>"001000000",
    5180=>"001000000",
    5181=>"101000101",
    5182=>"000000000",
    5183=>"110111000",
    5184=>"111111111",
    5185=>"000000000",
    5186=>"000000110",
    5187=>"011011011",
    5188=>"111011011",
    5189=>"000000001",
    5190=>"000000000",
    5191=>"011111111",
    5192=>"000000000",
    5193=>"111010110",
    5194=>"111111110",
    5195=>"000000000",
    5196=>"000110110",
    5197=>"000000010",
    5198=>"101000001",
    5199=>"011111010",
    5200=>"000000000",
    5201=>"111111111",
    5202=>"000000000",
    5203=>"110000001",
    5204=>"000000000",
    5205=>"000000000",
    5206=>"000100111",
    5207=>"111000011",
    5208=>"000000111",
    5209=>"111110100",
    5210=>"000000110",
    5211=>"111111111",
    5212=>"111100100",
    5213=>"011010110",
    5214=>"000000000",
    5215=>"100100110",
    5216=>"100000001",
    5217=>"100000000",
    5218=>"000000000",
    5219=>"111111110",
    5220=>"000001000",
    5221=>"111100100",
    5222=>"111111111",
    5223=>"000000000",
    5224=>"011111111",
    5225=>"011111011",
    5226=>"000000100",
    5227=>"110100100",
    5228=>"111111011",
    5229=>"111111111",
    5230=>"001011111",
    5231=>"000000000",
    5232=>"011000000",
    5233=>"101000001",
    5234=>"111111011",
    5235=>"111111110",
    5236=>"110111110",
    5237=>"111111111",
    5238=>"111111111",
    5239=>"110100001",
    5240=>"100100001",
    5241=>"110100101",
    5242=>"110101101",
    5243=>"111111011",
    5244=>"110111111",
    5245=>"000000000",
    5246=>"111111111",
    5247=>"101101001",
    5248=>"111001100",
    5249=>"001111000",
    5250=>"000000101",
    5251=>"000000101",
    5252=>"100110110",
    5253=>"100011001",
    5254=>"110111100",
    5255=>"011100100",
    5256=>"111101011",
    5257=>"010000000",
    5258=>"001101101",
    5259=>"110111011",
    5260=>"000111010",
    5261=>"001001001",
    5262=>"100110011",
    5263=>"011001100",
    5264=>"000000001",
    5265=>"001000101",
    5266=>"100110011",
    5267=>"001001001",
    5268=>"110110010",
    5269=>"000000000",
    5270=>"000110111",
    5271=>"001111111",
    5272=>"000000110",
    5273=>"000000000",
    5274=>"001001111",
    5275=>"100111100",
    5276=>"010110111",
    5277=>"000000001",
    5278=>"111111111",
    5279=>"111111111",
    5280=>"100100101",
    5281=>"111111110",
    5282=>"000111000",
    5283=>"000100101",
    5284=>"000100000",
    5285=>"111011011",
    5286=>"111111100",
    5287=>"100001101",
    5288=>"111111000",
    5289=>"111101000",
    5290=>"000110010",
    5291=>"000110111",
    5292=>"111111011",
    5293=>"111111100",
    5294=>"000110010",
    5295=>"100101010",
    5296=>"110111110",
    5297=>"011001011",
    5298=>"000000011",
    5299=>"110111110",
    5300=>"110110110",
    5301=>"110111001",
    5302=>"101100111",
    5303=>"001001111",
    5304=>"000111011",
    5305=>"000010110",
    5306=>"011111100",
    5307=>"011100100",
    5308=>"011001111",
    5309=>"001000101",
    5310=>"001000011",
    5311=>"001000110",
    5312=>"101000011",
    5313=>"010110011",
    5314=>"011100011",
    5315=>"110110000",
    5316=>"001101011",
    5317=>"001100101",
    5318=>"000111000",
    5319=>"101011111",
    5320=>"011001100",
    5321=>"000001111",
    5322=>"001010110",
    5323=>"010101111",
    5324=>"111111111",
    5325=>"110110000",
    5326=>"011101000",
    5327=>"111000010",
    5328=>"000110110",
    5329=>"011011111",
    5330=>"000001110",
    5331=>"000000110",
    5332=>"110100100",
    5333=>"101000000",
    5334=>"001101111",
    5335=>"000000110",
    5336=>"001011111",
    5337=>"011101011",
    5338=>"001011111",
    5339=>"011011011",
    5340=>"000001011",
    5341=>"001001110",
    5342=>"100000100",
    5343=>"110110000",
    5344=>"000010011",
    5345=>"011100110",
    5346=>"000000010",
    5347=>"001001101",
    5348=>"111100000",
    5349=>"011111100",
    5350=>"100101111",
    5351=>"011110110",
    5352=>"111011001",
    5353=>"110001000",
    5354=>"010001110",
    5355=>"111110000",
    5356=>"001001001",
    5357=>"001000010",
    5358=>"001001110",
    5359=>"110111010",
    5360=>"001001011",
    5361=>"001001111",
    5362=>"011001111",
    5363=>"000000101",
    5364=>"100110110",
    5365=>"001001010",
    5366=>"110010000",
    5367=>"000000000",
    5368=>"100000111",
    5369=>"001101011",
    5370=>"000001001",
    5371=>"001011001",
    5372=>"001001111",
    5373=>"001011111",
    5374=>"101110001",
    5375=>"110110000",
    5376=>"110110101",
    5377=>"000011100",
    5378=>"000000000",
    5379=>"110110100",
    5380=>"000000000",
    5381=>"111000000",
    5382=>"110111111",
    5383=>"000000000",
    5384=>"100000100",
    5385=>"100001001",
    5386=>"111111111",
    5387=>"000000100",
    5388=>"111111011",
    5389=>"011001000",
    5390=>"001101000",
    5391=>"111010011",
    5392=>"111110110",
    5393=>"000000001",
    5394=>"011100100",
    5395=>"001000011",
    5396=>"000100100",
    5397=>"011001001",
    5398=>"110000001",
    5399=>"000100011",
    5400=>"000001001",
    5401=>"001001101",
    5402=>"000010000",
    5403=>"111000001",
    5404=>"001100011",
    5405=>"011011010",
    5406=>"111111110",
    5407=>"100100100",
    5408=>"100110100",
    5409=>"111111111",
    5410=>"011101011",
    5411=>"011001001",
    5412=>"111111111",
    5413=>"000110000",
    5414=>"000000000",
    5415=>"011011111",
    5416=>"111111110",
    5417=>"000100000",
    5418=>"011001100",
    5419=>"111000111",
    5420=>"101101101",
    5421=>"111101101",
    5422=>"100110010",
    5423=>"111111101",
    5424=>"110110110",
    5425=>"000000001",
    5426=>"011000001",
    5427=>"111111110",
    5428=>"010110010",
    5429=>"000000000",
    5430=>"001101000",
    5431=>"101100000",
    5432=>"010110111",
    5433=>"100100000",
    5434=>"110111111",
    5435=>"110111111",
    5436=>"110010011",
    5437=>"000010000",
    5438=>"001001001",
    5439=>"001001000",
    5440=>"000000000",
    5441=>"000000000",
    5442=>"100010001",
    5443=>"001001111",
    5444=>"000000000",
    5445=>"111000111",
    5446=>"111111111",
    5447=>"100001011",
    5448=>"111001010",
    5449=>"000000000",
    5450=>"000000000",
    5451=>"101000000",
    5452=>"101101111",
    5453=>"101111111",
    5454=>"000101100",
    5455=>"100110110",
    5456=>"011110110",
    5457=>"111001000",
    5458=>"000100100",
    5459=>"100100111",
    5460=>"100000000",
    5461=>"111111111",
    5462=>"001000000",
    5463=>"111011101",
    5464=>"111011011",
    5465=>"000000000",
    5466=>"110000011",
    5467=>"101111000",
    5468=>"000101000",
    5469=>"111000100",
    5470=>"111111111",
    5471=>"000100111",
    5472=>"000111111",
    5473=>"000000000",
    5474=>"001000000",
    5475=>"000000000",
    5476=>"111001101",
    5477=>"001100100",
    5478=>"000000000",
    5479=>"100010010",
    5480=>"000001000",
    5481=>"000100000",
    5482=>"011101110",
    5483=>"000000000",
    5484=>"000000000",
    5485=>"111000111",
    5486=>"000000000",
    5487=>"111111110",
    5488=>"111100100",
    5489=>"000000000",
    5490=>"111011000",
    5491=>"111011111",
    5492=>"100111101",
    5493=>"000000000",
    5494=>"000000000",
    5495=>"100111111",
    5496=>"001100001",
    5497=>"111001001",
    5498=>"101010000",
    5499=>"100001000",
    5500=>"000011010",
    5501=>"000010010",
    5502=>"110111111",
    5503=>"000000000",
    5504=>"111011101",
    5505=>"011110111",
    5506=>"010000111",
    5507=>"101101101",
    5508=>"011111101",
    5509=>"110110100",
    5510=>"111011011",
    5511=>"011001001",
    5512=>"111100101",
    5513=>"001001111",
    5514=>"001011111",
    5515=>"111100100",
    5516=>"110000111",
    5517=>"011010011",
    5518=>"101100100",
    5519=>"011001001",
    5520=>"010110110",
    5521=>"110100000",
    5522=>"000001001",
    5523=>"011011011",
    5524=>"000110100",
    5525=>"000000000",
    5526=>"100111111",
    5527=>"000111111",
    5528=>"100110110",
    5529=>"110110010",
    5530=>"011011011",
    5531=>"001011010",
    5532=>"110010110",
    5533=>"000100111",
    5534=>"100100100",
    5535=>"101000010",
    5536=>"011001001",
    5537=>"110101100",
    5538=>"100110110",
    5539=>"001010001",
    5540=>"100100100",
    5541=>"100100111",
    5542=>"011011011",
    5543=>"111001001",
    5544=>"000000110",
    5545=>"100100000",
    5546=>"101100011",
    5547=>"100000010",
    5548=>"101100000",
    5549=>"100001001",
    5550=>"001001101",
    5551=>"000000011",
    5552=>"010010110",
    5553=>"010010111",
    5554=>"100100000",
    5555=>"111100100",
    5556=>"110011111",
    5557=>"001001000",
    5558=>"111001000",
    5559=>"110000000",
    5560=>"000011011",
    5561=>"101101001",
    5562=>"101101100",
    5563=>"101001001",
    5564=>"110111000",
    5565=>"110100100",
    5566=>"111000100",
    5567=>"001101111",
    5568=>"100111011",
    5569=>"111111011",
    5570=>"111101110",
    5571=>"011001111",
    5572=>"001110110",
    5573=>"000110110",
    5574=>"010101101",
    5575=>"110100101",
    5576=>"011000110",
    5577=>"101001000",
    5578=>"100011011",
    5579=>"001110100",
    5580=>"000101111",
    5581=>"011011000",
    5582=>"001111100",
    5583=>"100000100",
    5584=>"010000111",
    5585=>"010000110",
    5586=>"001100100",
    5587=>"110010001",
    5588=>"000000000",
    5589=>"010010000",
    5590=>"011010111",
    5591=>"011000001",
    5592=>"000000000",
    5593=>"010000000",
    5594=>"100000001",
    5595=>"100000101",
    5596=>"111111000",
    5597=>"101100111",
    5598=>"010111111",
    5599=>"000011000",
    5600=>"000000101",
    5601=>"111001001",
    5602=>"001010010",
    5603=>"000000101",
    5604=>"000000000",
    5605=>"000110110",
    5606=>"111111110",
    5607=>"011111101",
    5608=>"101000011",
    5609=>"000000010",
    5610=>"011000010",
    5611=>"000011011",
    5612=>"110111100",
    5613=>"100011001",
    5614=>"100100100",
    5615=>"110110000",
    5616=>"000010001",
    5617=>"011000000",
    5618=>"011001000",
    5619=>"110110010",
    5620=>"110101000",
    5621=>"100001001",
    5622=>"001011100",
    5623=>"000001000",
    5624=>"110010011",
    5625=>"110111001",
    5626=>"110011111",
    5627=>"110110001",
    5628=>"000010111",
    5629=>"000000100",
    5630=>"110111111",
    5631=>"010111000",
    5632=>"001101000",
    5633=>"011100010",
    5634=>"001000110",
    5635=>"101101100",
    5636=>"100110110",
    5637=>"001000001",
    5638=>"000100110",
    5639=>"111001101",
    5640=>"000000010",
    5641=>"011001011",
    5642=>"000100110",
    5643=>"000100100",
    5644=>"111111000",
    5645=>"011101110",
    5646=>"100110011",
    5647=>"011011010",
    5648=>"000100011",
    5649=>"011001001",
    5650=>"100110000",
    5651=>"000110111",
    5652=>"000001000",
    5653=>"100100110",
    5654=>"011011011",
    5655=>"100110011",
    5656=>"001001001",
    5657=>"011001011",
    5658=>"001001101",
    5659=>"100010110",
    5660=>"100111001",
    5661=>"011011001",
    5662=>"011001110",
    5663=>"001001011",
    5664=>"100100100",
    5665=>"000100100",
    5666=>"110110011",
    5667=>"001001100",
    5668=>"110011001",
    5669=>"101000010",
    5670=>"000001000",
    5671=>"000100110",
    5672=>"000110100",
    5673=>"000000011",
    5674=>"111110011",
    5675=>"011000001",
    5676=>"101010011",
    5677=>"100110110",
    5678=>"110111100",
    5679=>"000000110",
    5680=>"110011011",
    5681=>"100100000",
    5682=>"000100010",
    5683=>"100001000",
    5684=>"110001001",
    5685=>"000000100",
    5686=>"110110011",
    5687=>"100100110",
    5688=>"001100110",
    5689=>"100001100",
    5690=>"100110010",
    5691=>"101001011",
    5692=>"111010011",
    5693=>"010001011",
    5694=>"110101101",
    5695=>"000100100",
    5696=>"000001100",
    5697=>"111011110",
    5698=>"011000001",
    5699=>"011001011",
    5700=>"001011011",
    5701=>"001001001",
    5702=>"110110110",
    5703=>"000110110",
    5704=>"001001001",
    5705=>"011001001",
    5706=>"100100110",
    5707=>"001001001",
    5708=>"111000011",
    5709=>"111010010",
    5710=>"000001001",
    5711=>"100100101",
    5712=>"011011011",
    5713=>"000110011",
    5714=>"000000001",
    5715=>"110110110",
    5716=>"100001000",
    5717=>"000000111",
    5718=>"111111111",
    5719=>"110110100",
    5720=>"111010010",
    5721=>"111110110",
    5722=>"110110110",
    5723=>"110110101",
    5724=>"001111000",
    5725=>"111001001",
    5726=>"001011011",
    5727=>"000001010",
    5728=>"001100100",
    5729=>"001011111",
    5730=>"011011001",
    5731=>"101110110",
    5732=>"000001000",
    5733=>"100001001",
    5734=>"111110110",
    5735=>"000000000",
    5736=>"000000101",
    5737=>"100100101",
    5738=>"011011001",
    5739=>"010010010",
    5740=>"011110100",
    5741=>"100100110",
    5742=>"101100000",
    5743=>"001000110",
    5744=>"100100110",
    5745=>"000110110",
    5746=>"001011011",
    5747=>"010010000",
    5748=>"001010111",
    5749=>"000000101",
    5750=>"000000001",
    5751=>"100010011",
    5752=>"100110101",
    5753=>"100100101",
    5754=>"000000010",
    5755=>"100100100",
    5756=>"000100111",
    5757=>"000001011",
    5758=>"000101100",
    5759=>"000010001",
    5760=>"011010010",
    5761=>"111011011",
    5762=>"100100100",
    5763=>"101101001",
    5764=>"110100100",
    5765=>"001001101",
    5766=>"110100111",
    5767=>"010110100",
    5768=>"101100011",
    5769=>"111111000",
    5770=>"100100100",
    5771=>"010010110",
    5772=>"101000101",
    5773=>"110100111",
    5774=>"110010110",
    5775=>"100100100",
    5776=>"000000100",
    5777=>"001001001",
    5778=>"001001000",
    5779=>"000100001",
    5780=>"011011011",
    5781=>"011010010",
    5782=>"011011011",
    5783=>"001011010",
    5784=>"001011000",
    5785=>"010010010",
    5786=>"100110010",
    5787=>"110110110",
    5788=>"100100110",
    5789=>"001001011",
    5790=>"011000110",
    5791=>"011110000",
    5792=>"100100100",
    5793=>"000011110",
    5794=>"011010011",
    5795=>"000000111",
    5796=>"001001001",
    5797=>"001100000",
    5798=>"111001011",
    5799=>"100000111",
    5800=>"010010100",
    5801=>"011000000",
    5802=>"101010010",
    5803=>"011011011",
    5804=>"011010010",
    5805=>"111100000",
    5806=>"100100100",
    5807=>"010000100",
    5808=>"111011011",
    5809=>"000011110",
    5810=>"101110110",
    5811=>"110101110",
    5812=>"110110100",
    5813=>"010110111",
    5814=>"111110110",
    5815=>"011011111",
    5816=>"011001011",
    5817=>"010110000",
    5818=>"011010110",
    5819=>"010110100",
    5820=>"100100101",
    5821=>"001001001",
    5822=>"111110100",
    5823=>"110000100",
    5824=>"111001000",
    5825=>"011110110",
    5826=>"111110110",
    5827=>"001111111",
    5828=>"101111001",
    5829=>"000110111",
    5830=>"111111110",
    5831=>"011101001",
    5832=>"100011101",
    5833=>"011000110",
    5834=>"101011000",
    5835=>"011101110",
    5836=>"111111111",
    5837=>"011000000",
    5838=>"000010000",
    5839=>"110011000",
    5840=>"111110110",
    5841=>"001000111",
    5842=>"110010100",
    5843=>"111000000",
    5844=>"011000100",
    5845=>"101111001",
    5846=>"000000000",
    5847=>"111011111",
    5848=>"010000101",
    5849=>"000100000",
    5850=>"110010111",
    5851=>"110100111",
    5852=>"000000000",
    5853=>"011111010",
    5854=>"110111111",
    5855=>"000000110",
    5856=>"110111000",
    5857=>"011001000",
    5858=>"010011000",
    5859=>"100000100",
    5860=>"111111101",
    5861=>"001111110",
    5862=>"110000001",
    5863=>"001100110",
    5864=>"110111111",
    5865=>"011111000",
    5866=>"001001011",
    5867=>"100000000",
    5868=>"110110000",
    5869=>"111111111",
    5870=>"111000111",
    5871=>"110010000",
    5872=>"000101111",
    5873=>"000000000",
    5874=>"101000111",
    5875=>"101010001",
    5876=>"011010000",
    5877=>"100101100",
    5878=>"001001100",
    5879=>"000011000",
    5880=>"000000000",
    5881=>"111100001",
    5882=>"011011010",
    5883=>"000000000",
    5884=>"000001011",
    5885=>"010000001",
    5886=>"100011001",
    5887=>"010010000",
    5888=>"101000111",
    5889=>"101101001",
    5890=>"000001011",
    5891=>"111111111",
    5892=>"101101001",
    5893=>"011000100",
    5894=>"111001010",
    5895=>"001000001",
    5896=>"001000011",
    5897=>"011000000",
    5898=>"001001111",
    5899=>"000000000",
    5900=>"101100101",
    5901=>"000101111",
    5902=>"111111111",
    5903=>"110100100",
    5904=>"000101110",
    5905=>"111100100",
    5906=>"100111111",
    5907=>"011011011",
    5908=>"000000001",
    5909=>"000000000",
    5910=>"100100100",
    5911=>"000000000",
    5912=>"100100111",
    5913=>"100100100",
    5914=>"000000111",
    5915=>"000000000",
    5916=>"110110100",
    5917=>"101101110",
    5918=>"001001010",
    5919=>"000001011",
    5920=>"100110001",
    5921=>"001001000",
    5922=>"000100111",
    5923=>"111111100",
    5924=>"000110000",
    5925=>"000110000",
    5926=>"101100101",
    5927=>"010111111",
    5928=>"111110111",
    5929=>"011011111",
    5930=>"100000100",
    5931=>"100000000",
    5932=>"011011111",
    5933=>"110110110",
    5934=>"100100100",
    5935=>"100111110",
    5936=>"111111111",
    5937=>"000100000",
    5938=>"110100100",
    5939=>"000010000",
    5940=>"001001011",
    5941=>"000001101",
    5942=>"010101011",
    5943=>"000100001",
    5944=>"011011111",
    5945=>"111111111",
    5946=>"011101011",
    5947=>"000000000",
    5948=>"000001111",
    5949=>"110100000",
    5950=>"001000010",
    5951=>"101111110",
    5952=>"001000100",
    5953=>"100100000",
    5954=>"111111011",
    5955=>"111011000",
    5956=>"111011111",
    5957=>"110001000",
    5958=>"001100100",
    5959=>"000000000",
    5960=>"111001001",
    5961=>"111100110",
    5962=>"000000110",
    5963=>"101111011",
    5964=>"111011101",
    5965=>"111100101",
    5966=>"111011101",
    5967=>"000000101",
    5968=>"111100110",
    5969=>"110011000",
    5970=>"101111001",
    5971=>"000000100",
    5972=>"001111100",
    5973=>"001000101",
    5974=>"111011001",
    5975=>"100100100",
    5976=>"101101111",
    5977=>"001001000",
    5978=>"100000000",
    5979=>"001000100",
    5980=>"110111101",
    5981=>"110011001",
    5982=>"111111110",
    5983=>"011001100",
    5984=>"001100110",
    5985=>"111011011",
    5986=>"111110110",
    5987=>"000110011",
    5988=>"110011100",
    5989=>"000001001",
    5990=>"000100100",
    5991=>"001001111",
    5992=>"001100011",
    5993=>"000000100",
    5994=>"111011101",
    5995=>"111100100",
    5996=>"001100111",
    5997=>"001100100",
    5998=>"010011011",
    5999=>"001101111",
    6000=>"111011101",
    6001=>"100100100",
    6002=>"100110011",
    6003=>"011101101",
    6004=>"111100100",
    6005=>"001000100",
    6006=>"001100111",
    6007=>"000000100",
    6008=>"000100100",
    6009=>"100100001",
    6010=>"000000000",
    6011=>"001000100",
    6012=>"000000000",
    6013=>"000000000",
    6014=>"000000000",
    6015=>"001101111",
    6016=>"101100100",
    6017=>"011011110",
    6018=>"100100100",
    6019=>"011011111",
    6020=>"000001101",
    6021=>"011001011",
    6022=>"110110100",
    6023=>"100100100",
    6024=>"011011001",
    6025=>"100100100",
    6026=>"000100111",
    6027=>"100110100",
    6028=>"001100001",
    6029=>"101100101",
    6030=>"100100100",
    6031=>"011011011",
    6032=>"110000100",
    6033=>"011011011",
    6034=>"000010000",
    6035=>"111001110",
    6036=>"110111100",
    6037=>"100000100",
    6038=>"111111111",
    6039=>"010011011",
    6040=>"100100100",
    6041=>"000000000",
    6042=>"010011010",
    6043=>"100010100",
    6044=>"001101101",
    6045=>"111110000",
    6046=>"111011110",
    6047=>"100100100",
    6048=>"001000001",
    6049=>"000001111",
    6050=>"011011000",
    6051=>"001001001",
    6052=>"010010010",
    6053=>"100100100",
    6054=>"010011010",
    6055=>"000011001",
    6056=>"100100100",
    6057=>"001001000",
    6058=>"010110110",
    6059=>"011010010",
    6060=>"100100100",
    6061=>"001100100",
    6062=>"101100100",
    6063=>"100111100",
    6064=>"010110110",
    6065=>"011010010",
    6066=>"010010100",
    6067=>"111111111",
    6068=>"000100100",
    6069=>"100100100",
    6070=>"100000100",
    6071=>"011011010",
    6072=>"011011010",
    6073=>"101101110",
    6074=>"000001001",
    6075=>"100111100",
    6076=>"010011011",
    6077=>"011011011",
    6078=>"000001000",
    6079=>"000000100",
    6080=>"011011100",
    6081=>"111001101",
    6082=>"110100001",
    6083=>"111111000",
    6084=>"111111011",
    6085=>"010000111",
    6086=>"111111111",
    6087=>"111010000",
    6088=>"000000101",
    6089=>"100101111",
    6090=>"111111010",
    6091=>"100101001",
    6092=>"111101101",
    6093=>"111100111",
    6094=>"001000000",
    6095=>"100001010",
    6096=>"111000000",
    6097=>"101000111",
    6098=>"111111101",
    6099=>"000000000",
    6100=>"111111101",
    6101=>"111010000",
    6102=>"111100101",
    6103=>"110010000",
    6104=>"011010000",
    6105=>"101011010",
    6106=>"100000011",
    6107=>"001001001",
    6108=>"000000000",
    6109=>"001000111",
    6110=>"011111111",
    6111=>"111101011",
    6112=>"111110000",
    6113=>"110011111",
    6114=>"000000000",
    6115=>"000000000",
    6116=>"010110101",
    6117=>"111100000",
    6118=>"000110111",
    6119=>"000000000",
    6120=>"011111011",
    6121=>"000000010",
    6122=>"100111110",
    6123=>"111110110",
    6124=>"001001000",
    6125=>"001011010",
    6126=>"111111000",
    6127=>"011111000",
    6128=>"110100001",
    6129=>"000000000",
    6130=>"111001101",
    6131=>"000000001",
    6132=>"000111111",
    6133=>"111100010",
    6134=>"010010001",
    6135=>"011011011",
    6136=>"000100100",
    6137=>"000111111",
    6138=>"011111011",
    6139=>"001011011",
    6140=>"010010100",
    6141=>"001010000",
    6142=>"000000000",
    6143=>"011010000",
    6144=>"000001101",
    6145=>"011111011",
    6146=>"110111110",
    6147=>"100110110",
    6148=>"100100110",
    6149=>"011111111",
    6150=>"110100100",
    6151=>"111101000",
    6152=>"110110110",
    6153=>"110100100",
    6154=>"100110100",
    6155=>"000100100",
    6156=>"001001101",
    6157=>"011100011",
    6158=>"110000100",
    6159=>"110110100",
    6160=>"101101010",
    6161=>"011011011",
    6162=>"000000100",
    6163=>"110000100",
    6164=>"000000100",
    6165=>"010001000",
    6166=>"001011011",
    6167=>"111101111",
    6168=>"001001001",
    6169=>"001011011",
    6170=>"011011000",
    6171=>"100101001",
    6172=>"011111011",
    6173=>"001101101",
    6174=>"011110111",
    6175=>"110100110",
    6176=>"110100100",
    6177=>"110110100",
    6178=>"000010001",
    6179=>"111000001",
    6180=>"110010100",
    6181=>"100110111",
    6182=>"100100100",
    6183=>"011000000",
    6184=>"010011011",
    6185=>"000110000",
    6186=>"011100101",
    6187=>"001001001",
    6188=>"001101101",
    6189=>"100000011",
    6190=>"110100110",
    6191=>"111100100",
    6192=>"100101001",
    6193=>"110000110",
    6194=>"000011011",
    6195=>"000111001",
    6196=>"101100100",
    6197=>"000000101",
    6198=>"100001101",
    6199=>"011010001",
    6200=>"111011011",
    6201=>"100101100",
    6202=>"100110111",
    6203=>"100100100",
    6204=>"011011011",
    6205=>"001001011",
    6206=>"011110110",
    6207=>"110100001",
    6208=>"100100100",
    6209=>"001011101",
    6210=>"111111111",
    6211=>"011111000",
    6212=>"111111111",
    6213=>"001001100",
    6214=>"001000001",
    6215=>"110111111",
    6216=>"111111111",
    6217=>"001011011",
    6218=>"011000001",
    6219=>"111111111",
    6220=>"011111011",
    6221=>"000111110",
    6222=>"110110110",
    6223=>"000111010",
    6224=>"111111010",
    6225=>"111110100",
    6226=>"101111110",
    6227=>"100000000",
    6228=>"000111111",
    6229=>"000110110",
    6230=>"111001000",
    6231=>"000000001",
    6232=>"000000000",
    6233=>"110100100",
    6234=>"110111111",
    6235=>"000001000",
    6236=>"000110110",
    6237=>"010110100",
    6238=>"010111111",
    6239=>"111111011",
    6240=>"001011011",
    6241=>"110110111",
    6242=>"000100110",
    6243=>"111001100",
    6244=>"110101110",
    6245=>"000000001",
    6246=>"001001000",
    6247=>"111111111",
    6248=>"000100110",
    6249=>"000000000",
    6250=>"001110111",
    6251=>"000000000",
    6252=>"000100010",
    6253=>"000000000",
    6254=>"011011011",
    6255=>"100100011",
    6256=>"000110110",
    6257=>"001000001",
    6258=>"000000000",
    6259=>"100000000",
    6260=>"011111011",
    6261=>"100000100",
    6262=>"100110110",
    6263=>"001001001",
    6264=>"001001001",
    6265=>"000111011",
    6266=>"000000000",
    6267=>"100000000",
    6268=>"110110110",
    6269=>"000000000",
    6270=>"000000001",
    6271=>"001111100",
    6272=>"100000000",
    6273=>"111111111",
    6274=>"011111111",
    6275=>"111011010",
    6276=>"000100011",
    6277=>"000000001",
    6278=>"000000000",
    6279=>"011110110",
    6280=>"011111111",
    6281=>"110110000",
    6282=>"000111111",
    6283=>"001000111",
    6284=>"111011011",
    6285=>"101110010",
    6286=>"101011110",
    6287=>"001011000",
    6288=>"000111011",
    6289=>"111111000",
    6290=>"000000000",
    6291=>"101111110",
    6292=>"000000000",
    6293=>"000000000",
    6294=>"000000011",
    6295=>"110101011",
    6296=>"000001111",
    6297=>"110000010",
    6298=>"100000000",
    6299=>"010001000",
    6300=>"001000010",
    6301=>"000000000",
    6302=>"001100100",
    6303=>"000000000",
    6304=>"000000000",
    6305=>"111111000",
    6306=>"111111111",
    6307=>"000000000",
    6308=>"000000000",
    6309=>"001101011",
    6310=>"111111010",
    6311=>"110111111",
    6312=>"001101110",
    6313=>"110110110",
    6314=>"100100100",
    6315=>"000000000",
    6316=>"111011001",
    6317=>"100000000",
    6318=>"000000111",
    6319=>"000000000",
    6320=>"111111010",
    6321=>"100110111",
    6322=>"101001011",
    6323=>"111111111",
    6324=>"011111010",
    6325=>"000000001",
    6326=>"100100100",
    6327=>"101000000",
    6328=>"111111010",
    6329=>"000001111",
    6330=>"000000001",
    6331=>"111101011",
    6332=>"000001110",
    6333=>"000000000",
    6334=>"111111111",
    6335=>"000000000",
    6336=>"111111111",
    6337=>"000001111",
    6338=>"110010111",
    6339=>"110111010",
    6340=>"101000000",
    6341=>"000110000",
    6342=>"111000010",
    6343=>"100000100",
    6344=>"010011110",
    6345=>"000000011",
    6346=>"000010110",
    6347=>"100000110",
    6348=>"110110111",
    6349=>"010111111",
    6350=>"101011011",
    6351=>"000000000",
    6352=>"000110010",
    6353=>"110110100",
    6354=>"101000000",
    6355=>"110111011",
    6356=>"110110001",
    6357=>"111111000",
    6358=>"101100101",
    6359=>"000110000",
    6360=>"000000000",
    6361=>"001001011",
    6362=>"010110000",
    6363=>"001011111",
    6364=>"000000000",
    6365=>"100000000",
    6366=>"000000110",
    6367=>"000000000",
    6368=>"110110110",
    6369=>"000010000",
    6370=>"111111110",
    6371=>"000000000",
    6372=>"110111110",
    6373=>"001000000",
    6374=>"000010000",
    6375=>"111111111",
    6376=>"000001101",
    6377=>"000000101",
    6378=>"100100110",
    6379=>"001000000",
    6380=>"111110111",
    6381=>"000000000",
    6382=>"111000000",
    6383=>"001001101",
    6384=>"000000000",
    6385=>"000111111",
    6386=>"111011011",
    6387=>"011111111",
    6388=>"101000101",
    6389=>"010100000",
    6390=>"111111110",
    6391=>"000000010",
    6392=>"111111111",
    6393=>"000111111",
    6394=>"101111110",
    6395=>"011111111",
    6396=>"011110000",
    6397=>"100000001",
    6398=>"111111111",
    6399=>"111111110",
    6400=>"101001110",
    6401=>"000100111",
    6402=>"111110010",
    6403=>"111010000",
    6404=>"010000111",
    6405=>"100110111",
    6406=>"000001111",
    6407=>"111001000",
    6408=>"111100111",
    6409=>"111011000",
    6410=>"010010011",
    6411=>"100110110",
    6412=>"111100000",
    6413=>"011010000",
    6414=>"001000100",
    6415=>"111111000",
    6416=>"000110111",
    6417=>"011000000",
    6418=>"000100110",
    6419=>"100000100",
    6420=>"000100111",
    6421=>"001000000",
    6422=>"000101111",
    6423=>"100000100",
    6424=>"000110110",
    6425=>"111010000",
    6426=>"000011111",
    6427=>"001001011",
    6428=>"000010010",
    6429=>"111011000",
    6430=>"000110111",
    6431=>"000100111",
    6432=>"000100111",
    6433=>"110010111",
    6434=>"000000000",
    6435=>"001011000",
    6436=>"010100111",
    6437=>"111110000",
    6438=>"001001111",
    6439=>"000100111",
    6440=>"101111111",
    6441=>"111110000",
    6442=>"110110010",
    6443=>"000000111",
    6444=>"110010001",
    6445=>"000101011",
    6446=>"101110100",
    6447=>"010000001",
    6448=>"100000111",
    6449=>"010000000",
    6450=>"000100111",
    6451=>"000010010",
    6452=>"000000111",
    6453=>"000000010",
    6454=>"001001100",
    6455=>"000100111",
    6456=>"000011111",
    6457=>"110000011",
    6458=>"100001111",
    6459=>"100001111",
    6460=>"000100111",
    6461=>"100111100",
    6462=>"000101111",
    6463=>"101001111",
    6464=>"101111110",
    6465=>"111111111",
    6466=>"110111111",
    6467=>"000110110",
    6468=>"111111011",
    6469=>"011110110",
    6470=>"000000010",
    6471=>"111111111",
    6472=>"101111011",
    6473=>"111111111",
    6474=>"110111110",
    6475=>"001001010",
    6476=>"010111111",
    6477=>"010001011",
    6478=>"111100101",
    6479=>"000110010",
    6480=>"001000111",
    6481=>"111111010",
    6482=>"110111101",
    6483=>"111111110",
    6484=>"111101100",
    6485=>"001001000",
    6486=>"100000111",
    6487=>"110100111",
    6488=>"111110100",
    6489=>"111111010",
    6490=>"110111111",
    6491=>"001001111",
    6492=>"111111111",
    6493=>"010111010",
    6494=>"010010111",
    6495=>"100100111",
    6496=>"101001001",
    6497=>"111111011",
    6498=>"111111111",
    6499=>"100001111",
    6500=>"111111111",
    6501=>"111111111",
    6502=>"111111011",
    6503=>"111111111",
    6504=>"101101100",
    6505=>"000000000",
    6506=>"011000100",
    6507=>"111110111",
    6508=>"101101001",
    6509=>"111111011",
    6510=>"000111110",
    6511=>"000000001",
    6512=>"010111111",
    6513=>"111101001",
    6514=>"111111111",
    6515=>"000010001",
    6516=>"000000001",
    6517=>"001101111",
    6518=>"001001011",
    6519=>"000000000",
    6520=>"101000000",
    6521=>"100100001",
    6522=>"100101101",
    6523=>"111101001",
    6524=>"110000110",
    6525=>"011011111",
    6526=>"111111011",
    6527=>"111001001",
    6528=>"101100100",
    6529=>"000000000",
    6530=>"111111111",
    6531=>"110110110",
    6532=>"111111111",
    6533=>"001001111",
    6534=>"000000000",
    6535=>"110111110",
    6536=>"111111111",
    6537=>"110000000",
    6538=>"000000000",
    6539=>"111111111",
    6540=>"000100111",
    6541=>"111010011",
    6542=>"111111111",
    6543=>"111111011",
    6544=>"001000000",
    6545=>"111011101",
    6546=>"111101100",
    6547=>"001000000",
    6548=>"111101100",
    6549=>"111111000",
    6550=>"000000111",
    6551=>"001000100",
    6552=>"100110111",
    6553=>"110010011",
    6554=>"110010000",
    6555=>"001000000",
    6556=>"111111011",
    6557=>"110111111",
    6558=>"000000000",
    6559=>"010011010",
    6560=>"001100100",
    6561=>"111111111",
    6562=>"000001100",
    6563=>"000000110",
    6564=>"000000000",
    6565=>"111111111",
    6566=>"000000000",
    6567=>"111111111",
    6568=>"010001001",
    6569=>"111111110",
    6570=>"011001101",
    6571=>"001000000",
    6572=>"111111111",
    6573=>"000000000",
    6574=>"100110111",
    6575=>"001000000",
    6576=>"111111010",
    6577=>"111011000",
    6578=>"000000100",
    6579=>"011010101",
    6580=>"111110100",
    6581=>"000000000",
    6582=>"111111111",
    6583=>"011001001",
    6584=>"001001000",
    6585=>"100110011",
    6586=>"000000000",
    6587=>"000000000",
    6588=>"111111111",
    6589=>"111111111",
    6590=>"000000000",
    6591=>"001100100",
    6592=>"010010100",
    6593=>"000001000",
    6594=>"000010011",
    6595=>"000011111",
    6596=>"001100111",
    6597=>"111001110",
    6598=>"000111111",
    6599=>"110110110",
    6600=>"001001011",
    6601=>"000000010",
    6602=>"000001111",
    6603=>"011010110",
    6604=>"110000111",
    6605=>"000000010",
    6606=>"110111001",
    6607=>"001001111",
    6608=>"011111111",
    6609=>"000111000",
    6610=>"100001001",
    6611=>"001010110",
    6612=>"111000000",
    6613=>"000000000",
    6614=>"111101000",
    6615=>"010110110",
    6616=>"111000000",
    6617=>"000111111",
    6618=>"111100110",
    6619=>"000110010",
    6620=>"110111111",
    6621=>"000111111",
    6622=>"000111011",
    6623=>"000111111",
    6624=>"111101000",
    6625=>"011001110",
    6626=>"100111110",
    6627=>"010101000",
    6628=>"000000000",
    6629=>"100001001",
    6630=>"111000111",
    6631=>"000000110",
    6632=>"000110110",
    6633=>"000000111",
    6634=>"010110100",
    6635=>"110111111",
    6636=>"000000000",
    6637=>"100001000",
    6638=>"111101000",
    6639=>"011110110",
    6640=>"000011111",
    6641=>"000111111",
    6642=>"111001001",
    6643=>"111111110",
    6644=>"000000111",
    6645=>"011011111",
    6646=>"100000111",
    6647=>"111000000",
    6648=>"100001000",
    6649=>"110000011",
    6650=>"010111110",
    6651=>"010110111",
    6652=>"111011000",
    6653=>"101000000",
    6654=>"000000000",
    6655=>"110111100",
    6656=>"100000010",
    6657=>"001111101",
    6658=>"111111111",
    6659=>"110000100",
    6660=>"000000111",
    6661=>"000000000",
    6662=>"111111111",
    6663=>"000000000",
    6664=>"010000000",
    6665=>"110010010",
    6666=>"111111111",
    6667=>"101011010",
    6668=>"111101111",
    6669=>"111110111",
    6670=>"010101001",
    6671=>"000000000",
    6672=>"100001000",
    6673=>"000001100",
    6674=>"111111111",
    6675=>"111111111",
    6676=>"111100101",
    6677=>"000000000",
    6678=>"001101101",
    6679=>"011100100",
    6680=>"011111110",
    6681=>"001111100",
    6682=>"101111101",
    6683=>"100110111",
    6684=>"000111110",
    6685=>"111000010",
    6686=>"000000000",
    6687=>"000001111",
    6688=>"111000011",
    6689=>"001000000",
    6690=>"000000100",
    6691=>"001000100",
    6692=>"000000000",
    6693=>"111010011",
    6694=>"001111111",
    6695=>"111110111",
    6696=>"110010010",
    6697=>"000000000",
    6698=>"001110010",
    6699=>"011101101",
    6700=>"110111111",
    6701=>"111001010",
    6702=>"111000011",
    6703=>"010001011",
    6704=>"000101111",
    6705=>"010110001",
    6706=>"001000011",
    6707=>"010110111",
    6708=>"000101101",
    6709=>"000000101",
    6710=>"010000000",
    6711=>"111100100",
    6712=>"000111101",
    6713=>"111010111",
    6714=>"000000000",
    6715=>"111000100",
    6716=>"000001000",
    6717=>"100000000",
    6718=>"000000000",
    6719=>"000010100",
    6720=>"001001011",
    6721=>"111111111",
    6722=>"000000000",
    6723=>"110110100",
    6724=>"000000000",
    6725=>"011000110",
    6726=>"110110000",
    6727=>"000111001",
    6728=>"010010000",
    6729=>"001001111",
    6730=>"000000000",
    6731=>"001000101",
    6732=>"111101100",
    6733=>"110100101",
    6734=>"001001101",
    6735=>"000100000",
    6736=>"000000000",
    6737=>"110110110",
    6738=>"001101101",
    6739=>"100011111",
    6740=>"110100111",
    6741=>"000000111",
    6742=>"011011111",
    6743=>"001000111",
    6744=>"111110000",
    6745=>"000001001",
    6746=>"000000000",
    6747=>"001001111",
    6748=>"000100111",
    6749=>"111111110",
    6750=>"010001001",
    6751=>"000000001",
    6752=>"000000000",
    6753=>"000000000",
    6754=>"000100101",
    6755=>"111110000",
    6756=>"001111111",
    6757=>"000010000",
    6758=>"100000001",
    6759=>"111111111",
    6760=>"000000000",
    6761=>"110100100",
    6762=>"110100111",
    6763=>"111111111",
    6764=>"101001111",
    6765=>"000001001",
    6766=>"000000001",
    6767=>"001001011",
    6768=>"111011111",
    6769=>"100001111",
    6770=>"100000100",
    6771=>"101101011",
    6772=>"101000001",
    6773=>"001001011",
    6774=>"000000000",
    6775=>"111110000",
    6776=>"101001111",
    6777=>"001101011",
    6778=>"000001010",
    6779=>"000001010",
    6780=>"000100000",
    6781=>"110111010",
    6782=>"111111011",
    6783=>"000001001",
    6784=>"100100100",
    6785=>"100100100",
    6786=>"110100110",
    6787=>"000001111",
    6788=>"101101101",
    6789=>"001001001",
    6790=>"001010100",
    6791=>"001001000",
    6792=>"010011001",
    6793=>"111011000",
    6794=>"111000101",
    6795=>"111111111",
    6796=>"111110111",
    6797=>"101001100",
    6798=>"000000000",
    6799=>"001010010",
    6800=>"001001001",
    6801=>"101011001",
    6802=>"111001001",
    6803=>"111011111",
    6804=>"100000011",
    6805=>"001001011",
    6806=>"000001111",
    6807=>"011111111",
    6808=>"100000011",
    6809=>"110100100",
    6810=>"011011101",
    6811=>"100000000",
    6812=>"001001011",
    6813=>"010011011",
    6814=>"000101011",
    6815=>"100001011",
    6816=>"001001011",
    6817=>"001101001",
    6818=>"001101111",
    6819=>"100101111",
    6820=>"000000101",
    6821=>"100000010",
    6822=>"110011111",
    6823=>"110110100",
    6824=>"010010110",
    6825=>"111110100",
    6826=>"001000000",
    6827=>"000000100",
    6828=>"111110101",
    6829=>"001001001",
    6830=>"001001111",
    6831=>"001001011",
    6832=>"110110100",
    6833=>"000000000",
    6834=>"000001011",
    6835=>"000001100",
    6836=>"010100111",
    6837=>"110100111",
    6838=>"111110110",
    6839=>"100100000",
    6840=>"100000000",
    6841=>"111111111",
    6842=>"101000000",
    6843=>"111110111",
    6844=>"000001011",
    6845=>"100000001",
    6846=>"011110110",
    6847=>"110100100",
    6848=>"001100110",
    6849=>"111011101",
    6850=>"000000111",
    6851=>"111011000",
    6852=>"001001011",
    6853=>"000101001",
    6854=>"000000111",
    6855=>"111100111",
    6856=>"001001111",
    6857=>"111000000",
    6858=>"100100111",
    6859=>"000001011",
    6860=>"111101101",
    6861=>"000011000",
    6862=>"000000111",
    6863=>"010000100",
    6864=>"000010010",
    6865=>"011111000",
    6866=>"001001111",
    6867=>"010010010",
    6868=>"000011011",
    6869=>"000000111",
    6870=>"011111100",
    6871=>"011110000",
    6872=>"101101101",
    6873=>"100000010",
    6874=>"011111100",
    6875=>"100000111",
    6876=>"101000011",
    6877=>"111111000",
    6878=>"000000101",
    6879=>"000010111",
    6880=>"001001011",
    6881=>"000001011",
    6882=>"111011001",
    6883=>"000000100",
    6884=>"101111000",
    6885=>"100100011",
    6886=>"011110100",
    6887=>"000011111",
    6888=>"000000111",
    6889=>"000000011",
    6890=>"001011011",
    6891=>"110111000",
    6892=>"100000011",
    6893=>"000110111",
    6894=>"011101101",
    6895=>"010110111",
    6896=>"111000001",
    6897=>"000000101",
    6898=>"010011111",
    6899=>"000110111",
    6900=>"000010111",
    6901=>"000100111",
    6902=>"000001011",
    6903=>"001101000",
    6904=>"011010100",
    6905=>"000110110",
    6906=>"000010111",
    6907=>"000110111",
    6908=>"011111001",
    6909=>"110000000",
    6910=>"000000011",
    6911=>"010010010",
    6912=>"111111111",
    6913=>"000000000",
    6914=>"111111011",
    6915=>"010110010",
    6916=>"111111110",
    6917=>"000000000",
    6918=>"000100010",
    6919=>"110001011",
    6920=>"100000001",
    6921=>"000000000",
    6922=>"111011110",
    6923=>"111111111",
    6924=>"111110110",
    6925=>"000000000",
    6926=>"111110111",
    6927=>"100100110",
    6928=>"000000001",
    6929=>"011001000",
    6930=>"111101110",
    6931=>"000000100",
    6932=>"011011001",
    6933=>"110110011",
    6934=>"111111111",
    6935=>"101000000",
    6936=>"000000000",
    6937=>"111111010",
    6938=>"000000000",
    6939=>"011000010",
    6940=>"000010000",
    6941=>"111111000",
    6942=>"000000000",
    6943=>"100000111",
    6944=>"000000000",
    6945=>"000100000",
    6946=>"000000000",
    6947=>"000100111",
    6948=>"000000000",
    6949=>"111111111",
    6950=>"001001000",
    6951=>"111111111",
    6952=>"111111111",
    6953=>"000000000",
    6954=>"010000000",
    6955=>"100000000",
    6956=>"111111011",
    6957=>"010110111",
    6958=>"000000000",
    6959=>"110001101",
    6960=>"011011011",
    6961=>"000000000",
    6962=>"001001010",
    6963=>"000001000",
    6964=>"010110110",
    6965=>"111111111",
    6966=>"111111111",
    6967=>"010000011",
    6968=>"000000101",
    6969=>"010111111",
    6970=>"110101100",
    6971=>"111111111",
    6972=>"111111111",
    6973=>"100001101",
    6974=>"111011111",
    6975=>"100100100",
    6976=>"110111111",
    6977=>"000000100",
    6978=>"000000000",
    6979=>"111001111",
    6980=>"000000100",
    6981=>"011011000",
    6982=>"000000000",
    6983=>"111111011",
    6984=>"000000000",
    6985=>"000101111",
    6986=>"000000000",
    6987=>"101100110",
    6988=>"111100110",
    6989=>"111010111",
    6990=>"001000111",
    6991=>"111010001",
    6992=>"101101011",
    6993=>"111011000",
    6994=>"110101110",
    6995=>"101000001",
    6996=>"111111111",
    6997=>"000100100",
    6998=>"111111100",
    6999=>"101101110",
    7000=>"010111110",
    7001=>"000001111",
    7002=>"111111100",
    7003=>"000011011",
    7004=>"000111001",
    7005=>"111001001",
    7006=>"000000000",
    7007=>"000110000",
    7008=>"111100000",
    7009=>"000000100",
    7010=>"101101110",
    7011=>"111110000",
    7012=>"011111100",
    7013=>"011000010",
    7014=>"100000001",
    7015=>"000000000",
    7016=>"000000000",
    7017=>"111001101",
    7018=>"000110000",
    7019=>"111101111",
    7020=>"100100110",
    7021=>"100111111",
    7022=>"111111111",
    7023=>"001111111",
    7024=>"000000000",
    7025=>"000111110",
    7026=>"110111110",
    7027=>"000010010",
    7028=>"000000001",
    7029=>"000001110",
    7030=>"110110010",
    7031=>"111001111",
    7032=>"101001100",
    7033=>"111101110",
    7034=>"100101000",
    7035=>"010010010",
    7036=>"111000000",
    7037=>"001101000",
    7038=>"000000100",
    7039=>"001101111",
    7040=>"010110110",
    7041=>"000011110",
    7042=>"110110000",
    7043=>"100100111",
    7044=>"001100111",
    7045=>"100110111",
    7046=>"101111011",
    7047=>"100000100",
    7048=>"111110110",
    7049=>"011010100",
    7050=>"111101001",
    7051=>"001001100",
    7052=>"111110110",
    7053=>"011100110",
    7054=>"001010000",
    7055=>"000000011",
    7056=>"000101011",
    7057=>"100100000",
    7058=>"100100111",
    7059=>"110111000",
    7060=>"101000000",
    7061=>"010010000",
    7062=>"010011010",
    7063=>"000011011",
    7064=>"100100100",
    7065=>"111010000",
    7066=>"100101101",
    7067=>"100110111",
    7068=>"101111111",
    7069=>"100100111",
    7070=>"110110110",
    7071=>"000010000",
    7072=>"100000001",
    7073=>"110111111",
    7074=>"100100011",
    7075=>"100000001",
    7076=>"000111110",
    7077=>"110000001",
    7078=>"001011011",
    7079=>"111011001",
    7080=>"100101100",
    7081=>"000000000",
    7082=>"001001000",
    7083=>"000100111",
    7084=>"101101000",
    7085=>"011100001",
    7086=>"100010011",
    7087=>"010000110",
    7088=>"110100111",
    7089=>"111000000",
    7090=>"101100000",
    7091=>"000011011",
    7092=>"110110100",
    7093=>"100100111",
    7094=>"101001111",
    7095=>"001000000",
    7096=>"010010000",
    7097=>"110100000",
    7098=>"000001000",
    7099=>"110011100",
    7100=>"000000011",
    7101=>"100000000",
    7102=>"011110110",
    7103=>"100100111",
    7104=>"000000001",
    7105=>"001011001",
    7106=>"110111111",
    7107=>"101111101",
    7108=>"100111101",
    7109=>"001111000",
    7110=>"011001011",
    7111=>"110110101",
    7112=>"110111001",
    7113=>"000000111",
    7114=>"100100100",
    7115=>"000111011",
    7116=>"100100101",
    7117=>"000000001",
    7118=>"100111100",
    7119=>"000100000",
    7120=>"000001001",
    7121=>"101101101",
    7122=>"001100010",
    7123=>"011000011",
    7124=>"000110010",
    7125=>"001001001",
    7126=>"101101111",
    7127=>"001001001",
    7128=>"000001110",
    7129=>"111101100",
    7130=>"001001000",
    7131=>"111001100",
    7132=>"001001001",
    7133=>"100110110",
    7134=>"011011011",
    7135=>"001001001",
    7136=>"110100000",
    7137=>"001000111",
    7138=>"001001110",
    7139=>"100100110",
    7140=>"000110101",
    7141=>"100110111",
    7142=>"011010000",
    7143=>"001010110",
    7144=>"011010001",
    7145=>"001001000",
    7146=>"001001100",
    7147=>"110001000",
    7148=>"111011001",
    7149=>"001001000",
    7150=>"110110110",
    7151=>"111011001",
    7152=>"111100000",
    7153=>"001001001",
    7154=>"000001000",
    7155=>"011011001",
    7156=>"011001001",
    7157=>"111100000",
    7158=>"000000000",
    7159=>"100110011",
    7160=>"011001001",
    7161=>"110111001",
    7162=>"011001001",
    7163=>"110001001",
    7164=>"110100110",
    7165=>"110000000",
    7166=>"011110000",
    7167=>"001001001",
    7168=>"000000000",
    7169=>"000000111",
    7170=>"000001010",
    7171=>"011001001",
    7172=>"011111110",
    7173=>"001000010",
    7174=>"011111111",
    7175=>"000100000",
    7176=>"011111111",
    7177=>"010000011",
    7178=>"110111011",
    7179=>"001001100",
    7180=>"111101001",
    7181=>"101010111",
    7182=>"001001100",
    7183=>"100000101",
    7184=>"000000000",
    7185=>"111111101",
    7186=>"001001000",
    7187=>"111111111",
    7188=>"001001110",
    7189=>"111111110",
    7190=>"111111111",
    7191=>"110010111",
    7192=>"000000000",
    7193=>"111100000",
    7194=>"000000000",
    7195=>"100100001",
    7196=>"001001101",
    7197=>"011011101",
    7198=>"001111110",
    7199=>"101101111",
    7200=>"000000110",
    7201=>"111111111",
    7202=>"011000110",
    7203=>"001000000",
    7204=>"111111111",
    7205=>"000000000",
    7206=>"110110011",
    7207=>"111011111",
    7208=>"000010100",
    7209=>"000000000",
    7210=>"001011111",
    7211=>"110100001",
    7212=>"000000000",
    7213=>"100100011",
    7214=>"001000110",
    7215=>"101100011",
    7216=>"111111101",
    7217=>"111110010",
    7218=>"000000000",
    7219=>"111111111",
    7220=>"000000100",
    7221=>"110111111",
    7222=>"100011111",
    7223=>"101111111",
    7224=>"111101111",
    7225=>"001100100",
    7226=>"100100100",
    7227=>"100100010",
    7228=>"101111111",
    7229=>"000100000",
    7230=>"111110111",
    7231=>"111000000",
    7232=>"100110110",
    7233=>"100010000",
    7234=>"000111001",
    7235=>"000111111",
    7236=>"010011001",
    7237=>"011000110",
    7238=>"011011100",
    7239=>"100111011",
    7240=>"011001000",
    7241=>"100011000",
    7242=>"100100000",
    7243=>"010011000",
    7244=>"110111111",
    7245=>"001000000",
    7246=>"010011100",
    7247=>"011111101",
    7248=>"111011000",
    7249=>"111001100",
    7250=>"100111111",
    7251=>"000000100",
    7252=>"001110010",
    7253=>"000111000",
    7254=>"111000000",
    7255=>"110011000",
    7256=>"110110011",
    7257=>"100100110",
    7258=>"110100101",
    7259=>"111000000",
    7260=>"111001001",
    7261=>"001000111",
    7262=>"110011110",
    7263=>"010001001",
    7264=>"000111011",
    7265=>"110000000",
    7266=>"110110000",
    7267=>"000000100",
    7268=>"000100111",
    7269=>"000111101",
    7270=>"101100100",
    7271=>"000000010",
    7272=>"100111111",
    7273=>"010000000",
    7274=>"111110000",
    7275=>"100110110",
    7276=>"001101110",
    7277=>"100110000",
    7278=>"001001001",
    7279=>"100000000",
    7280=>"111011000",
    7281=>"001100000",
    7282=>"011001000",
    7283=>"111011010",
    7284=>"111011000",
    7285=>"000111111",
    7286=>"111011001",
    7287=>"000110111",
    7288=>"111111000",
    7289=>"101011000",
    7290=>"000110110",
    7291=>"000110011",
    7292=>"110100111",
    7293=>"000000011",
    7294=>"000000000",
    7295=>"000100010",
    7296=>"110001110",
    7297=>"000101000",
    7298=>"111101010",
    7299=>"101001001",
    7300=>"100000100",
    7301=>"000000001",
    7302=>"000000100",
    7303=>"011010110",
    7304=>"001101000",
    7305=>"010110110",
    7306=>"000011000",
    7307=>"111101111",
    7308=>"010000111",
    7309=>"101111101",
    7310=>"100111010",
    7311=>"001001001",
    7312=>"001001000",
    7313=>"101101001",
    7314=>"100101111",
    7315=>"101101000",
    7316=>"111101000",
    7317=>"000100110",
    7318=>"001001001",
    7319=>"001000000",
    7320=>"111000111",
    7321=>"001000101",
    7322=>"000000101",
    7323=>"010111011",
    7324=>"010001010",
    7325=>"100000101",
    7326=>"001001101",
    7327=>"110111111",
    7328=>"110111110",
    7329=>"011001001",
    7330=>"101001101",
    7331=>"101001001",
    7332=>"011000001",
    7333=>"110010011",
    7334=>"101000000",
    7335=>"100101100",
    7336=>"111111111",
    7337=>"000000100",
    7338=>"000011110",
    7339=>"001101101",
    7340=>"111011011",
    7341=>"110111101",
    7342=>"111010110",
    7343=>"111011010",
    7344=>"000001111",
    7345=>"001011000",
    7346=>"101101110",
    7347=>"011010010",
    7348=>"000000000",
    7349=>"010100100",
    7350=>"100100100",
    7351=>"000000000",
    7352=>"000000001",
    7353=>"110110110",
    7354=>"001111111",
    7355=>"011011101",
    7356=>"001001001",
    7357=>"011101100",
    7358=>"011000001",
    7359=>"000000000",
    7360=>"111101001",
    7361=>"000000000",
    7362=>"000000000",
    7363=>"000100110",
    7364=>"110100110",
    7365=>"111100111",
    7366=>"100011010",
    7367=>"111111001",
    7368=>"000000000",
    7369=>"011111010",
    7370=>"111011011",
    7371=>"001100100",
    7372=>"000000000",
    7373=>"111111101",
    7374=>"111001000",
    7375=>"100011110",
    7376=>"111101111",
    7377=>"001111011",
    7378=>"111111111",
    7379=>"110001011",
    7380=>"111111111",
    7381=>"011101010",
    7382=>"110100101",
    7383=>"001000101",
    7384=>"000000000",
    7385=>"111111010",
    7386=>"110101011",
    7387=>"001011111",
    7388=>"111011011",
    7389=>"111111000",
    7390=>"000000000",
    7391=>"001110111",
    7392=>"010100001",
    7393=>"101100110",
    7394=>"100110100",
    7395=>"110001010",
    7396=>"111111111",
    7397=>"111111100",
    7398=>"010111111",
    7399=>"000000000",
    7400=>"000000000",
    7401=>"001010000",
    7402=>"001000000",
    7403=>"111111111",
    7404=>"100110001",
    7405=>"110000001",
    7406=>"000100001",
    7407=>"011111111",
    7408=>"010111011",
    7409=>"101000000",
    7410=>"011101101",
    7411=>"001000101",
    7412=>"100101111",
    7413=>"111111111",
    7414=>"111101110",
    7415=>"000000000",
    7416=>"100001010",
    7417=>"100101111",
    7418=>"111110111",
    7419=>"000000001",
    7420=>"000000000",
    7421=>"110000001",
    7422=>"000000000",
    7423=>"001000001",
    7424=>"001100000",
    7425=>"111101111",
    7426=>"111101111",
    7427=>"101101001",
    7428=>"001100010",
    7429=>"111101000",
    7430=>"111111111",
    7431=>"001000000",
    7432=>"110111111",
    7433=>"000000000",
    7434=>"000011011",
    7435=>"111001000",
    7436=>"111101111",
    7437=>"111000110",
    7438=>"100110111",
    7439=>"111110101",
    7440=>"111110010",
    7441=>"001000000",
    7442=>"111111011",
    7443=>"111000101",
    7444=>"100001000",
    7445=>"100000000",
    7446=>"111101111",
    7447=>"111011011",
    7448=>"111111111",
    7449=>"000000000",
    7450=>"001100001",
    7451=>"101010000",
    7452=>"000000101",
    7453=>"000000000",
    7454=>"101111111",
    7455=>"000000000",
    7456=>"111111111",
    7457=>"010011000",
    7458=>"001010000",
    7459=>"000000000",
    7460=>"000000000",
    7461=>"000000000",
    7462=>"011010000",
    7463=>"111101111",
    7464=>"111011111",
    7465=>"111111111",
    7466=>"001111110",
    7467=>"011000000",
    7468=>"111101101",
    7469=>"111110111",
    7470=>"111111111",
    7471=>"111110111",
    7472=>"000011000",
    7473=>"001000000",
    7474=>"101101101",
    7475=>"000000000",
    7476=>"101111100",
    7477=>"001001001",
    7478=>"000001000",
    7479=>"111111111",
    7480=>"110011111",
    7481=>"111001100",
    7482=>"001010000",
    7483=>"101101110",
    7484=>"111111111",
    7485=>"000000000",
    7486=>"111111111",
    7487=>"111000101",
    7488=>"000000010",
    7489=>"110000110",
    7490=>"000011001",
    7491=>"111111111",
    7492=>"010011001",
    7493=>"111011000",
    7494=>"011110011",
    7495=>"111111111",
    7496=>"111010001",
    7497=>"000100101",
    7498=>"000110100",
    7499=>"011011001",
    7500=>"000010110",
    7501=>"000000010",
    7502=>"010011001",
    7503=>"111111111",
    7504=>"110111111",
    7505=>"111111100",
    7506=>"110011001",
    7507=>"011111100",
    7508=>"011001001",
    7509=>"000000000",
    7510=>"000111000",
    7511=>"111111000",
    7512=>"101111111",
    7513=>"111000000",
    7514=>"111111110",
    7515=>"100110000",
    7516=>"011110010",
    7517=>"101001111",
    7518=>"111011000",
    7519=>"111110000",
    7520=>"010011111",
    7521=>"000011011",
    7522=>"011001010",
    7523=>"001001111",
    7524=>"110111111",
    7525=>"011111111",
    7526=>"011110110",
    7527=>"000010011",
    7528=>"000000111",
    7529=>"111000000",
    7530=>"011111001",
    7531=>"111111101",
    7532=>"000000000",
    7533=>"100100100",
    7534=>"000101001",
    7535=>"000000100",
    7536=>"111000000",
    7537=>"111100000",
    7538=>"111111111",
    7539=>"000000010",
    7540=>"000000111",
    7541=>"000100000",
    7542=>"000000000",
    7543=>"000011111",
    7544=>"110111000",
    7545=>"110101000",
    7546=>"011110111",
    7547=>"000100100",
    7548=>"111111000",
    7549=>"111010101",
    7550=>"000100110",
    7551=>"110110010",
    7552=>"000011111",
    7553=>"111111000",
    7554=>"000101111",
    7555=>"011111111",
    7556=>"000100110",
    7557=>"111001100",
    7558=>"011111100",
    7559=>"000000111",
    7560=>"011011000",
    7561=>"101001101",
    7562=>"000111101",
    7563=>"000001110",
    7564=>"111111111",
    7565=>"100111001",
    7566=>"010000101",
    7567=>"000000111",
    7568=>"101111111",
    7569=>"111000000",
    7570=>"111011011",
    7571=>"000000111",
    7572=>"000000001",
    7573=>"110000000",
    7574=>"111111000",
    7575=>"111111000",
    7576=>"010111010",
    7577=>"010000000",
    7578=>"111100011",
    7579=>"101111000",
    7580=>"000010111",
    7581=>"111000000",
    7582=>"111111000",
    7583=>"000111011",
    7584=>"000000111",
    7585=>"111000000",
    7586=>"011000011",
    7587=>"100000111",
    7588=>"111000111",
    7589=>"000000111",
    7590=>"111100000",
    7591=>"000100111",
    7592=>"000111010",
    7593=>"000000101",
    7594=>"001000110",
    7595=>"010000110",
    7596=>"000111110",
    7597=>"000000010",
    7598=>"000000111",
    7599=>"110111000",
    7600=>"000111110",
    7601=>"000001000",
    7602=>"011101111",
    7603=>"101001100",
    7604=>"011111000",
    7605=>"000010011",
    7606=>"000000011",
    7607=>"010000101",
    7608=>"111101000",
    7609=>"000001111",
    7610=>"000000100",
    7611=>"000000111",
    7612=>"010000000",
    7613=>"111100100",
    7614=>"000010100",
    7615=>"110010000",
    7616=>"000000010",
    7617=>"100100000",
    7618=>"000001010",
    7619=>"110011001",
    7620=>"000011011",
    7621=>"000011111",
    7622=>"011110000",
    7623=>"111101000",
    7624=>"000011111",
    7625=>"001000111",
    7626=>"111110000",
    7627=>"000000111",
    7628=>"110011111",
    7629=>"100000000",
    7630=>"001000111",
    7631=>"010000000",
    7632=>"001100001",
    7633=>"110110000",
    7634=>"111111110",
    7635=>"011111100",
    7636=>"001011010",
    7637=>"000010100",
    7638=>"111100110",
    7639=>"011110000",
    7640=>"000001111",
    7641=>"011110001",
    7642=>"111100000",
    7643=>"111110000",
    7644=>"010100001",
    7645=>"000001111",
    7646=>"000011111",
    7647=>"001110100",
    7648=>"111011110",
    7649=>"001011000",
    7650=>"111000001",
    7651=>"100000001",
    7652=>"011100000",
    7653=>"000001111",
    7654=>"110100000",
    7655=>"111011110",
    7656=>"000100000",
    7657=>"001110000",
    7658=>"000011110",
    7659=>"001010100",
    7660=>"000110100",
    7661=>"011110000",
    7662=>"100001111",
    7663=>"001100000",
    7664=>"110110000",
    7665=>"010100001",
    7666=>"000001111",
    7667=>"111110000",
    7668=>"111100000",
    7669=>"011100000",
    7670=>"011100100",
    7671=>"100001111",
    7672=>"011110000",
    7673=>"001000000",
    7674=>"011010100",
    7675=>"011110100",
    7676=>"111111000",
    7677=>"000001011",
    7678=>"011000000",
    7679=>"111100000",
    7680=>"100100011",
    7681=>"010110001",
    7682=>"010010111",
    7683=>"111011000",
    7684=>"111101111",
    7685=>"100000111",
    7686=>"010010000",
    7687=>"100110110",
    7688=>"000000000",
    7689=>"110100001",
    7690=>"110010111",
    7691=>"111111111",
    7692=>"111000111",
    7693=>"010110111",
    7694=>"000000000",
    7695=>"010111011",
    7696=>"000100110",
    7697=>"010000100",
    7698=>"011100111",
    7699=>"110000001",
    7700=>"010000100",
    7701=>"111100000",
    7702=>"100110111",
    7703=>"000000000",
    7704=>"000000100",
    7705=>"001000001",
    7706=>"101000111",
    7707=>"100000100",
    7708=>"111011000",
    7709=>"000000000",
    7710=>"000010000",
    7711=>"000110111",
    7712=>"110100110",
    7713=>"011001100",
    7714=>"011111111",
    7715=>"000000100",
    7716=>"001000110",
    7717=>"010010010",
    7718=>"010000000",
    7719=>"001110000",
    7720=>"100011111",
    7721=>"111110000",
    7722=>"111001100",
    7723=>"010100011",
    7724=>"110001010",
    7725=>"111011100",
    7726=>"100110111",
    7727=>"011011010",
    7728=>"111111001",
    7729=>"110100110",
    7730=>"111001001",
    7731=>"111110010",
    7732=>"000100111",
    7733=>"000001110",
    7734=>"011010100",
    7735=>"000000110",
    7736=>"111111111",
    7737=>"110000000",
    7738=>"010000000",
    7739=>"000010011",
    7740=>"101000011",
    7741=>"110010000",
    7742=>"010011000",
    7743=>"000110111",
    7744=>"000001001",
    7745=>"001000010",
    7746=>"011111111",
    7747=>"000001110",
    7748=>"000110010",
    7749=>"111000000",
    7750=>"101000110",
    7751=>"000111111",
    7752=>"000111111",
    7753=>"000000101",
    7754=>"000111110",
    7755=>"001111110",
    7756=>"000111111",
    7757=>"011001111",
    7758=>"000000111",
    7759=>"000111111",
    7760=>"111000000",
    7761=>"111100000",
    7762=>"001001000",
    7763=>"111100100",
    7764=>"111100011",
    7765=>"111010000",
    7766=>"111000000",
    7767=>"111000000",
    7768=>"110000000",
    7769=>"111000010",
    7770=>"110000000",
    7771=>"110000000",
    7772=>"111000101",
    7773=>"000111111",
    7774=>"001000010",
    7775=>"001000000",
    7776=>"000111111",
    7777=>"111010000",
    7778=>"111000000",
    7779=>"000111111",
    7780=>"101000000",
    7781=>"000111111",
    7782=>"111110000",
    7783=>"000000001",
    7784=>"111111111",
    7785=>"000000111",
    7786=>"111000000",
    7787=>"111110001",
    7788=>"000000100",
    7789=>"110000100",
    7790=>"000111111",
    7791=>"011010010",
    7792=>"111000011",
    7793=>"111000000",
    7794=>"101001010",
    7795=>"110110110",
    7796=>"111010000",
    7797=>"000000100",
    7798=>"100111111",
    7799=>"000110111",
    7800=>"111000000",
    7801=>"000101111",
    7802=>"100101110",
    7803=>"000001111",
    7804=>"010110010",
    7805=>"000111101",
    7806=>"000011111",
    7807=>"111000000",
    7808=>"111111111",
    7809=>"110111101",
    7810=>"000000010",
    7811=>"101001010",
    7812=>"111011011",
    7813=>"111011100",
    7814=>"000000000",
    7815=>"011000111",
    7816=>"111011000",
    7817=>"111010010",
    7818=>"001010110",
    7819=>"000111000",
    7820=>"111100111",
    7821=>"110111111",
    7822=>"011001011",
    7823=>"001000000",
    7824=>"001100111",
    7825=>"100111001",
    7826=>"000000000",
    7827=>"000000000",
    7828=>"011000101",
    7829=>"000000000",
    7830=>"100101101",
    7831=>"001000000",
    7832=>"010111011",
    7833=>"110111000",
    7834=>"100000000",
    7835=>"001101100",
    7836=>"001011000",
    7837=>"100000000",
    7838=>"111111111",
    7839=>"110000101",
    7840=>"000000111",
    7841=>"110111111",
    7842=>"111111111",
    7843=>"001000111",
    7844=>"111000111",
    7845=>"000000000",
    7846=>"000000010",
    7847=>"000000000",
    7848=>"011010111",
    7849=>"101000100",
    7850=>"101101101",
    7851=>"010101001",
    7852=>"000000010",
    7853=>"111010110",
    7854=>"011000111",
    7855=>"001000000",
    7856=>"000111101",
    7857=>"000011100",
    7858=>"000110001",
    7859=>"011011110",
    7860=>"001001111",
    7861=>"011111111",
    7862=>"011010110",
    7863=>"111001111",
    7864=>"101111010",
    7865=>"001010110",
    7866=>"111101111",
    7867=>"111000111",
    7868=>"000000000",
    7869=>"100100000",
    7870=>"111111111",
    7871=>"000111011",
    7872=>"101001011",
    7873=>"111111111",
    7874=>"000000000",
    7875=>"100111000",
    7876=>"000110110",
    7877=>"110111001",
    7878=>"101110110",
    7879=>"000001001",
    7880=>"001000100",
    7881=>"000000001",
    7882=>"010000001",
    7883=>"110000011",
    7884=>"111101000",
    7885=>"010001000",
    7886=>"010000000",
    7887=>"000000110",
    7888=>"000001011",
    7889=>"000111111",
    7890=>"111000100",
    7891=>"000010110",
    7892=>"101100111",
    7893=>"110110111",
    7894=>"111111111",
    7895=>"111111011",
    7896=>"000010101",
    7897=>"010110000",
    7898=>"001010100",
    7899=>"011001111",
    7900=>"111111000",
    7901=>"000000001",
    7902=>"111011011",
    7903=>"111101000",
    7904=>"000000001",
    7905=>"011111011",
    7906=>"000000101",
    7907=>"000100000",
    7908=>"100101111",
    7909=>"001000100",
    7910=>"111010110",
    7911=>"010000100",
    7912=>"000000000",
    7913=>"010000000",
    7914=>"010100000",
    7915=>"111111100",
    7916=>"111100111",
    7917=>"111001010",
    7918=>"000000000",
    7919=>"100111110",
    7920=>"000111010",
    7921=>"000101111",
    7922=>"000000110",
    7923=>"111111010",
    7924=>"111111111",
    7925=>"111001111",
    7926=>"011111011",
    7927=>"000000000",
    7928=>"110111111",
    7929=>"000001011",
    7930=>"010000001",
    7931=>"000000101",
    7932=>"110111111",
    7933=>"000000011",
    7934=>"000000000",
    7935=>"000011111",
    7936=>"110110110",
    7937=>"100110110",
    7938=>"011011011",
    7939=>"101001001",
    7940=>"011011011",
    7941=>"101101101",
    7942=>"101000011",
    7943=>"001001001",
    7944=>"111011111",
    7945=>"010011001",
    7946=>"011011011",
    7947=>"010010011",
    7948=>"111111111",
    7949=>"011011011",
    7950=>"110010011",
    7951=>"000001001",
    7952=>"000000011",
    7953=>"101101100",
    7954=>"100110010",
    7955=>"100110011",
    7956=>"000010010",
    7957=>"000010110",
    7958=>"111110110",
    7959=>"100100100",
    7960=>"000100100",
    7961=>"000000011",
    7962=>"101100100",
    7963=>"101100110",
    7964=>"000010011",
    7965=>"000011101",
    7966=>"111101110",
    7967=>"110010010",
    7968=>"010010000",
    7969=>"011010001",
    7970=>"111100100",
    7971=>"001000000",
    7972=>"101101100",
    7973=>"010011001",
    7974=>"100100110",
    7975=>"100110010",
    7976=>"010000001",
    7977=>"100000000",
    7978=>"110100110",
    7979=>"100100100",
    7980=>"110111010",
    7981=>"010110010",
    7982=>"011011011",
    7983=>"011111011",
    7984=>"101110110",
    7985=>"000110111",
    7986=>"000000000",
    7987=>"000001011",
    7988=>"001001001",
    7989=>"111011011",
    7990=>"011011011",
    7991=>"100100100",
    7992=>"101100100",
    7993=>"110011111",
    7994=>"001100000",
    7995=>"010010010",
    7996=>"001100100",
    7997=>"000101101",
    7998=>"011011011",
    7999=>"100100010",
    8000=>"100000011",
    8001=>"000000011",
    8002=>"111110000",
    8003=>"000000111",
    8004=>"000001111",
    8005=>"100000110",
    8006=>"101111011",
    8007=>"011000001",
    8008=>"000000010",
    8009=>"111110000",
    8010=>"100000111",
    8011=>"111011000",
    8012=>"111000111",
    8013=>"000101011",
    8014=>"111001100",
    8015=>"001000000",
    8016=>"111101101",
    8017=>"001100111",
    8018=>"000110111",
    8019=>"001100110",
    8020=>"000001000",
    8021=>"000000000",
    8022=>"000101111",
    8023=>"101000010",
    8024=>"110000000",
    8025=>"001110110",
    8026=>"001010011",
    8027=>"101010000",
    8028=>"000000010",
    8029=>"100001000",
    8030=>"001011010",
    8031=>"100111010",
    8032=>"111000000",
    8033=>"011011010",
    8034=>"001010000",
    8035=>"100000000",
    8036=>"001001111",
    8037=>"110011100",
    8038=>"000011010",
    8039=>"000111011",
    8040=>"010011000",
    8041=>"111010000",
    8042=>"001010110",
    8043=>"000000110",
    8044=>"011001100",
    8045=>"101110111",
    8046=>"111111000",
    8047=>"110101100",
    8048=>"001000111",
    8049=>"001000000",
    8050=>"100101001",
    8051=>"001110111",
    8052=>"010000111",
    8053=>"000100001",
    8054=>"110111001",
    8055=>"000000100",
    8056=>"001110010",
    8057=>"010000101",
    8058=>"001001100",
    8059=>"010010111",
    8060=>"000001111",
    8061=>"101000000",
    8062=>"011011001",
    8063=>"110000000",
    8064=>"100101000",
    8065=>"000000010",
    8066=>"000010000",
    8067=>"111100111",
    8068=>"001110100",
    8069=>"001000000",
    8070=>"111000111",
    8071=>"100100000",
    8072=>"011011000",
    8073=>"100000010",
    8074=>"100100001",
    8075=>"001111001",
    8076=>"101101111",
    8077=>"011111010",
    8078=>"011111100",
    8079=>"000010111",
    8080=>"101000000",
    8081=>"111010000",
    8082=>"010101100",
    8083=>"111011101",
    8084=>"111001101",
    8085=>"000100111",
    8086=>"110110111",
    8087=>"110000011",
    8088=>"001001001",
    8089=>"011101000",
    8090=>"110000000",
    8091=>"100001000",
    8092=>"111111000",
    8093=>"011111000",
    8094=>"011100111",
    8095=>"010000100",
    8096=>"111000001",
    8097=>"011010010",
    8098=>"101110111",
    8099=>"010000001",
    8100=>"111001111",
    8101=>"000001000",
    8102=>"110010010",
    8103=>"111101101",
    8104=>"000101000",
    8105=>"000000000",
    8106=>"010001101",
    8107=>"000000100",
    8108=>"000101100",
    8109=>"111100100",
    8110=>"100111101",
    8111=>"101100000",
    8112=>"111110000",
    8113=>"111000000",
    8114=>"011000000",
    8115=>"001000000",
    8116=>"000011010",
    8117=>"000011111",
    8118=>"000000110",
    8119=>"110100100",
    8120=>"110010011",
    8121=>"001100100",
    8122=>"110110000",
    8123=>"110111001",
    8124=>"111000100",
    8125=>"100000000",
    8126=>"110001001",
    8127=>"111000101",
    8128=>"010110111",
    8129=>"100101101",
    8130=>"010000010",
    8131=>"001000101",
    8132=>"010000000",
    8133=>"100001001",
    8134=>"011010110",
    8135=>"001010010",
    8136=>"110011011",
    8137=>"010010010",
    8138=>"011010111",
    8139=>"000010100",
    8140=>"111111111",
    8141=>"110101001",
    8142=>"001010000",
    8143=>"000010010",
    8144=>"001001100",
    8145=>"100101001",
    8146=>"110100111",
    8147=>"011000000",
    8148=>"111010011",
    8149=>"000010010",
    8150=>"100101111",
    8151=>"011010110",
    8152=>"100101001",
    8153=>"101010100",
    8154=>"001001000",
    8155=>"011110110",
    8156=>"000011111",
    8157=>"100101001",
    8158=>"111111111",
    8159=>"011010110",
    8160=>"011010000",
    8161=>"010110110",
    8162=>"110101001",
    8163=>"000000000",
    8164=>"110111100",
    8165=>"100000001",
    8166=>"010110110",
    8167=>"110000000",
    8168=>"001010110",
    8169=>"000000000",
    8170=>"010011001",
    8171=>"000001000",
    8172=>"101011111",
    8173=>"011010100",
    8174=>"110111010",
    8175=>"110110110",
    8176=>"100100100",
    8177=>"000001001",
    8178=>"110100001",
    8179=>"011110111",
    8180=>"010111100",
    8181=>"010111100",
    8182=>"011010110",
    8183=>"100000000",
    8184=>"110001011",
    8185=>"011100110",
    8186=>"011010010",
    8187=>"011010100",
    8188=>"100001001",
    8189=>"100001001",
    8190=>"011010110",
    8191=>"010100110");

BEGIN
    weight <= ROM_content(to_integer(address));
END RTL;