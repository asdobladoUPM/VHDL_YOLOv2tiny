LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L5BNROM IS
    PORT (
        coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); -- Instruction bus
        address : IN unsigned(9 DOWNTO 0));
END L5BNROM;

ARCHITECTURE RTL OF L5BNROM IS

    TYPE ROM_mem IS ARRAY (0 TO 1023) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem :=
    (0=>"1011101101010100"&"0100011101000000",
    1=>"0000011000110000"&"0101001000010001",
    2=>"1111110100111000"&"0101011011110010",
    3=>"1110101100110010"&"0100001100101100",
    4=>"1110010010000001"&"0100100010101011",
    5=>"1101101101111111"&"0100111010110010",
    6=>"1101110101111111"&"0100100111010101",
    7=>"1101000001011100"&"0101001111100010",
    8=>"1101100000010001"&"0101000011001000",
    9=>"1100010010111110"&"0100101000111000",
    10=>"1110000000100100"&"0100010010111001",
    11=>"1111101100001000"&"0100011001111001",
    12=>"1101001000101010"&"0100010100111011",
    13=>"1110001011001110"&"0100101000101111",
    14=>"1110100111001110"&"0100011001000110",
    15=>"1100110101010001"&"0101010111011001",
    16=>"1101100011001101"&"0100101000101000",
    17=>"1101100100101010"&"0100101010101001",
    18=>"1110001000000110"&"0100101111110000",
    19=>"1110000101101010"&"0100100001000110",
    20=>"1011111111000011"&"0101000010010111",
    21=>"1100001011110101"&"0100100010101111",
    22=>"1110101110000110"&"0100101110111011",
    23=>"1011011100000100"&"0011111111000001",
    24=>"1100000110010101"&"0100111110110010",
    25=>"1110110111001100"&"0100101001000010",
    26=>"1101001100010000"&"0100001000010010",
    27=>"1110101110010010"&"0100101010001011",
    28=>"1101110000111100"&"0100010010101101",
    29=>"1111100100110011"&"0100101110100010",
    30=>"1110011100101001"&"0100101100101011",
    31=>"1101101101111110"&"0100001110011110",
    32=>"1100011011100011"&"0101000100001110",
    33=>"1101111110011111"&"0100101111011001",
    34=>"1110100111000111"&"0101011010010110",
    35=>"1100111101100001"&"0101001000101011",
    36=>"1101010101101011"&"0101111100111111",
    37=>"1100111100101101"&"0100110111000000",
    38=>"1101000011100001"&"0100100100000100",
    39=>"0000001011000000"&"0100101111100011",
    40=>"1100100111011011"&"0100110111101100",
    41=>"1110101011000111"&"0100100110001010",
    42=>"1100011001101010"&"0101000100001000",
    43=>"1110101000011100"&"0100010111000100",
    44=>"1011010101000001"&"0101000011110111",
    45=>"1101101001111110"&"0100101111000101",
    46=>"1100110011001010"&"0100101100111001",
    47=>"1011100010100100"&"0100101100000111",
    48=>"1101110011100111"&"0101011111010111",
    49=>"1110110010000000"&"0100000000101011",
    50=>"1110101110010001"&"0101100010000011",
    51=>"1101000011001110"&"0100100111000010",
    52=>"1110111110000110"&"0100010100101111",
    53=>"1100010010010100"&"0100011001100110",
    54=>"1101011011110110"&"0100100000100010",
    55=>"1101111111100001"&"0100100100001100",
    56=>"1110001010100011"&"0110001101111000",
    57=>"1100101011111101"&"0100110011000000",
    58=>"1100000110001001"&"0101010001000110",
    59=>"1100011110010101"&"0101011001111010",
    60=>"1110000011111010"&"0100100111011001",
    61=>"1101011000001100"&"0100101011110110",
    62=>"1100110011111111"&"0100100001110101",
    63=>"1110000100111000"&"0011111101000001",
    64=>"1101001100010111"&"0100100000001100",
    65=>"1101011001010111"&"0011100100001011",
    66=>"1111101001000110"&"0100101001100001",
    67=>"1110101001110101"&"0100010110011100",
    68=>"0000011100001101"&"0100000001110101",
    69=>"1100111100101010"&"0101000000010001",
    70=>"1011010101001001"&"0101100110011000",
    71=>"1101010101001001"&"0100111100111000",
    72=>"1111000101111100"&"0100010010110000",
    73=>"1110000101111100"&"0101000000011111",
    74=>"1110111101100000"&"0100011111101101",
    75=>"1101001011101010"&"0101001000001101",
    76=>"1100110000111001"&"0100010101101001",
    77=>"1011000111100101"&"0101010111110011",
    78=>"1110010111100111"&"0100010111000110",
    79=>"1110010110010001"&"0100011110110110",
    80=>"1101000000011100"&"0101010000010010",
    81=>"1011110111000101"&"0100011111010111",
    82=>"1110100111010111"&"0101010001001110",
    83=>"1110000110010001"&"0101000010110111",
    84=>"1110100010011101"&"0100010110101001",
    85=>"1101101011111011"&"0101101101100000",
    86=>"0000101111010011"&"0100100110011000",
    87=>"1110001100010100"&"0100100110110111",
    88=>"1110111001111111"&"0100101000111000",
    89=>"1101101011010000"&"0100110110000101",
    90=>"1100110101110111"&"0100100111110011",
    91=>"1110010001011001"&"0100000011010100",
    92=>"1101110110101111"&"0100111101010010",
    93=>"1100011001010110"&"0101000100000111",
    94=>"1101111111110100"&"0100110101110110",
    95=>"1100111000111100"&"0101011101010110",
    96=>"1010101110011001"&"0100100111010111",
    97=>"1110100010001100"&"0100001011000110",
    98=>"1101011011101111"&"0100101111011011",
    99=>"1110000100011000"&"0100010011000111",
    100=>"1101100010010111"&"0100000110001011",
    101=>"1110011111100010"&"0101001111010101",
    102=>"0000010010011101"&"0100100011010001",
    103=>"1110100100100011"&"0100000100011001",
    104=>"1101101101100101"&"0100011011001100",
    105=>"1010000010110110"&"0101000010110000",
    106=>"1111000111011000"&"0100100001000011",
    107=>"1110111100010110"&"0100000101110110",
    108=>"1110001000101111"&"0100110000000000",
    109=>"1101110010000001"&"0100100000111011",
    110=>"1100010001111111"&"0100001110111110",
    111=>"1011001101111011"&"0101010101001100",
    112=>"1111001100111010"&"0101111101111000",
    113=>"1111101100011100"&"0100000010010111",
    114=>"1100000000011001"&"0101100010011000",
    115=>"1010110011001100"&"0101101010011111",
    116=>"1101110001101000"&"0100111100101110",
    117=>"1110011011010001"&"0100101001101010",
    118=>"1110111110000001"&"0101011001010100",
    119=>"1110101001110010"&"0100111010101100",
    120=>"1101010100011001"&"0100010011000110",
    121=>"1110010000110110"&"0100100000111100",
    122=>"1111101011101111"&"0100101000100001",
    123=>"1111000000110001"&"0100111000010101",
    124=>"1100011100111110"&"0100010101000011",
    125=>"1101000010010111"&"0101000100110010",
    126=>"1101101101110010"&"0100101100011100",
    127=>"1101001111000010"&"0100100100001001",
    128=>"1101110101101110"&"0100001000110011",
    129=>"1110110001010010"&"0100010101110111",
    130=>"1110011011011110"&"0100010101110001",
    131=>"1011100111101111"&"0101101000000100",
    132=>"1100110101111011"&"0100101010100010",
    133=>"1100011011110010"&"0110000110000100",
    134=>"1101111110001001"&"0100110100111100",
    135=>"1111010011001010"&"0100011100110001",
    136=>"0000000000011001"&"0100101011110110",
    137=>"1110111011010111"&"0100000001011001",
    138=>"1101000100011101"&"0100010110111111",
    139=>"1110001111011010"&"0100101010011111",
    140=>"1011110001101111"&"0100110110100011",
    141=>"1101001101011000"&"0100011001000000",
    142=>"1101101010001100"&"0100010101011111",
    143=>"1111000001000001"&"0100100010011000",
    144=>"1101001010000010"&"0101010100110011",
    145=>"1111111111111010"&"0100001110010101",
    146=>"1101001110101100"&"0100101100011010",
    147=>"1101110111110001"&"0100111011100001",
    148=>"1110110110101111"&"0100110101110001",
    149=>"1110100010100001"&"0100110011011101",
    150=>"1101110100101000"&"0100001100111010",
    151=>"1101011101110010"&"0101001011001110",
    152=>"1110010100010100"&"0101011001100001",
    153=>"1101011010110001"&"0101010100001001",
    154=>"1100010000001101"&"0101011000010100",
    155=>"1110000000010101"&"0100100110001100",
    156=>"1100100100100110"&"0100101010111010",
    157=>"1101110000011010"&"0101000001001100",
    158=>"1101000101110000"&"0100101111101101",
    159=>"1111101000110110"&"0110000000110101",
    160=>"1011111011001111"&"0101011001001010",
    161=>"1110111000000100"&"0100101010010110",
    162=>"1100010000110110"&"0100100101101111",
    163=>"1011000011110111"&"0101101110001110",
    164=>"1111010000110011"&"0100100000011111",
    165=>"1010011000000001"&"0101010111110000",
    166=>"1111001111010110"&"0100101001000010",
    167=>"1100110001011000"&"0100100111010100",
    168=>"1111010000111010"&"0100100100111011",
    169=>"1101001100101110"&"0100111101110100",
    170=>"1101110100000110"&"0100101111100000",
    171=>"1111111011001001"&"0100100101111011",
    172=>"1110100010011100"&"0100010010110100",
    173=>"1010110010000100"&"0101001100000011",
    174=>"1100011001101001"&"0100110000010011",
    175=>"1110110010101011"&"0100101000000011",
    176=>"1110000101010010"&"0100110001010011",
    177=>"1011101110100101"&"0100110111110110",
    178=>"1110100110000000"&"0100110000100111",
    179=>"1110001110101100"&"0100001011010000",
    180=>"0000010001110010"&"0100100011011001",
    181=>"1110001011000111"&"0100011111100110",
    182=>"1110111110011100"&"0011111110110000",
    183=>"1111100000011111"&"0100010011000001",
    184=>"1111011001110110"&"0100000010111101",
    185=>"1111100111010101"&"0101000101100001",
    186=>"1101000101011000"&"0100000111010010",
    187=>"1100000001000001"&"0100110101011000",
    188=>"1110111000100100"&"0101101001100011",
    189=>"1100111110000010"&"0100011011101101",
    190=>"1110001011010001"&"0101000100000011",
    191=>"1101111011001101"&"0100011111011000",
    192=>"1011011110000100"&"0101010111100110",
    193=>"1111101101101100"&"0100100001011101",
    194=>"1100111110011111"&"0100010100101011",
    195=>"1011111000000011"&"0100111111001110",
    196=>"1101110001011011"&"0100110011101110",
    197=>"1101100100101000"&"0101011001010000",
    198=>"1101010001001100"&"0101001100001001",
    199=>"1100100010110110"&"0101101000110011",
    200=>"1101101100011011"&"0100001111000011",
    201=>"1110010001001000"&"0101111001001100",
    202=>"1011110110000001"&"0100101011011111",
    203=>"1100011000000001"&"0101000110010100",
    204=>"1101000110110001"&"0100111101101111",
    205=>"1111001011011001"&"0101101001100010",
    206=>"1110010011000111"&"0100010111110011",
    207=>"1100011101000101"&"0100011101011011",
    208=>"1101101000000011"&"0101011000110000",
    209=>"1110000111010011"&"0100111111101101",
    210=>"1101000110110001"&"0100110010100001",
    211=>"1111001011011010"&"0101000101001001",
    212=>"1100101111000011"&"0100101001011010",
    213=>"1101111001010011"&"0100100000111100",
    214=>"1101100110001101"&"0100101101100010",
    215=>"1101001011110010"&"0101001000110010",
    216=>"1101100111101001"&"0100100010111001",
    217=>"1110101101001100"&"0100110011110100",
    218=>"1100011011001001"&"0100000010111000",
    219=>"1101011101000010"&"0100001001001100",
    220=>"1101000111011000"&"0100001010000011",
    221=>"1011100000000000"&"0101010001011100",
    222=>"1011101000110100"&"0101111001001001",
    223=>"1101011101100011"&"0101011011011110",
    224=>"1011101010011000"&"0101010101010111",
    225=>"1101010000010010"&"0100101010100000",
    226=>"1101001110010101"&"0100110011010000",
    227=>"1010110110001101"&"0100100110010010",
    228=>"1110011011111111"&"0100111001001111",
    229=>"1110101011001100"&"0100000001011100",
    230=>"1111001110000110"&"0010011001111100",
    231=>"1111110111110001"&"0101010010110111",
    232=>"1110000100000011"&"0101000110011011",
    233=>"1101010010010101"&"0100111110010011",
    234=>"1110000100011111"&"0100100110111110",
    235=>"1100110101100010"&"0101011000010111",
    236=>"0000011111110101"&"0100111000111110",
    237=>"1101010101001000"&"0100100001111011",
    238=>"1011110011111000"&"0100100111000101",
    239=>"1100110100100111"&"0100110001010011",
    240=>"1110101101111000"&"0100011110000111",
    241=>"1101100001110001"&"0100100101011001",
    242=>"1110100111000001"&"0101010010111010",
    243=>"1100101111110110"&"0100100110111111",
    244=>"1110111010111000"&"0101000010000001",
    245=>"1101111111111000"&"0101111000000100",
    246=>"1111100010000011"&"0100010100000001",
    247=>"1110010010000001"&"0100100001111001",
    248=>"1101110010111110"&"0100001110001011",
    249=>"1110000010100001"&"0100001001100111",
    250=>"1110011110010010"&"0100100111000101",
    251=>"1110011111010010"&"0011101011100111",
    252=>"1110010001001101"&"0100001000011111",
    253=>"1110011110110011"&"0100011111010110",
    254=>"1100101110001110"&"0101010000100110",
    255=>"1011110011000101"&"0101010000000111",
    256=>"1110001101101110"&"0101100001110000",
    257=>"1110100101110100"&"0100101111000111",
    258=>"1110011111000101"&"0100110000000111",
    259=>"1110011010001001"&"0101100000010001",
    260=>"1111100101001110"&"0100011001001101",
    261=>"1110001010111011"&"0100111101100100",
    262=>"1110111000010101"&"0100111111110101",
    263=>"1110011101000000"&"0100011000111111",
    264=>"1111010001111101"&"0100011100101111",
    265=>"1101101111111001"&"0100110010001000",
    266=>"1101110101100110"&"0101100101111101",
    267=>"1101010001110111"&"0100110000110010",
    268=>"1110011101011011"&"0100011101001000",
    269=>"1101110101100101"&"0100100011100100",
    270=>"1110100010100010"&"0100110100100011",
    271=>"1100101010101110"&"0100100101110000",
    272=>"1110011000111000"&"0100101101101101",
    273=>"1110111101100100"&"0100001111111110",
    274=>"1100111110011100"&"0101000111100000",
    275=>"1100101101001110"&"0100111110111101",
    276=>"1110010011100100"&"0100110010010100",
    277=>"1110001100000111"&"0100010010111011",
    278=>"1111100101110010"&"0100010000111110",
    279=>"1100101111111111"&"0101001000110100",
    280=>"1100010111111011"&"0100110111001101",
    281=>"1100011111101111"&"0101011001010100",
    282=>"1101110101100000"&"0100010111001110",
    283=>"1101010110011101"&"0100110000011101",
    284=>"1110111111111010"&"0100011000100010",
    285=>"1101000110011111"&"0101001010100000",
    286=>"1111001100100011"&"0100100100111011",
    287=>"1110100011111101"&"0100101001100010",
    288=>"1100000010011111"&"0101011100001011",
    289=>"1101110011100000"&"0100011001001101",
    290=>"1101100001001000"&"0100111111001010",
    291=>"1111011011100011"&"0100100111000110",
    292=>"1110000101010101"&"0100011110010100",
    293=>"1111101001100110"&"0100011111101101",
    294=>"0001000011001111"&"0100001110110110",
    295=>"1110011100011011"&"0100101011011111",
    296=>"1101010111101110"&"0101010011101011",
    297=>"1101100010001110"&"0100110100101111",
    298=>"1110110101110001"&"0100011011111110",
    299=>"1110001010000111"&"0100000011101000",
    300=>"1110101111001101"&"0100110001010011",
    301=>"1110011001010011"&"0100110011111011",
    302=>"1100110010000011"&"0100101110110111",
    303=>"0000000110001101"&"0100101110110110",
    304=>"1111110100011011"&"0100101001011011",
    305=>"1100110110001101"&"0100110000110100",
    306=>"1101101000001110"&"0100010101110000",
    307=>"1101101001010101"&"0100111010101011",
    308=>"1110010100101100"&"0100010111001011",
    309=>"1101101001000101"&"0101000111100100",
    310=>"1110110000010010"&"0101000101000011",
    311=>"1101000111011110"&"0100011110110010",
    312=>"1101000100101010"&"0100001010001000",
    313=>"1110100110001111"&"0100110110001000",
    314=>"1110111011001110"&"0100010011101100",
    315=>"1111110111110100"&"0101001010011000",
    316=>"1110101111101100"&"0100100011100010",
    317=>"1110101110001010"&"0101001010101110",
    318=>"1110100100110101"&"0100101000000001",
    319=>"1110111111110011"&"0100011011001111",
    320=>"1111010110110111"&"0100001111000110",
    321=>"1100111110001001"&"0100111101001001",
    322=>"1111100011110000"&"0100101111001100",
    323=>"1100101001111011"&"0100001011011010",
    324=>"1111010011011110"&"0100001000110011",
    325=>"1101101100111011"&"0101011000101000",
    326=>"1101001000001010"&"0100111001111110",
    327=>"1110101100000010"&"0100110011001100",
    328=>"1101111100001101"&"0101000011101100",
    329=>"1100011111011100"&"0011111100011100",
    330=>"1110100110101010"&"0100011100010110",
    331=>"1100110110100011"&"0100010110001101",
    332=>"1101100111001011"&"0101001000001110",
    333=>"1100100000010101"&"0101111011010000",
    334=>"1110001010011011"&"0011111111110101",
    335=>"1100110100001001"&"0011111101001101",
    336=>"1101000111010100"&"0100100001000001",
    337=>"1100011111100011"&"0101110101000001",
    338=>"1110101011100011"&"0100101010101001",
    339=>"1111111110011100"&"0100101100100110",
    340=>"1110001111000111"&"0101100101011100",
    341=>"1101101111000000"&"0100000001111110",
    342=>"1100111101001000"&"0100110010101101",
    343=>"1110010011011101"&"0100110100101110",
    344=>"1111010101010001"&"0100100111001000",
    345=>"1101000111110000"&"0100000010010011",
    346=>"1101000100001011"&"0100010100101111",
    347=>"1110000011100000"&"0100100111001100",
    348=>"1101000000011101"&"0100010100000100",
    349=>"1110010000010011"&"0101010100010110",
    350=>"1101101100110010"&"0100111000000110",
    351=>"1110010111011000"&"0101000111000010",
    352=>"1110001101100000"&"0100001011011000",
    353=>"0000001000010011"&"0100110000010010",
    354=>"1101110100010110"&"0101011001001110",
    355=>"1101001111110100"&"0100110011101111",
    356=>"1110111001001000"&"0101001101000100",
    357=>"1110010001111011"&"0100111101000110",
    358=>"1101111000100111"&"0101010101101110",
    359=>"1101011011011000"&"0100100110001101",
    360=>"1111010001110100"&"0100011100110001",
    361=>"1101011010111011"&"0100100000011100",
    362=>"1110111000011110"&"0100101001110110",
    363=>"1101101101010010"&"0101011011110101",
    364=>"1101100001100100"&"0100010110011110",
    365=>"1100010001010010"&"0110000011111111",
    366=>"1100010001101101"&"0101000101101000",
    367=>"1110011001111101"&"0100111100111110",
    368=>"1101101000110111"&"0100101011110001",
    369=>"1100010111110110"&"0101010010100000",
    370=>"1110010001100110"&"0101000010100100",
    371=>"0000000100011110"&"0100011100000110",
    372=>"1101011001010010"&"0101111000110000",
    373=>"1100001110110011"&"0100011011011111",
    374=>"1011111110100111"&"0100111010011101",
    375=>"1110011000110101"&"0100101101001111",
    376=>"1110011010001111"&"0100111011001010",
    377=>"1100110110011111"&"0100010100110100",
    378=>"1110100011100101"&"0101010001100011",
    379=>"1101011111001110"&"0100110011111001",
    380=>"1100111110011011"&"0100010011000000",
    381=>"1111000010100111"&"0100111010010111",
    382=>"1111000001000100"&"0101101010110000",
    383=>"1100100101011010"&"0100010110000110",
    384=>"1111110000000101"&"0100100010001100",
    385=>"1111101010100010"&"0011110010111110",
    386=>"0001000011011001"&"0100111010110000",
    387=>"1101111100001011"&"0011011010010001",
    388=>"1110101110100110"&"0101010011000010",
    389=>"1100110011100010"&"0100111011111011",
    390=>"1100100111110001"&"0101100100100011",
    391=>"1111100010111000"&"0100010100110011",
    392=>"1010101101111011"&"0101011001010110",
    393=>"1011100000010011"&"0100101101110001",
    394=>"1110111011110011"&"0011111111011110",
    395=>"1101000110011101"&"0100100110110111",
    396=>"1110111011111001"&"0100001010011010",
    397=>"1100001000100001"&"0101011011110000",
    398=>"1110000111111011"&"0100100111011001",
    399=>"1110001101110010"&"0101000011101101",
    400=>"1101101010010110"&"0100100010001010",
    401=>"1101000101011110"&"0100101000100010",
    402=>"1100010001001000"&"0100010011110110",
    403=>"1110010001010010"&"0100110010000001",
    404=>"1101011100101000"&"0100101001110001",
    405=>"1100010010101100"&"0100101010000011",
    406=>"0000001011111001"&"0100011000110101",
    407=>"1101000011010001"&"0100101110101101",
    408=>"1011011110000101"&"0100110000011000",
    409=>"1100110011111010"&"0101011101011101",
    410=>"0000000000100101"&"0100100011110110",
    411=>"1100000010100101"&"0100101110010000",
    412=>"1111100100110011"&"0100111010001100",
    413=>"1101111000110101"&"0100011011110000",
    414=>"1101100001000111"&"0101000100100110",
    415=>"1110100000010100"&"0101110110101011",
    416=>"1100101111111110"&"0100011010101100",
    417=>"1101000001110011"&"0101010110010101",
    418=>"1110101001011010"&"0100001111110111",
    419=>"1101101101010001"&"0100010110101000",
    420=>"1010110000100100"&"0100110111011110",
    421=>"1111001011111110"&"0011111011010100",
    422=>"1011011001010101"&"0101001011001011",
    423=>"1100111000100101"&"0100110011010101",
    424=>"1111000111111000"&"0101000001111001",
    425=>"1111010010001111"&"0100001010111101",
    426=>"1111100011001101"&"0100000001100001",
    427=>"1101011111111110"&"0100101100000001",
    428=>"1011101100100010"&"0100111100100111",
    429=>"1101100110110001"&"0100110001100101",
    430=>"1110110110001001"&"0100111001001110",
    431=>"1101110000000110"&"0100010011100001",
    432=>"1110100110010100"&"0100010011100010",
    433=>"1110111010010101"&"0100010001110101",
    434=>"1100000111100011"&"0100011011001100",
    435=>"1110110100001011"&"0100011100011110",
    436=>"1100011100111111"&"0100110100111001",
    437=>"0000000110100001"&"0100010101010011",
    438=>"1110101100100001"&"0100011111111110",
    439=>"1101101011001100"&"0100011011001011",
    440=>"1101111101100111"&"0100101111101000",
    441=>"1101100011001010"&"0100100100111111",
    442=>"1101110010000011"&"0100101100101010",
    443=>"1101011010000001"&"0101100101110000",
    444=>"1111100001110110"&"0101011000001001",
    445=>"1101111111011100"&"0100110100001100",
    446=>"1110001000010100"&"0100011011010001",
    447=>"1101001011000110"&"0101001000110110",
    448=>"1100111101110010"&"0101001101011111",
    449=>"1101111010000000"&"0100100111100001",
    450=>"1111000111011001"&"0100010000000011",
    451=>"1110010100110110"&"0101001010101001",
    452=>"1110100110010101"&"0100100111010000",
    453=>"1100010100010011"&"0100111010001110",
    454=>"1110101101011001"&"0101000111011110",
    455=>"1011101000100001"&"0100010111101100",
    456=>"1110001101010100"&"0101010100010110",
    457=>"1110000010101000"&"0100110001111110",
    458=>"1110111011110111"&"0100100101100100",
    459=>"1111000100100011"&"0100100000011100",
    460=>"1011101011010111"&"0100011011111111",
    461=>"1100100000000000"&"0101001001001001",
    462=>"1101100111100011"&"0100111100000101",
    463=>"1101010111011100"&"0100010100001000",
    464=>"1110010001100011"&"0100100010010101",
    465=>"1111110011010110"&"0001111000100011",
    466=>"1101111011010001"&"0100110100000100",
    467=>"1101001010011101"&"0100111000101111",
    468=>"1101011011100001"&"0100010110110110",
    469=>"1101011111000110"&"0101011110111101",
    470=>"1101001011010111"&"0100000001000010",
    471=>"1101110010010110"&"0100011111010001",
    472=>"1101001110001000"&"0100110110000011",
    473=>"1100100001101111"&"0100111100110101",
    474=>"1101111101110010"&"0100100011010000",
    475=>"1100100101100011"&"0101011011111001",
    476=>"1110101100001111"&"0100010101011101",
    477=>"1110011100010100"&"0100101000001101",
    478=>"1110010110101001"&"0100011110101110",
    479=>"1101100011101110"&"0101101000111000",
    480=>"1110011100011110"&"0101010111100110",
    481=>"1111011001011010"&"0100001110010000",
    482=>"1111111111110110"&"0100001001110110",
    483=>"1111000101100010"&"0101100011100111",
    484=>"1110100100101110"&"0100100110100111",
    485=>"1111101100110110"&"0100101001010101",
    486=>"1100011100111001"&"0100101011001010",
    487=>"1100111001000101"&"0101011010101000",
    488=>"1111000011101011"&"0100001011111001",
    489=>"1110111001011110"&"0110010101110001",
    490=>"1100111001000001"&"0100010010001100",
    491=>"1101111111100011"&"0101011111101000",
    492=>"1111110110011111"&"0100110101111111",
    493=>"1100000110010100"&"0101000000110101",
    494=>"1101011000110100"&"0100100011100001",
    495=>"1100011001001101"&"0100100010100111",
    496=>"1111000001011010"&"0100100001010010",
    497=>"1100000010000110"&"0101110001000111",
    498=>"1100111001101111"&"0100011111110001",
    499=>"1101000111101101"&"0100010011110100",
    500=>"1110111100111111"&"0100011110001010",
    501=>"1110010000011101"&"0101100011110010",
    502=>"1101101000100100"&"0100110101111101",
    503=>"1101111111100100"&"0101101010011101",
    504=>"1011100101110010"&"0101000110111100",
    505=>"1110010011101111"&"0100101111100100",
    506=>"1110010011111110"&"0100110010000010",
    507=>"1111100101000010"&"0100011101011001",
    508=>"1101000101101111"&"0100011101101101",
    509=>"1100101011101100"&"0100111100001000",
    510=>"1101100111010000"&"0101101101111110",
    511=>"1110011001010001"&"0100101100001011",
    512=>"1100110011011101"&"0101100111011100",
    513=>"1101110101000110"&"0100011010111010",
    514=>"1110001110001100"&"0100010100010110",
    515=>"1111001100010110"&"0011011010100010",
    516=>"1100101000000100"&"0100100010100111",
    517=>"1101110011111001"&"0100011010100100",
    518=>"1101101100000001"&"0101000010001010",
    519=>"1101110110001100"&"0100000111001011",
    520=>"1011100111010101"&"0100011001011111",
    521=>"1101010000111001"&"0100010101010000",
    522=>"1110100000111100"&"0101000010100001",
    523=>"1101101000001000"&"0100101011011111",
    524=>"1101010011010011"&"0100111100101110",
    525=>"1110110011000011"&"0100110101010101",
    526=>"1111110001001001"&"0100011001100111",
    527=>"1101111010100100"&"0100110001100001",
    528=>"1111000111000111"&"0100101011010010",
    529=>"1110001001000100"&"0100100001100010",
    530=>"1101100010110110"&"0100110110100111",
    531=>"1101111101001110"&"0100111100110111",
    532=>"1101001101000010"&"0011101101101010",
    533=>"1111010001010000"&"0100100001000010",
    534=>"1110010011010011"&"0110001110001110",
    535=>"1101001011101101"&"0100111111000001",
    536=>"1110010111100010"&"0100110010100111",
    537=>"1110010000100110"&"0100101011011110",
    538=>"1110001001000011"&"0100000110110011",
    539=>"1110001000001101"&"0100101010101000",
    540=>"1110110111100011"&"0101000110000011",
    541=>"1100011010001000"&"0100111000101101",
    542=>"1101110001011111"&"0100110101100101",
    543=>"1111010011000000"&"0100010001110110",
    544=>"1111001011101011"&"0100000100011001",
    545=>"1101000000100110"&"0100110010001111",
    546=>"1011010010100011"&"0100110111011001",
    547=>"1011111110001111"&"0100010101010001",
    548=>"1110101001010011"&"0100001110100000",
    549=>"1101110101101101"&"0100101010010111",
    550=>"1101011101011101"&"0100110110001010",
    551=>"1110111011000100"&"0101000011101100",
    552=>"1100101101000011"&"0011101111000011",
    553=>"1111000001011100"&"0100010110100100",
    554=>"1100111010100001"&"0101011001011101",
    555=>"1110001001100110"&"0100101100100011",
    556=>"1110001011010111"&"0100010011110001",
    557=>"1110000000011100"&"0100100010000000",
    558=>"1110110101100110"&"0101011000110001",
    559=>"1110000001100111"&"0100011100110010",
    560=>"1101111010011111"&"0100111011000010",
    561=>"1101110111101101"&"0100000000011100",
    562=>"1101000101111101"&"0110001011101100",
    563=>"1101001100010000"&"0100110111011011",
    564=>"1100111101010010"&"0100100011001001",
    565=>"1111010001001000"&"0100101000000000",
    566=>"1101001011000111"&"0100011101001110",
    567=>"1111010100011100"&"0101010010101101",
    568=>"1110001000001111"&"0100100101001011",
    569=>"1100010101100010"&"0100101111010111",
    570=>"1101101110001110"&"0101010110001111",
    571=>"1110010100110011"&"0100100111001011",
    572=>"1110111010000100"&"0101001101100110",
    573=>"1110001010101001"&"0100001100010000",
    574=>"1110010101110111"&"0100001110001000",
    575=>"1100011000100000"&"0100110001000100",
    576=>"1011100111010100"&"0101010100100001",
    577=>"1110000111010000"&"0100100100011001",
    578=>"1101000110111100"&"0101010010011100",
    579=>"1101011010100100"&"0101101100010111",
    580=>"1110011100011110"&"0100010001010000",
    581=>"1101110010001001"&"0100101111011110",
    582=>"1111000111011011"&"0100011000001111",
    583=>"1111101110001111"&"0101001000111111",
    584=>"1111010010100011"&"0100110100111101",
    585=>"1111000101001100"&"0101100101011000",
    586=>"1110000001001101"&"0101000101011001",
    587=>"1111000101001000"&"0100000000100111",
    588=>"1011010001101110"&"0101011001100100",
    589=>"1101000111000001"&"0100001001000001",
    590=>"1101110011100001"&"0100111110101100",
    591=>"1101000010011100"&"0101001011011000",
    592=>"1111110010110111"&"0100111101011000",
    593=>"1101110010110011"&"0100100100011100",
    594=>"1110011101110010"&"0100110010010011",
    595=>"1101010011011101"&"0100010111111001",
    596=>"1110011001000011"&"0101001000011101",
    597=>"1011011111110001"&"0100100100010011",
    598=>"1100000000101000"&"0100000100000101",
    599=>"1110110110011111"&"0100111111111111",
    600=>"1101011000010100"&"0101101011001000",
    601=>"1110011000000001"&"0101011010001111",
    602=>"1110111100010101"&"0100010001101101",
    603=>"1110011010111000"&"0100011010000011",
    604=>"1100110010100110"&"0100101110111010",
    605=>"1110101101101101"&"0100000110010001",
    606=>"1011011101001110"&"0101011101010111",
    607=>"1101110100000010"&"0101111110100110",
    608=>"1110000101110001"&"0100101101101000",
    609=>"1101110001010111"&"0011101100010111",
    610=>"1110110110110110"&"0100011111011111",
    611=>"1101111101000011"&"0100110010001000",
    612=>"1110010100100100"&"0100100010011011",
    613=>"1101011101001010"&"0101000110000011",
    614=>"0000011111011111"&"0101101110110110",
    615=>"1110010111100001"&"0100111011101010",
    616=>"1100000011011011"&"0100010011001100",
    617=>"1110100011000100"&"0101100010110000",
    618=>"1110111010000001"&"0100111111010100",
    619=>"1101010001010101"&"0100010010001100",
    620=>"1111000000010100"&"0100100011001100",
    621=>"1101010011010100"&"0101001101110000",
    622=>"1011100100001110"&"0101100010000101",
    623=>"1110000010010100"&"0101101011001011",
    624=>"1110000001110101"&"0100010011001111",
    625=>"1110011010100100"&"0011111101011001",
    626=>"1110010000100011"&"0100111011110011",
    627=>"1110010100011000"&"0100010100001010",
    628=>"1101110110011100"&"0100101000100110",
    629=>"1111000001111010"&"0100001110100011",
    630=>"1101111010010101"&"0100111000101111",
    631=>"1100101010011100"&"0101001000111100",
    632=>"1101010100110011"&"0100000100101000",
    633=>"1110010000101010"&"0101000000101001",
    634=>"1110000111000100"&"0100101001000110",
    635=>"1110110000011011"&"0100100001000001",
    636=>"1100000001111111"&"0100100111000111",
    637=>"1111000110101100"&"0100100111000010",
    638=>"1101110110110000"&"0011111100100110",
    639=>"1110101100101011"&"0100011010011110",
    640=>"1111110110101100"&"0100010101110111",
    641=>"1100111000011111"&"0100100110001011",
    642=>"1101110111010000"&"0101001000010100",
    643=>"1011100100001001"&"0101101000001100",
    644=>"1101101011101110"&"0101111011110000",
    645=>"1100111010011110"&"0100001010111010",
    646=>"1110010000001110"&"0100101100011100",
    647=>"0000000111001111"&"0101000000100101",
    648=>"1101110001001011"&"0100100010001111",
    649=>"1100100101100110"&"0101100101101111",
    650=>"1110000010010100"&"0101000101111100",
    651=>"1111000111001101"&"0100110110001110",
    652=>"1110011010001101"&"0100101000001101",
    653=>"1110011000100000"&"0100011100001000",
    654=>"1101111100110001"&"0100011010011001",
    655=>"0000010000010100"&"0100100100111001",
    656=>"1110011111001010"&"0101111000110001",
    657=>"1110000010100111"&"0100111001011001",
    658=>"1110101111100011"&"0100001000100010",
    659=>"1111001110001000"&"0100010011011101",
    660=>"1101010010001010"&"0101111101011011",
    661=>"1111100010011100"&"0100100000011001",
    662=>"1111001010110000"&"0101011000011100",
    663=>"1100101000001111"&"0100001011010010",
    664=>"1101011010001110"&"0100101011110000",
    665=>"1111101011101010"&"0100110011101010",
    666=>"1101000000101110"&"0100100011001111",
    667=>"1111011011111010"&"0100011011101011",
    668=>"1110101001100100"&"0100001011000100",
    669=>"1011101101110101"&"0100110101001111",
    670=>"1110101000101101"&"0100111000110111",
    671=>"1111000001010010"&"0100000001010111",
    672=>"1110010101010101"&"0100000110111001",
    673=>"1110011000001000"&"0100111110101100",
    674=>"1110101101001010"&"0101001111011100",
    675=>"1101111110110000"&"0101000100111101",
    676=>"1110000001011000"&"0100001001101010",
    677=>"1101111011011111"&"0101001111000000",
    678=>"1110001000111011"&"0101000111011011",
    679=>"1101010000010111"&"0100101111011100",
    680=>"1101000110110111"&"0101001110010000",
    681=>"1111101001110101"&"0011110110110001",
    682=>"1101011111000001"&"0100011100111111",
    683=>"1011110000000101"&"0101000001111100",
    684=>"1111000100101000"&"0100101011010110",
    685=>"1110011000100100"&"0100011000011110",
    686=>"1110010100000110"&"0100101010110011",
    687=>"1100111000111010"&"0101000111101011",
    688=>"1100100100011001"&"0100110000100100",
    689=>"1111011101111100"&"0101010100000110",
    690=>"1111000001001111"&"0100001011101101",
    691=>"1110100101110010"&"0011101110111101",
    692=>"1011111001010100"&"0100100100110101",
    693=>"1110101111111010"&"0100011111010011",
    694=>"1110110000010111"&"0100101110110010",
    695=>"1110100001101000"&"0100110000110110",
    696=>"1101011101101101"&"0100001100110101",
    697=>"1110101110110101"&"0101010110101110",
    698=>"0000001110000001"&"0100011011110011",
    699=>"1101101111111110"&"0100110010101011",
    700=>"1101110010010111"&"0100010001011001",
    701=>"1111000010101100"&"0011001101111100",
    702=>"1111000011011011"&"0101001010111011",
    703=>"1110001111011110"&"0100110010110011",
    704=>"1101001010100010"&"0100010000100001",
    705=>"1100000110111011"&"0101010001101000",
    706=>"1111000101010111"&"0100110101101100",
    707=>"1110110110001110"&"0101000110100100",
    708=>"1110010111101011"&"0100110110001010",
    709=>"1111000110010010"&"0101001010101110",
    710=>"1101100101110000"&"0100010000110010",
    711=>"1111010000011000"&"0100100010110000",
    712=>"1110110100100111"&"0100110011110110",
    713=>"1110111101001010"&"0100011100100111",
    714=>"1111000110000010"&"0100011000001100",
    715=>"1100000010001001"&"0100111011011101",
    716=>"1110000111110111"&"0100101110100110",
    717=>"1100011000010101"&"0100111000111100",
    718=>"1101101111000101"&"0100101101101010",
    719=>"1101100110010010"&"0100010111111010",
    720=>"1101011101110111"&"0100101011101000",
    721=>"1101011101011000"&"0100101010011111",
    722=>"1101000101100001"&"0100111111011101",
    723=>"1111010101100001"&"0100101101110100",
    724=>"1100110101001100"&"0100100100110000",
    725=>"1111010101001011"&"0100000110001001",
    726=>"0000000000101001"&"0101000101010010",
    727=>"1110101001010110"&"0100011011001011",
    728=>"1101011000000010"&"0101000111010011",
    729=>"1101111011001010"&"0100001011111101",
    730=>"1101100111101011"&"0100111011010000",
    731=>"1101100010010010"&"0100110011010101",
    732=>"1100001111010100"&"0101111111101010",
    733=>"1011011100111001"&"0100011111001111",
    734=>"1111001110010010"&"0100110101100101",
    735=>"1101111000110100"&"0100100110000011",
    736=>"1110100010110100"&"0100010100000011",
    737=>"1101000111111011"&"0011110111101000",
    738=>"1101101010111111"&"0100111111111110",
    739=>"1101110011101010"&"0100111101111111",
    740=>"1110101010111011"&"0100100101101001",
    741=>"1100111010000100"&"0101001000111011",
    742=>"1110101000101100"&"0100101011111110",
    743=>"1100110111010111"&"0100101101011001",
    744=>"1101000010011111"&"0100001111100000",
    745=>"1101110101101011"&"0100011111011001",
    746=>"1100101101010100"&"0100110100010001",
    747=>"1101101111101001"&"0100101100101111",
    748=>"1011001011001100"&"0100110111100000",
    749=>"1111001000101000"&"0100101111001000",
    750=>"1111000110001110"&"0100010101011000",
    751=>"1101111111110101"&"0101101101000100",
    752=>"1101101100011110"&"0100110101111010",
    753=>"1101011110000100"&"0100101001110001",
    754=>"1100110110100101"&"0101000000111100",
    755=>"1110000011111011"&"0101000011010010",
    756=>"1110110001101111"&"0101000011110000",
    757=>"1110000000011110"&"0100101111011010",
    758=>"0000110110111011"&"0101110110010000",
    759=>"1110000111000110"&"0100011011000010",
    760=>"1100110100110011"&"0100100000110100",
    761=>"1110001110101100"&"0101110010001101",
    762=>"1011100101011101"&"0101001100101010",
    763=>"1011000100001000"&"0100101110010110",
    764=>"1101010111001001"&"0100100011101001",
    765=>"1110000110100111"&"0100110011000100",
    766=>"1110001111000001"&"0100011010100011",
    767=>"1101001011100001"&"0100111000101011",
    768=>"1110111111001000"&"0100001010100100",
    769=>"1100010100011010"&"0101001101010011",
    770=>"1101100011111010"&"0101000110110000",
    771=>"1011010000001111"&"0101010100010101",
    772=>"1110001111011001"&"0100100110111101",
    773=>"1110011010001111"&"0100000110101011",
    774=>"1101110100000111"&"0101001110111000",
    775=>"1100010011001100"&"0101001110011101",
    776=>"1101011011001001"&"0100100000001011",
    777=>"1101101001110010"&"0101010100100010",
    778=>"1111100000111001"&"0101000000000001",
    779=>"1100111101111000"&"0100110010100110",
    780=>"1101001101111011"&"0100011000001010",
    781=>"1101010101111101"&"0101010010010011",
    782=>"1111010000011001"&"0100010110110110",
    783=>"1110111001101110"&"0100011010111100",
    784=>"1101011011100011"&"0101111011110101",
    785=>"1100110011011010"&"0011111101011110",
    786=>"1110110111011100"&"0100011011100000",
    787=>"1111100101001000"&"0101100001010011",
    788=>"0000000011101001"&"0100100101011110",
    789=>"1110110000110110"&"0100110110000101",
    790=>"1101001010111011"&"0011111110101000",
    791=>"1101010110000101"&"0100011011111001",
    792=>"1101101100111100"&"0100110010100100",
    793=>"1100111110001001"&"0100101001111010",
    794=>"1100110001111010"&"0101100100001101",
    795=>"1100110001000110"&"0101011010100101",
    796=>"1101111010111001"&"0100100001110100",
    797=>"1110110011001011"&"0100010010101111",
    798=>"1111001101110110"&"0010111001001100",
    799=>"1111101100010111"&"0100101011100100",
    800=>"1110001010010001"&"0100011010010110",
    801=>"1110100011010110"&"0101011001001100",
    802=>"1011011100110101"&"0101011000101000",
    803=>"1100001001110110"&"0100111101100000",
    804=>"1101110111011011"&"0100111011010100",
    805=>"1011000101101000"&"0100111101101110",
    806=>"1100001110011111"&"0110000110011110",
    807=>"1110000100111001"&"0101010101100100",
    808=>"1111100011000001"&"0100100001000111",
    809=>"1101000010110111"&"0101101000111010",
    810=>"1111110010100100"&"0100111000010101",
    811=>"1100101101011111"&"0100100110111001",
    812=>"1011110100001110"&"0101001000010111",
    813=>"1100101101011010"&"0100011111100011",
    814=>"1011111011110100"&"0011110111100111",
    815=>"1100101011010011"&"0100110011010101",
    816=>"1110001010000110"&"0100010100000110",
    817=>"1100101101100011"&"0101110001100000",
    818=>"1100111001111011"&"0100111000010010",
    819=>"1110100101111100"&"0100001100100000",
    820=>"1110000110110010"&"0100110101001001",
    821=>"1101010111011100"&"0100110011001011",
    822=>"1110011001010011"&"0100011001110010",
    823=>"1110011110011001"&"0100100111000111",
    824=>"1110011010101010"&"0100111000011101",
    825=>"1110110110111111"&"0100100010000110",
    826=>"1100101011100011"&"0110001111010111",
    827=>"1110111111010100"&"0100011111101101",
    828=>"1101111011011101"&"0101000100110111",
    829=>"1101100101101010"&"0100101101011011",
    830=>"1110111011001101"&"0100011011111010",
    831=>"1111001000001011"&"0101011011110101",
    832=>"1110110111111000"&"0100010001100110",
    833=>"1100100111101011"&"0101011001100000",
    834=>"1100111001001110"&"0100101110000000",
    835=>"1110001010101110"&"0011111110101010",
    836=>"1101000100110100"&"0101000101010001",
    837=>"0000011000011100"&"0100101001111101",
    838=>"1100001011001011"&"0100011101100001",
    839=>"1110010111010010"&"0100110000110001",
    840=>"1110011001000011"&"0100001100101101",
    841=>"1101110001000110"&"0100111001101001",
    842=>"1110000111101001"&"0100101000111100",
    843=>"1110100011110000"&"0100101101010101",
    844=>"1100111001001010"&"0100110110111000",
    845=>"0000001000111001"&"0100001011101000",
    846=>"1101101001100110"&"0100000100111010",
    847=>"1101010000001111"&"0100111101001011",
    848=>"1100110101001001"&"0100111100000011",
    849=>"1100100101100100"&"0100101001001111",
    850=>"1110010100011010"&"0100111111100101",
    851=>"1110100010101101"&"0011111110000101",
    852=>"1111001011010111"&"0100011010011111",
    853=>"1110100001101010"&"0100100100001110",
    854=>"1100000110001011"&"0101100001101100",
    855=>"1110011111001001"&"0101000010001101",
    856=>"1101110001100010"&"0100101001100010",
    857=>"1101101110100100"&"0101011111100101",
    858=>"1111011010000010"&"0100010000001100",
    859=>"1100011101010000"&"0101101000011110",
    860=>"1100100001100101"&"0100111001011101",
    861=>"1100010011000100"&"0101010101011001",
    862=>"1101010000111001"&"0100010111010000",
    863=>"1011010101110100"&"0100010101110001",
    864=>"1111011011101100"&"0100011001000001",
    865=>"1101110101100000"&"0100100101110111",
    866=>"1101001011110001"&"0100011100001010",
    867=>"1110000010010011"&"0100101011011011",
    868=>"1110110111010001"&"0100001100100000",
    869=>"1101000101111100"&"0100101100011001",
    870=>"1100101001000000"&"0101001110000111",
    871=>"1110010101010111"&"0100111010001101",
    872=>"1011010100001101"&"0100111001001011",
    873=>"0000010001001010"&"0100011000000110",
    874=>"1111100100011001"&"0100010010100001",
    875=>"1110101011010110"&"0101010011100010",
    876=>"1011000111111110"&"0101010110100001",
    877=>"1111100001100101"&"0101110101000000",
    878=>"1101011111101011"&"0100011101000110",
    879=>"1111010010001110"&"0101000000101011",
    880=>"1100010100100100"&"0101011101110110",
    881=>"1110000101100100"&"0100011010110001",
    882=>"1101111110000100"&"0101000111101101",
    883=>"1100111100110110"&"0100100111000010",
    884=>"1101000110011010"&"0100011100001001",
    885=>"1101010000111110"&"0100101111010011",
    886=>"1110010010110011"&"0011110111100011",
    887=>"1100001100010001"&"0101110111100001",
    888=>"1110010111011101"&"0101010010111010",
    889=>"1111000001110110"&"0100010110101010",
    890=>"1111110110010111"&"0100011011111101",
    891=>"1100010010110000"&"0101100110010000",
    892=>"1110010010000101"&"0001100001101000",
    893=>"1100100011111011"&"0100110100011011",
    894=>"1101110010001000"&"0101000010001111",
    895=>"1101101101100110"&"0100100100011010",
    896=>"1111101011010011"&"0100100110100001",
    897=>"1110110010000011"&"0101100110111011",
    898=>"1101101001000010"&"0100110110101001",
    899=>"1101100011011000"&"0100011101111011",
    900=>"1110000001011011"&"0100011010001001",
    901=>"1100101101111100"&"0100101111000110",
    902=>"1101100001101110"&"0100101011010111",
    903=>"1110011000100000"&"0100010010100100",
    904=>"1101110111110010"&"0100011100100010",
    905=>"1110100100100001"&"0101011110010011",
    906=>"1011011000111110"&"0101001101111111",
    907=>"1100111111110001"&"0101010100111111",
    908=>"1011111010110000"&"0100111000000001",
    909=>"1110010010000010"&"0101000011001000",
    910=>"1011101111000000"&"0101011000101110",
    911=>"1101110100011111"&"0101000110101101",
    912=>"1110101011100111"&"0101011100011000",
    913=>"1110111110100001"&"0101000011001110",
    914=>"1101100111110001"&"0011010100011111",
    915=>"1110000110010111"&"0100010010100110",
    916=>"1111110100100011"&"0100010111110100",
    917=>"1110111110001010"&"0100100111010111",
    918=>"0000111010101111"&"0101011111001110",
    919=>"1011111101001111"&"0101100100100100",
    920=>"1100101001011101"&"0101010010111001",
    921=>"1001010010001001"&"0100100010011111",
    922=>"1110100000010111"&"0100111010011000",
    923=>"1111010101101001"&"0100010001101000",
    924=>"1101011011111000"&"0101101001101011",
    925=>"1101010011101000"&"0100010100011011",
    926=>"1101011000111110"&"0101000001010000",
    927=>"1111000010101101"&"0101010101010001",
    928=>"1101110111111001"&"0100000110101010",
    929=>"1101110111010001"&"0100110111100010",
    930=>"1101101000011000"&"0101010000011111",
    931=>"1100111110100111"&"0100101000010011",
    932=>"1011111101001110"&"0011111100100100",
    933=>"1010111100011010"&"0110001001000000",
    934=>"1110001001000101"&"0100101011100000",
    935=>"1101110001101101"&"0101001101000001",
    936=>"1101111101010100"&"0100001011100101",
    937=>"1010010101011110"&"0100001000111000",
    938=>"1110101111101000"&"0100110001011011",
    939=>"1101010100110100"&"0101111110101000",
    940=>"1101010000101011"&"0100011100101001",
    941=>"1110000100000101"&"0100100010100101",
    942=>"1101111101101100"&"0100100000010100",
    943=>"1100101010010100"&"0101000100010110",
    944=>"1111011111011111"&"0100101001001011",
    945=>"1011101100000110"&"0100111001011100",
    946=>"1101110101001000"&"0101000111110100",
    947=>"1110111010010111"&"0101001101100101",
    948=>"1101011100000100"&"0101011100100100",
    949=>"1101100110110010"&"0100100110111000",
    950=>"1101000011100000"&"0101001011000011",
    951=>"1110110001000001"&"0100111111100100",
    952=>"1101010110010000"&"0100110100001101",
    953=>"1111111111110111"&"0100101101111101",
    954=>"1110001010110100"&"0100000111101111",
    955=>"1101111100110000"&"0100100110101100",
    956=>"1101011001100100"&"0101001100001110",
    957=>"1111001000100100"&"0100010000011011",
    958=>"1110110001100000"&"0101000011101110",
    959=>"1101101011100101"&"0100111011111100",
    960=>"1110010101011011"&"0101010011100011",
    961=>"1101110000100101"&"0100001011011001",
    962=>"1100110100011010"&"0101100100110100",
    963=>"0000010100110010"&"0100110001101111",
    964=>"1110000010010001"&"0100111011010001",
    965=>"1100100010001001"&"0101100000001100",
    966=>"1111110100101110"&"0011111110101011",
    967=>"0000000111000001"&"0100110010010010",
    968=>"1101011111010011"&"0011101110101000",
    969=>"1101100100110101"&"0100100100101110",
    970=>"1101100100010000"&"0100101101100110",
    971=>"1111010000000101"&"0100101000010100",
    972=>"1101110101000011"&"0100110011000010",
    973=>"1010000111100001"&"0101001101101001",
    974=>"1101101101001101"&"0011101001101010",
    975=>"1110101010000001"&"0100101001000001",
    976=>"1101111111010010"&"0100100010100101",
    977=>"1110000111101110"&"0100011110101101",
    978=>"1110000111001110"&"0101001010100111",
    979=>"1110111111001111"&"0100001100010110",
    980=>"1011111100001110"&"0101000110001010",
    981=>"1101011010101010"&"0100111011011100",
    982=>"1110001011111010"&"0100100101110000",
    983=>"1011011010110110"&"0101000110110001",
    984=>"1110001010110010"&"0100101000111001",
    985=>"1110001100011100"&"0100010010010110",
    986=>"1110001100100111"&"0100101001110110",
    987=>"1100011010100111"&"0100100111000111",
    988=>"1110101111000001"&"0100101010010101",
    989=>"1110101001101101"&"0101010111100111",
    990=>"1101100000000110"&"0101010001110100",
    991=>"1101100010110100"&"0101001011110111",
    992=>"1101100000010110"&"0101000101011111",
    993=>"1101111011100101"&"0100011110010001",
    994=>"1110111001101011"&"0011100111001010",
    995=>"1110100111011011"&"0100000011100000",
    996=>"1101011100100101"&"0010100111000010",
    997=>"1101111101111100"&"0101010100100011",
    998=>"1110010011010011"&"0100110000011110",
    999=>"1110100001110011"&"0100101000010000",
    1000=>"1100010010111001"&"0100011010110101",
    1001=>"1110110000100010"&"0100010101011000",
    1002=>"1110001001011011"&"0100100100110110",
    1003=>"1111001001100011"&"0100010101111100",
    1004=>"1110100110101111"&"0100000111111001",
    1005=>"1110011000000111"&"0100111100101001",
    1006=>"1100110001100100"&"0100001101011100",
    1007=>"1101001101001101"&"0101000001010000",
    1008=>"1111110000001000"&"0100000000101110",
    1009=>"1101111101100000"&"0100110011110000",
    1010=>"1110100110101100"&"0100101100100000",
    1011=>"1100110100111011"&"0100110001011011",
    1012=>"0000111010101000"&"0100110000110100",
    1013=>"1011101001110010"&"0100000111001001",
    1014=>"1110101111010111"&"0100101110111011",
    1015=>"1110001001001000"&"0101001111100100",
    1016=>"1101001010101001"&"0100111111010000",
    1017=>"1110000100101010"&"0100000000111110",
    1018=>"1111011000010100"&"0100110101110101",
    1019=>"1101011111001000"&"0101011101110011",
    1020=>"1111000111100010"&"0100110000001000",
    1021=>"1110110001101111"&"0100111000110000",
    1022=>"1101010111000101"&"0101011101000111",
    1023=>"0000000000011110"&"0100111011101010");
    
BEGIN
    coefs <= ROM_content(to_integer(address));
END RTL;